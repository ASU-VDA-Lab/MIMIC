module fake_ariane_2477_n_367 (n_83, n_8, n_56, n_60, n_64, n_90, n_38, n_47, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_72, n_105, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_93, n_23, n_61, n_102, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_35, n_54, n_25, n_367);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_90;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_72;
input n_105;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_93;
input n_23;
input n_61;
input n_102;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_367;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_347;
wire n_183;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_109;
wire n_245;
wire n_319;
wire n_283;
wire n_187;
wire n_345;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_189;
wire n_286;
wire n_117;
wire n_139;
wire n_130;
wire n_349;
wire n_346;
wire n_214;
wire n_348;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_327;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_339;
wire n_167;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_115;
wire n_320;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_128;
wire n_224;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_108;
wire n_303;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_333;
wire n_221;
wire n_321;
wire n_361;
wire n_149;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_199;
wire n_107;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_343;
wire n_287;
wire n_302;
wire n_284;
wire n_249;
wire n_212;
wire n_123;
wire n_355;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_216;
wire n_223;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_150;
wire n_113;
wire n_114;
wire n_324;
wire n_337;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_159;
wire n_358;
wire n_131;
wire n_263;
wire n_360;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_118;
wire n_121;
wire n_353;
wire n_241;
wire n_357;
wire n_191;
wire n_211;
wire n_322;
wire n_251;
wire n_116;
wire n_351;
wire n_359;
wire n_155;
wire n_127;

INVx1_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_6),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_25),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_14),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_37),
.B(n_29),
.Y(n_115)
);

INVxp33_ASAP7_75t_SL g116 ( 
.A(n_34),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_15),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_23),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_16),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_26),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_42),
.B(n_87),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_3),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_70),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

INVxp33_ASAP7_75t_SL g134 ( 
.A(n_8),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_83),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_20),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_78),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_38),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_32),
.Y(n_146)
);

INVxp33_ASAP7_75t_SL g147 ( 
.A(n_67),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_49),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_31),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_35),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVxp33_ASAP7_75t_SL g154 ( 
.A(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_44),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_12),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_41),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_45),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_21),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_36),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_R g168 ( 
.A(n_108),
.B(n_58),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_0),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_145),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_0),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_112),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_1),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_2),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

OR2x6_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_125),
.Y(n_188)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_117),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_116),
.Y(n_190)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_109),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_182),
.Y(n_192)
);

OR2x6_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_130),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_135),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_175),
.B(n_115),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_117),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_134),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_124),
.B1(n_109),
.B2(n_129),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_129),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_140),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_173),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_179),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_143),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_190),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_200),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_184),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_181),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_142),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_142),
.Y(n_227)
);

AND3x1_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_155),
.C(n_149),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_193),
.A2(n_154),
.B1(n_147),
.B2(n_164),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_201),
.B(n_111),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_160),
.B1(n_157),
.B2(n_158),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_193),
.A2(n_188),
.B1(n_194),
.B2(n_191),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g235 ( 
.A1(n_196),
.A2(n_207),
.B1(n_210),
.B2(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_194),
.B(n_114),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_188),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_204),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_136),
.B1(n_138),
.B2(n_151),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_144),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_153),
.B(n_156),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_195),
.B(n_123),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_117),
.B1(n_163),
.B2(n_162),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_152),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_4),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_5),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_161),
.B(n_159),
.C(n_137),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_214),
.A2(n_133),
.B(n_132),
.C(n_126),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_168),
.B1(n_9),
.B2(n_11),
.Y(n_260)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_7),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_217),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_19),
.B(n_22),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_242),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_233),
.A2(n_24),
.B1(n_33),
.B2(n_39),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_224),
.B(n_40),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_230),
.A2(n_242),
.B1(n_241),
.B2(n_216),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_228),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_231),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_271),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_226),
.B(n_234),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_229),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_243),
.B1(n_235),
.B2(n_232),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_249),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_50),
.Y(n_282)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_265),
.B(n_271),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_51),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_52),
.B(n_53),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_54),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

OA21x2_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_55),
.B(n_56),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_258),
.A2(n_57),
.B(n_59),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_254),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_64),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_282),
.A2(n_273),
.B1(n_266),
.B2(n_261),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_260),
.B(n_273),
.C(n_272),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_285),
.Y(n_301)
);

OAI221xp5_ASAP7_75t_L g302 ( 
.A1(n_276),
.A2(n_267),
.B1(n_264),
.B2(n_248),
.C(n_259),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_253),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_275),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_285),
.Y(n_307)
);

OAI221xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_269),
.B1(n_256),
.B2(n_263),
.C(n_262),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_R g310 ( 
.A1(n_299),
.A2(n_279),
.B(n_280),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

NOR2x1_ASAP7_75t_R g312 ( 
.A(n_305),
.B(n_285),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_303),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_307),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_295),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_298),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_301),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

OAI221xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_302),
.B1(n_286),
.B2(n_294),
.C(n_308),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

NAND4xp25_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_294),
.C(n_277),
.D(n_309),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_263),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_317),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_287),
.Y(n_332)
);

AND2x4_ASAP7_75t_SL g333 ( 
.A(n_321),
.B(n_287),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_322),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_327),
.B(n_292),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_292),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_292),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_284),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_330),
.A2(n_284),
.B1(n_288),
.B2(n_291),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_284),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_284),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_334),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_335),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_283),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_68),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

NOR2x1_ASAP7_75t_R g350 ( 
.A(n_348),
.B(n_343),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_343),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_344),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_351),
.Y(n_354)
);

OAI31xp33_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_349),
.A3(n_345),
.B(n_338),
.Y(n_355)
);

A2O1A1Ixp33_ASAP7_75t_L g356 ( 
.A1(n_353),
.A2(n_339),
.B(n_350),
.C(n_340),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_333),
.B1(n_341),
.B2(n_326),
.Y(n_357)
);

AOI311xp33_ASAP7_75t_L g358 ( 
.A1(n_355),
.A2(n_347),
.A3(n_326),
.B(n_336),
.C(n_291),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_357),
.B(n_347),
.Y(n_359)
);

NAND4xp25_ASAP7_75t_SL g360 ( 
.A(n_358),
.B(n_337),
.C(n_291),
.D(n_341),
.Y(n_360)
);

NOR3x1_ASAP7_75t_L g361 ( 
.A(n_359),
.B(n_278),
.C(n_71),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_361),
.Y(n_362)
);

AOI221xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_360),
.B1(n_73),
.B2(n_74),
.C(n_77),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_363),
.A2(n_69),
.B1(n_79),
.B2(n_81),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_364),
.A2(n_82),
.B(n_84),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_365),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_96),
.B(n_98),
.Y(n_367)
);


endmodule