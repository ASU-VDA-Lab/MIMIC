module fake_netlist_1_6137_n_717 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_717);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_717;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx2_ASAP7_75t_L g87 ( .A(n_74), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_31), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_26), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_7), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_67), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_12), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_25), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_40), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_33), .Y(n_96) );
BUFx10_ASAP7_75t_L g97 ( .A(n_84), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_2), .Y(n_98) );
BUFx5_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_36), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_57), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_62), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_59), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_19), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_64), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_60), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_61), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_29), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_11), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_53), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_72), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_69), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_32), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_11), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_56), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_101), .Y(n_124) );
NOR2x1_ASAP7_75t_L g125 ( .A(n_90), .B(n_0), .Y(n_125) );
AND2x6_ASAP7_75t_L g126 ( .A(n_95), .B(n_20), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_100), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_106), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_103), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_95), .B(n_0), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_88), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_131) );
INVx6_ASAP7_75t_L g132 ( .A(n_97), .Y(n_132) );
INVx5_ASAP7_75t_L g133 ( .A(n_101), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_107), .B(n_1), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_97), .B(n_3), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_116), .B(n_113), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_101), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_104), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_97), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_117), .B(n_4), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_116), .B(n_4), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_105), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
INVx4_ASAP7_75t_SL g145 ( .A(n_126), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_124), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_137), .A2(n_93), .B1(n_110), .B2(n_109), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_124), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_135), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_130), .B(n_119), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_137), .A2(n_93), .B1(n_101), .B2(n_99), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_135), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_124), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
INVxp33_ASAP7_75t_SL g157 ( .A(n_123), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_126), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
OR2x2_ASAP7_75t_L g161 ( .A(n_123), .B(n_98), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
INVxp33_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_127), .B(n_129), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_128), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
OAI21xp33_ASAP7_75t_SL g167 ( .A1(n_127), .A2(n_94), .B(n_99), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_140), .B(n_93), .Y(n_169) );
NOR3xp33_ASAP7_75t_L g170 ( .A(n_134), .B(n_121), .C(n_122), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_129), .B(n_99), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_140), .B(n_89), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
NOR2xp33_ASAP7_75t_SL g176 ( .A(n_126), .B(n_88), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_140), .B(n_92), .Y(n_177) );
OR2x2_ASAP7_75t_L g178 ( .A(n_140), .B(n_93), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_132), .B(n_99), .Y(n_179) );
NOR3xp33_ASAP7_75t_L g180 ( .A(n_141), .B(n_120), .C(n_118), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_168), .B(n_132), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_168), .B(n_132), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_163), .B(n_139), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_161), .B(n_136), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_178), .Y(n_185) );
NAND3xp33_ASAP7_75t_SL g186 ( .A(n_165), .B(n_131), .C(n_114), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_157), .B(n_139), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_168), .B(n_143), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_146), .B(n_142), .Y(n_189) );
NAND2x1_ASAP7_75t_L g190 ( .A(n_151), .B(n_126), .Y(n_190) );
INVx8_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_170), .A2(n_142), .B1(n_114), .B2(n_144), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_151), .A2(n_126), .B1(n_143), .B2(n_144), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_161), .A2(n_91), .B1(n_125), .B2(n_102), .Y(n_194) );
INVx8_ASAP7_75t_L g195 ( .A(n_151), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_146), .B(n_99), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_168), .B(n_126), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_172), .B(n_125), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_178), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_172), .B(n_96), .Y(n_200) );
NOR3xp33_ASAP7_75t_L g201 ( .A(n_170), .B(n_111), .C(n_112), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_151), .A2(n_91), .B1(n_115), .B2(n_133), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_172), .B(n_133), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_174), .B(n_133), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_146), .B(n_133), .Y(n_205) );
O2A1O1Ixp5_ASAP7_75t_L g206 ( .A1(n_146), .A2(n_133), .B(n_138), .C(n_45), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_150), .Y(n_207) );
INVxp33_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_175), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_179), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_172), .B(n_133), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_178), .Y(n_212) );
BUFx8_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_179), .B(n_138), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_171), .B(n_5), .Y(n_216) );
OAI22xp33_ASAP7_75t_L g217 ( .A1(n_176), .A2(n_138), .B1(n_6), .B2(n_7), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_179), .B(n_138), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_153), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_151), .B(n_138), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
BUFx2_ASAP7_75t_L g222 ( .A(n_213), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_190), .B(n_159), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_187), .A2(n_176), .B1(n_151), .B2(n_180), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_184), .B(n_180), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_183), .A2(n_160), .B(n_158), .C(n_154), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_197), .A2(n_159), .B(n_154), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_208), .B(n_177), .Y(n_228) );
NOR2x1_ASAP7_75t_L g229 ( .A(n_186), .B(n_164), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_207), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_184), .B(n_151), .Y(n_231) );
NOR2xp67_ASAP7_75t_L g232 ( .A(n_192), .B(n_167), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_SL g233 ( .A1(n_201), .A2(n_158), .B(n_160), .C(n_152), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_208), .B(n_167), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_210), .B(n_164), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_185), .B(n_145), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_199), .B(n_169), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_212), .B(n_169), .Y(n_238) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_196), .A2(n_158), .B(n_160), .C(n_169), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_213), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_191), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_198), .B(n_158), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_189), .B(n_145), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_189), .B(n_160), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_220), .A2(n_171), .B(n_152), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_188), .A2(n_148), .B(n_159), .C(n_166), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_193), .B(n_145), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_196), .A2(n_145), .B(n_148), .Y(n_248) );
NAND3xp33_ASAP7_75t_L g249 ( .A(n_202), .B(n_216), .C(n_213), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_205), .A2(n_145), .B(n_173), .Y(n_250) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_206), .A2(n_156), .B(n_173), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_191), .A2(n_175), .B1(n_145), .B2(n_166), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_207), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_209), .B(n_175), .Y(n_254) );
NOR2xp67_ASAP7_75t_L g255 ( .A(n_232), .B(n_216), .Y(n_255) );
INVx3_ASAP7_75t_SL g256 ( .A(n_240), .Y(n_256) );
AO21x1_ASAP7_75t_L g257 ( .A1(n_234), .A2(n_217), .B(n_218), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_225), .B(n_194), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_251), .A2(n_214), .B(n_219), .Y(n_259) );
AO22x2_ASAP7_75t_L g260 ( .A1(n_249), .A2(n_221), .B1(n_219), .B2(n_215), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_234), .A2(n_221), .B1(n_215), .B2(n_182), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
AOI22xp33_ASAP7_75t_SL g263 ( .A1(n_222), .A2(n_191), .B1(n_195), .B2(n_209), .Y(n_263) );
INVx5_ASAP7_75t_L g264 ( .A(n_241), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g265 ( .A(n_240), .B(n_191), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_228), .B(n_200), .Y(n_266) );
BUFx8_ASAP7_75t_L g267 ( .A(n_241), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_224), .A2(n_195), .B1(n_181), .B2(n_203), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_230), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_238), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_226), .A2(n_204), .B(n_195), .C(n_211), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_253), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_250), .A2(n_205), .B(n_173), .Y(n_273) );
OAI22xp5_ASAP7_75t_SL g274 ( .A1(n_228), .A2(n_195), .B1(n_6), .B2(n_8), .Y(n_274) );
NAND3xp33_ASAP7_75t_SL g275 ( .A(n_233), .B(n_166), .C(n_162), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_231), .B(n_175), .Y(n_276) );
AOI21x1_ASAP7_75t_L g277 ( .A1(n_260), .A2(n_247), .B(n_227), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_259), .A2(n_245), .B(n_252), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_272), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_271), .A2(n_233), .B(n_247), .Y(n_280) );
AND2x6_ASAP7_75t_L g281 ( .A(n_269), .B(n_241), .Y(n_281) );
BUFx8_ASAP7_75t_SL g282 ( .A(n_262), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_270), .B(n_244), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_257), .A2(n_239), .B(n_248), .Y(n_285) );
INVx4_ASAP7_75t_L g286 ( .A(n_264), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_258), .A2(n_229), .B1(n_244), .B2(n_242), .Y(n_287) );
AO31x2_ASAP7_75t_L g288 ( .A1(n_268), .A2(n_242), .A3(n_235), .B(n_149), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_255), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_264), .B(n_254), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_275), .A2(n_266), .B(n_246), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_267), .B(n_243), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_275), .A2(n_254), .B(n_243), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_261), .A2(n_162), .B(n_156), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_256), .A2(n_236), .B(n_223), .C(n_156), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_261), .B(n_236), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_273), .A2(n_162), .B(n_155), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_299), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_279), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_299), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_280), .A2(n_276), .B(n_155), .Y(n_304) );
AO21x1_ASAP7_75t_SL g305 ( .A1(n_297), .A2(n_264), .B(n_274), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_297), .B(n_256), .Y(n_307) );
INVxp67_ASAP7_75t_SL g308 ( .A(n_295), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_300), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_279), .B(n_263), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_288), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_290), .B(n_265), .Y(n_312) );
OA21x2_ASAP7_75t_L g313 ( .A1(n_278), .A2(n_155), .B(n_149), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_285), .B(n_263), .Y(n_314) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_292), .A2(n_276), .B(n_149), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_295), .A2(n_223), .B(n_265), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_298), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_286), .Y(n_320) );
NOR2xp33_ASAP7_75t_SL g321 ( .A(n_286), .B(n_241), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_282), .B(n_175), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_285), .B(n_5), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
OAI21x1_ASAP7_75t_L g325 ( .A1(n_278), .A2(n_147), .B(n_47), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_285), .B(n_8), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_295), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_288), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_281), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_284), .B(n_9), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_285), .B(n_10), .Y(n_333) );
AO21x2_ASAP7_75t_L g334 ( .A1(n_277), .A2(n_10), .B(n_12), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_300), .B(n_288), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_300), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_284), .B(n_13), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_289), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_289), .B(n_14), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_335), .B(n_288), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_317), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_335), .B(n_288), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_335), .B(n_283), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_301), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_317), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_319), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_319), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_331), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_324), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_302), .B(n_287), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_336), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_323), .B(n_277), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_330), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_286), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_310), .B(n_294), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_303), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_323), .B(n_326), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_331), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_326), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_326), .B(n_286), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_325), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_333), .B(n_283), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_14), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_333), .B(n_15), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_303), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_320), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_303), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_316), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_314), .B(n_15), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_316), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_327), .Y(n_382) );
NOR2x1_ASAP7_75t_R g383 ( .A(n_320), .B(n_293), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_307), .B(n_291), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_314), .B(n_16), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_327), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_327), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_331), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_310), .B(n_281), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_328), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_328), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_307), .B(n_16), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_306), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_328), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_314), .B(n_17), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_306), .B(n_17), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_310), .B(n_281), .Y(n_397) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_334), .B(n_296), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_311), .B(n_281), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_329), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_338), .B(n_18), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_312), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_312), .B(n_281), .Y(n_403) );
INVx5_ASAP7_75t_L g404 ( .A(n_312), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_338), .B(n_18), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_358), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_348), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_343), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_365), .B(n_311), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_365), .B(n_329), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_358), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_342), .B(n_368), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_343), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_340), .B(n_329), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_403), .B(n_312), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_342), .B(n_308), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_379), .B(n_332), .Y(n_417) );
NOR2xp67_ASAP7_75t_L g418 ( .A(n_404), .B(n_322), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_348), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_379), .B(n_332), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_341), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_368), .B(n_308), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_340), .B(n_334), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_341), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_348), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_381), .B(n_339), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_385), .B(n_337), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_345), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g429 ( .A1(n_404), .A2(n_321), .B1(n_334), .B2(n_281), .Y(n_429) );
CKINVDCx14_ASAP7_75t_R g430 ( .A(n_371), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_344), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_362), .B(n_334), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_345), .Y(n_433) );
AND2x4_ASAP7_75t_L g434 ( .A(n_403), .B(n_312), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_346), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_362), .B(n_334), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_361), .B(n_315), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_385), .B(n_337), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_403), .B(n_312), .Y(n_440) );
OR2x6_ASAP7_75t_SL g441 ( .A(n_396), .B(n_305), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_380), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_361), .B(n_315), .Y(n_443) );
BUFx3_ASAP7_75t_L g444 ( .A(n_375), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_404), .B(n_321), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_355), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_346), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_369), .B(n_315), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_347), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_369), .B(n_315), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_347), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_357), .B(n_315), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_352), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_403), .B(n_304), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_352), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_357), .B(n_304), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_404), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_353), .B(n_304), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_364), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_380), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_371), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_393), .B(n_304), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_353), .B(n_304), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_393), .B(n_339), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_364), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_380), .B(n_305), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_356), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_359), .B(n_305), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_383), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_359), .B(n_313), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_396), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_395), .B(n_281), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_344), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_383), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_404), .B(n_318), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_404), .B(n_318), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_360), .B(n_313), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_395), .B(n_19), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_392), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_360), .B(n_313), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_367), .B(n_313), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_392), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_356), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_367), .B(n_313), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_344), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_377), .B(n_325), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_377), .B(n_325), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_401), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_402), .A2(n_147), .B1(n_23), .B2(n_24), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_401), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_378), .B(n_22), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_405), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_404), .B(n_27), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_389), .B(n_28), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_405), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_350), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_372), .B(n_30), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_446), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_408), .B(n_389), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_461), .B(n_397), .Y(n_500) );
AND2x2_ASAP7_75t_SL g501 ( .A(n_469), .B(n_373), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_413), .B(n_414), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_430), .B(n_349), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_412), .B(n_409), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_406), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_412), .B(n_366), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_409), .B(n_366), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_458), .B(n_386), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_426), .B(n_384), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_444), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_479), .B(n_354), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_406), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_416), .B(n_388), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_431), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_416), .B(n_386), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_410), .B(n_388), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_411), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_421), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_458), .B(n_354), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_410), .B(n_382), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_424), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_428), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_419), .B(n_399), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_433), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_482), .B(n_399), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_435), .Y(n_526) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_418), .B(n_398), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_464), .B(n_376), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_419), .B(n_382), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_425), .B(n_376), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_471), .B(n_376), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_415), .B(n_387), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_415), .B(n_387), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_447), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_463), .B(n_374), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_449), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_451), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_407), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_453), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_407), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_438), .B(n_374), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_455), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_467), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_469), .A2(n_398), .B(n_374), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_463), .B(n_350), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_488), .B(n_490), .Y(n_546) );
OR2x6_ASAP7_75t_L g547 ( .A(n_474), .B(n_350), .Y(n_547) );
OR2x6_ASAP7_75t_L g548 ( .A(n_474), .B(n_363), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_483), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_492), .B(n_363), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_459), .B(n_351), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_432), .B(n_351), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_459), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_457), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_432), .B(n_400), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_465), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_465), .B(n_400), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_443), .B(n_400), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_495), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_423), .B(n_394), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_448), .B(n_394), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_431), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_436), .B(n_394), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_436), .B(n_391), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_452), .B(n_391), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_452), .B(n_391), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_422), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_456), .B(n_390), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_422), .Y(n_569) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_429), .A2(n_390), .B(n_370), .Y(n_570) );
NAND2x1_ASAP7_75t_L g571 ( .A(n_466), .B(n_370), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_450), .B(n_370), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_473), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_485), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_496), .Y(n_575) );
AND3x1_ASAP7_75t_L g576 ( .A(n_466), .B(n_370), .C(n_34), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_496), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_450), .B(n_370), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_441), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_504), .B(n_456), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_503), .B(n_468), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_506), .B(n_468), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_519), .B(n_427), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_519), .B(n_439), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_502), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_540), .B(n_454), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_543), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_515), .B(n_462), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_540), .B(n_478), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_498), .B(n_417), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_507), .B(n_454), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_549), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_579), .A2(n_441), .B1(n_420), .B2(n_475), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_520), .B(n_437), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_538), .B(n_415), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_547), .B(n_454), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_501), .A2(n_434), .B1(n_440), .B2(n_445), .Y(n_597) );
AOI222xp33_ASAP7_75t_L g598 ( .A1(n_509), .A2(n_434), .B1(n_440), .B2(n_457), .C1(n_497), .C2(n_476), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_517), .Y(n_599) );
NOR2xp67_ASAP7_75t_SL g600 ( .A(n_554), .B(n_494), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_511), .B(n_486), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_565), .B(n_460), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_516), .B(n_523), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_576), .A2(n_434), .B1(n_440), .B2(n_472), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_567), .B(n_569), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g606 ( .A1(n_544), .A2(n_494), .B(n_493), .C(n_475), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_559), .B(n_486), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_565), .B(n_460), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_513), .B(n_460), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_525), .B(n_487), .Y(n_610) );
OAI21xp5_ASAP7_75t_L g611 ( .A1(n_576), .A2(n_493), .B(n_491), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_551), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_510), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_546), .B(n_437), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_566), .B(n_442), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_570), .A2(n_442), .B(n_437), .C(n_487), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_541), .B(n_480), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_528), .B(n_475), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_518), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_521), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_566), .B(n_480), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_557), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_553), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_522), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_544), .A2(n_493), .B(n_489), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_558), .B(n_484), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_524), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_568), .B(n_484), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_526), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_568), .B(n_481), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_529), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_552), .B(n_481), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_561), .B(n_477), .Y(n_633) );
A2O1A1O1Ixp25_ASAP7_75t_L g634 ( .A1(n_570), .A2(n_370), .B(n_477), .C(n_470), .D(n_38), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_552), .B(n_470), .Y(n_635) );
OAI22xp33_ASAP7_75t_SL g636 ( .A1(n_547), .A2(n_35), .B1(n_37), .B2(n_39), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_534), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_556), .A2(n_147), .B(n_42), .Y(n_638) );
OAI32xp33_ASAP7_75t_L g639 ( .A1(n_593), .A2(n_527), .A3(n_499), .B1(n_508), .B2(n_500), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_597), .A2(n_547), .B1(n_548), .B2(n_527), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_602), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_599), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_596), .B(n_548), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_619), .Y(n_644) );
AOI321xp33_ASAP7_75t_L g645 ( .A1(n_597), .A2(n_578), .A3(n_572), .B1(n_532), .B2(n_533), .C(n_555), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_634), .B(n_548), .C(n_531), .Y(n_646) );
NOR2xp67_ASAP7_75t_SL g647 ( .A(n_611), .B(n_562), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_608), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_615), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_583), .B(n_542), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_586), .B(n_533), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_587), .B(n_508), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_598), .A2(n_532), .B1(n_555), .B2(n_564), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_620), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_634), .A2(n_539), .B(n_536), .C(n_537), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_598), .A2(n_563), .B1(n_564), .B2(n_545), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_612), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_611), .A2(n_571), .B(n_550), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_584), .A2(n_563), .B(n_535), .Y(n_659) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_604), .B(n_545), .C(n_535), .D(n_560), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_594), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_636), .A2(n_574), .B(n_573), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_636), .A2(n_530), .B(n_505), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_585), .B(n_512), .Y(n_664) );
OAI21xp33_ASAP7_75t_L g665 ( .A1(n_601), .A2(n_577), .B(n_575), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_606), .A2(n_514), .B(n_147), .C(n_43), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_607), .B(n_624), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_623), .B(n_41), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_604), .A2(n_147), .B1(n_44), .B2(n_46), .C(n_50), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_589), .A2(n_147), .B1(n_51), .B2(n_52), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_627), .Y(n_671) );
BUFx4f_ASAP7_75t_SL g672 ( .A(n_581), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_655), .A2(n_592), .B(n_590), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_639), .A2(n_637), .B1(n_629), .B2(n_595), .C(n_613), .Y(n_674) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_662), .A2(n_625), .B(n_600), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_663), .A2(n_638), .B(n_616), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_662), .A2(n_638), .B(n_618), .C(n_614), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_672), .A2(n_588), .B1(n_596), .B2(n_580), .Y(n_678) );
AOI311xp33_ASAP7_75t_L g679 ( .A1(n_640), .A2(n_610), .A3(n_605), .B(n_617), .C(n_626), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_656), .B(n_603), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_660), .A2(n_622), .B1(n_631), .B2(n_582), .C(n_591), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_659), .A2(n_609), .B1(n_633), .B2(n_632), .C(n_635), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_663), .A2(n_630), .B(n_628), .C(n_621), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_653), .A2(n_147), .B1(n_54), .B2(n_58), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_646), .B(n_63), .Y(n_685) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_647), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_650), .B(n_66), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_665), .A2(n_68), .B1(n_70), .B2(n_73), .C(n_75), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_658), .A2(n_76), .B1(n_78), .B2(n_79), .C(n_80), .Y(n_689) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_645), .A2(n_81), .B(n_82), .C(n_83), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_667), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_658), .B(n_85), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_667), .A2(n_86), .B1(n_652), .B2(n_642), .C(n_644), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_666), .A2(n_669), .B(n_670), .C(n_664), .Y(n_694) );
AOI221x1_ASAP7_75t_L g695 ( .A1(n_668), .A2(n_654), .B1(n_671), .B2(n_643), .C(n_649), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_643), .A2(n_657), .B(n_648), .C(n_641), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g697 ( .A1(n_651), .A2(n_640), .B(n_663), .C(n_662), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_661), .B(n_669), .C(n_662), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_673), .B(n_691), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_697), .A2(n_675), .B1(n_683), .B2(n_674), .C(n_686), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_680), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_685), .B(n_689), .C(n_694), .Y(n_702) );
NOR2xp67_ASAP7_75t_L g703 ( .A(n_676), .B(n_677), .Y(n_703) );
AOI211x1_ASAP7_75t_L g704 ( .A1(n_701), .A2(n_678), .B(n_679), .C(n_692), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_703), .B(n_690), .C(n_688), .Y(n_705) );
NAND4xp75_ASAP7_75t_L g706 ( .A(n_700), .B(n_695), .C(n_684), .D(n_687), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_704), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_706), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_708), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_708), .Y(n_710) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_709), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_711), .Y(n_713) );
OAI21x1_ASAP7_75t_SL g714 ( .A1(n_713), .A2(n_712), .B(n_707), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_SL g715 ( .A1(n_714), .A2(n_699), .B(n_696), .C(n_705), .Y(n_715) );
AO21x2_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_702), .B(n_698), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_681), .B1(n_682), .B2(n_693), .Y(n_717) );
endmodule