module fake_netlist_6_2931_n_1565 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1565);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1565;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_142;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_141;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_140;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_167;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_143;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_67),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

BUFx8_ASAP7_75t_SL g143 ( 
.A(n_119),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_44),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_42),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_45),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_14),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_73),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_28),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_36),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_78),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_40),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_84),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_33),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_7),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_22),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_112),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_89),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_79),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_76),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_74),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_132),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_26),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_28),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_3),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_72),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_136),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_62),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_69),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_47),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_41),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_12),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_113),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_63),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_51),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_97),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_101),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_1),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_30),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_99),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_30),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_3),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_87),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_31),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_38),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_68),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_129),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_24),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_122),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_20),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_61),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_15),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_54),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_22),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_13),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_27),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_43),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_128),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_23),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_52),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_39),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_11),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_65),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_34),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_85),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_6),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_12),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_10),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_15),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_75),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_34),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_0),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_13),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_137),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_32),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_48),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_60),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_46),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_123),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_19),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_29),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_33),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_96),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_107),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_29),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_105),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_126),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_6),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_8),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_82),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_90),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_20),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_56),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_21),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_55),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_16),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_50),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_80),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_100),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_86),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_58),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_114),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_71),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_25),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_229),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_142),
.Y(n_283)
);

BUFx6f_ASAP7_75t_SL g284 ( 
.A(n_185),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_229),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_274),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_229),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_229),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_197),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_213),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_251),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_146),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_198),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_147),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_159),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_147),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_152),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_157),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_180),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_216),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_168),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_170),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_147),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_147),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_177),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_211),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_171),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_278),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_175),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_220),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_251),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_146),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_171),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_232),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_236),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_188),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_256),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_237),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_268),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_189),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_144),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_155),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_144),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_191),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_268),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_177),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_177),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_177),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_275),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_155),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_169),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_307),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_199),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_183),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_303),
.B(n_140),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_289),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_307),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_169),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_303),
.B(n_230),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_306),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_289),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_R g363 ( 
.A(n_312),
.B(n_275),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_141),
.Y(n_365)
);

BUFx8_ASAP7_75t_L g366 ( 
.A(n_284),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_281),
.B(n_185),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_230),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_300),
.B(n_151),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_288),
.B(n_151),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_308),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_300),
.B(n_185),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_282),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_285),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_290),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_290),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_173),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g380 ( 
.A1(n_341),
.A2(n_292),
.B(n_291),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_313),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_291),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_283),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_294),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_292),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_293),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_293),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_313),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_297),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_297),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_299),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_299),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_302),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_302),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_173),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_281),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_304),
.B(n_145),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_305),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_305),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g401 ( 
.A(n_287),
.B(n_238),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_318),
.B(n_264),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_301),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_316),
.B(n_264),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_317),
.B(n_148),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_344),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_320),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_286),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_344),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_326),
.B(n_149),
.Y(n_413)
);

CKINVDCx8_ASAP7_75t_R g414 ( 
.A(n_396),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_373),
.B(n_276),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_359),
.B(n_276),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_357),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_359),
.B(n_320),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_363),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_327),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_150),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_383),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_397),
.B(n_150),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_364),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_371),
.B(n_150),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_364),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_367),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_365),
.B(n_327),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_371),
.B(n_150),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

OR2x6_ASAP7_75t_L g441 ( 
.A(n_410),
.B(n_310),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_365),
.B(n_333),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_411),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_408),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_375),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_386),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_371),
.B(n_192),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_377),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_384),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_377),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_372),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_354),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_401),
.B(n_298),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_353),
.B(n_382),
.Y(n_456)
);

OAI22xp33_ASAP7_75t_L g457 ( 
.A1(n_372),
.A2(n_295),
.B1(n_241),
.B2(n_239),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_R g458 ( 
.A(n_381),
.B(n_311),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_353),
.B(n_333),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_361),
.B(n_342),
.Y(n_464)
);

AND3x2_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_208),
.C(n_154),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_357),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_407),
.B(n_342),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_369),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_354),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_369),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_369),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_407),
.B(n_284),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_394),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_371),
.B(n_192),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_368),
.B(n_321),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_386),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_403),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_405),
.B(n_192),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_413),
.B(n_284),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_380),
.A2(n_405),
.B1(n_391),
.B2(n_400),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_405),
.B(n_192),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_R g487 ( 
.A(n_388),
.B(n_319),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_409),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_357),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_366),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_370),
.B(n_337),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_366),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_405),
.B(n_263),
.Y(n_494)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_366),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_393),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_386),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_357),
.B(n_329),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_413),
.B(n_286),
.Y(n_500)
);

NOR2x1p5_ASAP7_75t_L g501 ( 
.A(n_366),
.B(n_207),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_412),
.B(n_331),
.Y(n_502)
);

NAND3xp33_ASAP7_75t_L g503 ( 
.A(n_351),
.B(n_218),
.C(n_217),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_378),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_378),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_376),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_378),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_386),
.Y(n_508)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_370),
.B(n_263),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_378),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_376),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_370),
.B(n_263),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_399),
.B(n_336),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_374),
.B(n_263),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_408),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_408),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_399),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_356),
.B(n_338),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_374),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_387),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_374),
.Y(n_525)
);

NOR2x1p5_ASAP7_75t_L g526 ( 
.A(n_406),
.B(n_222),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_374),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_374),
.B(n_273),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_374),
.Y(n_529)
);

NAND3xp33_ASAP7_75t_L g530 ( 
.A(n_356),
.B(n_244),
.C(n_243),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_387),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_380),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_387),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_387),
.B(n_205),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_352),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_387),
.B(n_273),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_379),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_387),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_389),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_352),
.A2(n_172),
.B1(n_279),
.B2(n_200),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_389),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_389),
.B(n_273),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_389),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_389),
.B(n_156),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_350),
.B(n_338),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_392),
.Y(n_547)
);

AND3x2_ASAP7_75t_L g548 ( 
.A(n_379),
.B(n_153),
.C(n_209),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_402),
.B(n_322),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_392),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_402),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_423),
.B(n_380),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_454),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_420),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_423),
.B(n_380),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_485),
.B(n_392),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_467),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_419),
.B(n_380),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_417),
.B(n_177),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_419),
.B(n_392),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_438),
.B(n_392),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_424),
.B(n_469),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_438),
.B(n_392),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_532),
.B(n_398),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_489),
.Y(n_568)
);

NOR3xp33_ASAP7_75t_L g569 ( 
.A(n_421),
.B(n_500),
.C(n_503),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_451),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_451),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_426),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_532),
.B(n_398),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_468),
.B(n_247),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_476),
.B(n_482),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_476),
.B(n_482),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_456),
.B(n_398),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_470),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_468),
.B(n_398),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_537),
.B(n_398),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_489),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_435),
.B(n_398),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

AND2x6_ASAP7_75t_SL g584 ( 
.A(n_441),
.B(n_478),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_551),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_435),
.B(n_379),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_442),
.B(n_160),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_455),
.B(n_406),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_442),
.B(n_252),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_422),
.B(n_143),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_471),
.B(n_273),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_535),
.B(n_395),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_415),
.B(n_395),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_445),
.B(n_395),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_460),
.B(n_261),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_472),
.B(n_177),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_500),
.B(n_269),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_424),
.A2(n_210),
.B1(n_262),
.B2(n_226),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_450),
.B(n_402),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_464),
.B(n_277),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_452),
.B(n_350),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_519),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_453),
.B(n_210),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_526),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_504),
.A2(n_228),
.B(n_162),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_519),
.B(n_177),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_549),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_521),
.B(n_158),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_502),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_459),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_462),
.B(n_143),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_466),
.B(n_355),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_491),
.B(n_358),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_496),
.B(n_161),
.Y(n_615)
);

INVx8_ASAP7_75t_L g616 ( 
.A(n_417),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_498),
.B(n_163),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_418),
.B(n_491),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_491),
.B(n_360),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_427),
.B(n_328),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_521),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_505),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_478),
.A2(n_418),
.B1(n_484),
.B2(n_473),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_513),
.A2(n_484),
.B(n_473),
.C(n_507),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_534),
.B(n_510),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_513),
.B(n_164),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_520),
.B(n_165),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_417),
.B(n_176),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_417),
.B(n_428),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_441),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_417),
.B(n_184),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_428),
.A2(n_262),
.B1(n_224),
.B2(n_242),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_533),
.B(n_186),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_533),
.B(n_190),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_539),
.B(n_204),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_502),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_416),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_429),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_478),
.B(n_166),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_425),
.B(n_214),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_441),
.B(n_330),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_425),
.B(n_215),
.Y(n_643)
);

NOR2xp67_ASAP7_75t_L g644 ( 
.A(n_490),
.B(n_360),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_425),
.B(n_223),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_512),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_488),
.B(n_414),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_546),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_432),
.A2(n_246),
.B1(n_259),
.B2(n_235),
.Y(n_649)
);

BUFx6f_ASAP7_75t_SL g650 ( 
.A(n_522),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_425),
.B(n_240),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_425),
.B(n_245),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_440),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_430),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_465),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_444),
.B(n_248),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_509),
.B(n_167),
.Y(n_657)
);

BUFx12f_ASAP7_75t_SL g658 ( 
.A(n_522),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_509),
.B(n_174),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_539),
.B(n_249),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_530),
.B(n_178),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_546),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_522),
.B(n_318),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_517),
.A2(n_255),
.B(n_258),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_545),
.A2(n_345),
.B(n_346),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_490),
.B(n_332),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_548),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_547),
.B(n_179),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_547),
.B(n_181),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_457),
.B(n_182),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_432),
.Y(n_671)
);

OAI22x1_ASAP7_75t_SL g672 ( 
.A1(n_488),
.A2(n_347),
.B1(n_343),
.B2(n_231),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_458),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_506),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_492),
.B(n_187),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_458),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_440),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_487),
.B(n_324),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_506),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_431),
.Y(n_680)
);

NOR2xp67_ASAP7_75t_L g681 ( 
.A(n_481),
.B(n_193),
.Y(n_681)
);

AND2x2_ASAP7_75t_SL g682 ( 
.A(n_550),
.B(n_345),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_511),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_481),
.A2(n_346),
.B(n_233),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_486),
.B(n_201),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_440),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_437),
.A2(n_449),
.B1(n_477),
.B2(n_509),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_511),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_540),
.B(n_544),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_497),
.B(n_250),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_433),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_531),
.B(n_206),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_487),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_434),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_497),
.B(n_260),
.Y(n_695)
);

A2O1A1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_474),
.A2(n_475),
.B(n_483),
.C(n_486),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_437),
.B(n_194),
.C(n_196),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_440),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_574),
.A2(n_589),
.B(n_598),
.C(n_618),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_608),
.Y(n_700)
);

BUFx12f_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_588),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_623),
.B(n_515),
.Y(n_703)
);

CKINVDCx6p67_ASAP7_75t_R g704 ( 
.A(n_572),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_553),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_552),
.B(n_474),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_629),
.B(n_495),
.Y(n_707)
);

BUFx5_ASAP7_75t_L g708 ( 
.A(n_682),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_553),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_574),
.B(n_495),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_570),
.Y(n_712)
);

NOR2x2_ASAP7_75t_L g713 ( 
.A(n_599),
.B(n_633),
.Y(n_713)
);

NOR2x2_ASAP7_75t_L g714 ( 
.A(n_599),
.B(n_495),
.Y(n_714)
);

NAND2x1p5_ASAP7_75t_L g715 ( 
.A(n_581),
.B(n_448),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_611),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_589),
.B(n_541),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_558),
.A2(n_494),
.B(n_448),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_557),
.B(n_475),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_586),
.B(n_515),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_565),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_653),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_648),
.B(n_483),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_649),
.A2(n_501),
.B1(n_494),
.B2(n_477),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_680),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_598),
.B(n_508),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_569),
.A2(n_449),
.B1(n_509),
.B2(n_523),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_678),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_662),
.B(n_434),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_569),
.B(n_515),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_649),
.A2(n_509),
.B1(n_525),
.B2(n_527),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_618),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_581),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_653),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_595),
.A2(n_517),
.B(n_529),
.C(n_538),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_614),
.B(n_508),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_653),
.Y(n_737)
);

INVx5_ASAP7_75t_L g738 ( 
.A(n_616),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_592),
.Y(n_739)
);

BUFx12f_ASAP7_75t_L g740 ( 
.A(n_655),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_620),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_616),
.B(n_515),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_622),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_680),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_597),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_663),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_571),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_597),
.B(n_516),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_689),
.A2(n_436),
.B1(n_439),
.B2(n_443),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_610),
.B(n_436),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_610),
.B(n_439),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_601),
.B(n_334),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_693),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_637),
.B(n_443),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_555),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_556),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_658),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_559),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_653),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_686),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_568),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_616),
.B(n_516),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_673),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_SL g764 ( 
.A(n_604),
.B(n_266),
.C(n_221),
.Y(n_764)
);

AND2x6_ASAP7_75t_L g765 ( 
.A(n_630),
.B(n_646),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_579),
.B(n_446),
.Y(n_766)
);

NOR2x1_ASAP7_75t_L g767 ( 
.A(n_644),
.B(n_524),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_601),
.B(n_335),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_582),
.B(n_446),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_638),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_558),
.B(n_447),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_603),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_560),
.B(n_624),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_577),
.B(n_447),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_603),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_585),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_577),
.B(n_543),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_595),
.B(n_543),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_670),
.B(n_538),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_603),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_670),
.B(n_524),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_676),
.B(n_516),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_593),
.B(n_448),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_567),
.A2(n_542),
.B(n_536),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_674),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_614),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_647),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_594),
.B(n_493),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_587),
.B(n_493),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_600),
.B(n_493),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_679),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_683),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_619),
.B(n_335),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_686),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_663),
.B(n_518),
.Y(n_795)
);

O2A1O1Ixp5_ASAP7_75t_L g796 ( 
.A1(n_596),
.A2(n_626),
.B(n_625),
.C(n_591),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_619),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_688),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_639),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_671),
.B(n_518),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_682),
.B(n_518),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_603),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_575),
.B(n_518),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_691),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_689),
.A2(n_542),
.B1(n_536),
.B2(n_528),
.Y(n_805)
);

AND2x6_ASAP7_75t_L g806 ( 
.A(n_621),
.B(n_227),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_605),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_576),
.B(n_528),
.Y(n_808)
);

INVx5_ASAP7_75t_L g809 ( 
.A(n_686),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_633),
.B(n_227),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_615),
.B(n_202),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_694),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_615),
.B(n_270),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_567),
.B(n_514),
.Y(n_814)
);

NAND3xp33_ASAP7_75t_L g815 ( 
.A(n_612),
.B(n_271),
.C(n_219),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_677),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_602),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_642),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_631),
.B(n_514),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_573),
.B(n_479),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_612),
.B(n_272),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_596),
.A2(n_227),
.B1(n_195),
.B2(n_212),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_621),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_667),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_613),
.Y(n_825)
);

OR2x2_ASAP7_75t_L g826 ( 
.A(n_640),
.B(n_203),
.Y(n_826)
);

INVx5_ASAP7_75t_L g827 ( 
.A(n_686),
.Y(n_827)
);

AND2x6_ASAP7_75t_SL g828 ( 
.A(n_661),
.B(n_195),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_573),
.B(n_479),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_554),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_621),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_617),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_621),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_697),
.A2(n_606),
.B1(n_625),
.B2(n_661),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_580),
.B(n_479),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_697),
.A2(n_195),
.B1(n_479),
.B2(n_463),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_666),
.B(n_0),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_675),
.B(n_103),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_677),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_681),
.B(n_108),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_591),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_561),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_627),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_672),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_685),
.B(n_463),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_628),
.B(n_1),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_660),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_563),
.A2(n_463),
.B(n_118),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_609),
.Y(n_849)
);

AND3x2_ASAP7_75t_SL g850 ( 
.A(n_650),
.B(n_2),
.C(n_5),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_698),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_590),
.B(n_2),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_564),
.B(n_117),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_578),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_650),
.B(n_5),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_583),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_783),
.A2(n_566),
.B(n_698),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_745),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_707),
.Y(n_859)
);

OAI21xp33_ASAP7_75t_L g860 ( 
.A1(n_810),
.A2(n_632),
.B(n_609),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_716),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_710),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_699),
.B(n_698),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_834),
.A2(n_687),
.B1(n_698),
.B2(n_656),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_817),
.B(n_692),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_R g866 ( 
.A(n_763),
.B(n_562),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_783),
.A2(n_664),
.B(n_659),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_788),
.A2(n_657),
.B(n_668),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_722),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_712),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_732),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.Y(n_871)
);

AO21x1_ASAP7_75t_L g872 ( 
.A1(n_703),
.A2(n_634),
.B(n_635),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_788),
.A2(n_669),
.B(n_695),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_722),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_732),
.A2(n_636),
.B(n_607),
.C(n_696),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_790),
.A2(n_690),
.B(n_665),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_787),
.B(n_607),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_825),
.B(n_752),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_768),
.B(n_684),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_728),
.B(n_652),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_708),
.B(n_645),
.Y(n_881)
);

BUFx8_ASAP7_75t_L g882 ( 
.A(n_757),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_702),
.B(n_651),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_790),
.A2(n_643),
.B(n_641),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_725),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_739),
.B(n_116),
.Y(n_886)
);

NOR2x1_ASAP7_75t_L g887 ( 
.A(n_745),
.B(n_102),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_779),
.A2(n_781),
.B1(n_717),
.B2(n_711),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_739),
.B(n_8),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_722),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_744),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_776),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_787),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_809),
.A2(n_98),
.B(n_94),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_721),
.B(n_16),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_721),
.B(n_18),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_SL g897 ( 
.A1(n_837),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_747),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_832),
.B(n_31),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_809),
.A2(n_49),
.B(n_57),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_741),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_708),
.B(n_59),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_734),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_708),
.B(n_32),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_734),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_718),
.A2(n_35),
.B(n_37),
.Y(n_906)
);

CKINVDCx16_ASAP7_75t_R g907 ( 
.A(n_753),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_816),
.B(n_839),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_724),
.A2(n_813),
.B(n_811),
.C(n_821),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_708),
.B(n_746),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_796),
.A2(n_726),
.B(n_849),
.C(n_841),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_826),
.B(n_700),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_809),
.A2(n_827),
.B(n_719),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_750),
.B(n_751),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_734),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_750),
.B(n_751),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_754),
.B(n_843),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_724),
.A2(n_730),
.B(n_754),
.C(n_723),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_770),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_786),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_793),
.B(n_818),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_793),
.B(n_818),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_708),
.B(n_797),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_827),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_827),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_704),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_827),
.A2(n_719),
.B(n_706),
.Y(n_927)
);

OR2x6_ASAP7_75t_SL g928 ( 
.A(n_815),
.B(n_713),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_740),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_723),
.B(n_743),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_799),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_824),
.Y(n_932)
);

OAI22x1_ASAP7_75t_L g933 ( 
.A1(n_852),
.A2(n_855),
.B1(n_850),
.B2(n_714),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_706),
.A2(n_769),
.B(n_766),
.Y(n_934)
);

BUFx8_ASAP7_75t_L g935 ( 
.A(n_844),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_766),
.A2(n_769),
.B(n_762),
.Y(n_936)
);

AND2x6_ASAP7_75t_L g937 ( 
.A(n_814),
.B(n_705),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_729),
.A2(n_761),
.B(n_758),
.C(n_756),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_736),
.B(n_807),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_796),
.A2(n_718),
.B(n_778),
.C(n_789),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_742),
.A2(n_803),
.B(n_778),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_847),
.B(n_755),
.Y(n_942)
);

OAI22x1_ASAP7_75t_L g943 ( 
.A1(n_850),
.A2(n_836),
.B1(n_736),
.B2(n_782),
.Y(n_943)
);

OAI21xp33_ASAP7_75t_L g944 ( 
.A1(n_822),
.A2(n_764),
.B(n_773),
.Y(n_944)
);

CKINVDCx10_ASAP7_75t_R g945 ( 
.A(n_707),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_707),
.B(n_846),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_846),
.A2(n_773),
.B(n_795),
.C(n_720),
.Y(n_947)
);

AO22x1_ASAP7_75t_L g948 ( 
.A1(n_838),
.A2(n_806),
.B1(n_840),
.B2(n_765),
.Y(n_948)
);

AO31x2_ASAP7_75t_L g949 ( 
.A1(n_735),
.A2(n_853),
.A3(n_848),
.B(n_808),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_819),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_737),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_737),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_814),
.A2(n_801),
.B1(n_731),
.B2(n_705),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_701),
.Y(n_954)
);

O2A1O1Ixp5_ASAP7_75t_L g955 ( 
.A1(n_853),
.A2(n_845),
.B(n_784),
.C(n_748),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_784),
.A2(n_803),
.B(n_835),
.Y(n_956)
);

NAND2x1_ASAP7_75t_L g957 ( 
.A(n_759),
.B(n_794),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_737),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_846),
.B(n_819),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_808),
.A2(n_715),
.B(n_835),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_709),
.B(n_733),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_805),
.A2(n_804),
.B(n_791),
.C(n_792),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_709),
.B(n_733),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_715),
.A2(n_801),
.B(n_771),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_760),
.Y(n_965)
);

AO31x2_ASAP7_75t_L g966 ( 
.A1(n_848),
.A2(n_777),
.A3(n_771),
.B(n_774),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_800),
.B(n_812),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_708),
.B(n_785),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_840),
.Y(n_969)
);

BUFx2_ASAP7_75t_SL g970 ( 
.A(n_738),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_806),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_798),
.B(n_765),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_774),
.A2(n_777),
.B(n_820),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_830),
.B(n_856),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_842),
.B(n_854),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_SL g976 ( 
.A(n_738),
.B(n_760),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_820),
.A2(n_829),
.B(n_738),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_760),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_759),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_772),
.B(n_780),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_861),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_878),
.B(n_828),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_917),
.B(n_765),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_973),
.A2(n_829),
.B(n_749),
.Y(n_984)
);

AOI221x1_ASAP7_75t_L g985 ( 
.A1(n_888),
.A2(n_838),
.B1(n_802),
.B2(n_833),
.C(n_831),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_921),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_863),
.A2(n_941),
.B(n_927),
.Y(n_987)
);

OAI21x1_ASAP7_75t_L g988 ( 
.A1(n_977),
.A2(n_802),
.B(n_833),
.Y(n_988)
);

AOI221x1_ASAP7_75t_L g989 ( 
.A1(n_944),
.A2(n_831),
.B1(n_823),
.B2(n_780),
.C(n_772),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_870),
.Y(n_990)
);

NAND2x1_ASAP7_75t_L g991 ( 
.A(n_924),
.B(n_794),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_867),
.A2(n_738),
.B(n_727),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_918),
.A2(n_767),
.B(n_775),
.Y(n_993)
);

O2A1O1Ixp5_ASAP7_75t_SL g994 ( 
.A1(n_904),
.A2(n_775),
.B(n_823),
.C(n_851),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_934),
.A2(n_851),
.B(n_806),
.Y(n_995)
);

NOR2x1_ASAP7_75t_L g996 ( 
.A(n_979),
.B(n_806),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_873),
.A2(n_936),
.B(n_868),
.Y(n_997)
);

INVx6_ASAP7_75t_L g998 ( 
.A(n_882),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_922),
.B(n_877),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_914),
.B(n_916),
.Y(n_1000)
);

O2A1O1Ixp5_ASAP7_75t_SL g1001 ( 
.A1(n_886),
.A2(n_902),
.B(n_923),
.C(n_910),
.Y(n_1001)
);

OR2x6_ASAP7_75t_L g1002 ( 
.A(n_892),
.B(n_932),
.Y(n_1002)
);

AND2x6_ASAP7_75t_SL g1003 ( 
.A(n_912),
.B(n_889),
.Y(n_1003)
);

AO21x1_ASAP7_75t_L g1004 ( 
.A1(n_947),
.A2(n_864),
.B(n_972),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_907),
.Y(n_1005)
);

CKINVDCx6p67_ASAP7_75t_R g1006 ( 
.A(n_945),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_901),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_895),
.Y(n_1008)
);

AOI21x1_ASAP7_75t_L g1009 ( 
.A1(n_960),
.A2(n_857),
.B(n_964),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_930),
.B(n_967),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_859),
.B(n_939),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_859),
.B(n_969),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_928),
.B(n_959),
.Y(n_1013)
);

AO31x2_ASAP7_75t_L g1014 ( 
.A1(n_940),
.A2(n_872),
.A3(n_911),
.B(n_962),
.Y(n_1014)
);

INVx8_ASAP7_75t_L g1015 ( 
.A(n_859),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_L g1016 ( 
.A(n_942),
.B(n_883),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_879),
.A2(n_884),
.B(n_881),
.Y(n_1017)
);

CKINVDCx14_ASAP7_75t_R g1018 ( 
.A(n_929),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_876),
.A2(n_860),
.B(n_955),
.Y(n_1019)
);

AO31x2_ASAP7_75t_L g1020 ( 
.A1(n_953),
.A2(n_943),
.A3(n_968),
.B(n_913),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_906),
.A2(n_875),
.B(n_963),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_938),
.A2(n_858),
.B(n_887),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_858),
.A2(n_887),
.B(n_957),
.Y(n_1023)
);

NAND2x1_ASAP7_75t_L g1024 ( 
.A(n_924),
.B(n_925),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_974),
.B(n_975),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_L g1026 ( 
.A(n_919),
.B(n_931),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_950),
.B(n_946),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_894),
.A2(n_900),
.B(n_980),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_948),
.A2(n_880),
.B(n_961),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_925),
.A2(n_956),
.B(n_961),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_871),
.A2(n_862),
.B(n_891),
.Y(n_1031)
);

NAND3x1_ASAP7_75t_L g1032 ( 
.A(n_896),
.B(n_899),
.C(n_897),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_866),
.B(n_885),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_956),
.A2(n_951),
.B(n_979),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_966),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_920),
.B(n_926),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_933),
.B(n_966),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_905),
.A2(n_937),
.B(n_966),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_905),
.A2(n_937),
.B(n_949),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_937),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_971),
.B(n_937),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_893),
.B(n_949),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_SL g1043 ( 
.A1(n_945),
.A2(n_935),
.B(n_954),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_949),
.A2(n_978),
.B(n_976),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_970),
.A2(n_978),
.B(n_874),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_869),
.A2(n_874),
.B(n_965),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_890),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_903),
.A2(n_915),
.B(n_952),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_915),
.B(n_952),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_915),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_958),
.B(n_965),
.Y(n_1051)
);

NAND3x1_ASAP7_75t_L g1052 ( 
.A(n_935),
.B(n_882),
.C(n_958),
.Y(n_1052)
);

AO31x2_ASAP7_75t_L g1053 ( 
.A1(n_940),
.A2(n_872),
.A3(n_699),
.B(n_888),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_909),
.A2(n_699),
.B(n_589),
.C(n_574),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_867),
.A2(n_934),
.B(n_873),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_878),
.B(n_328),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_878),
.B(n_917),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_859),
.Y(n_1058)
);

INVx3_ASAP7_75t_SL g1059 ( 
.A(n_929),
.Y(n_1059)
);

INVxp67_ASAP7_75t_SL g1060 ( 
.A(n_908),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_878),
.B(n_328),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_878),
.B(n_917),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_863),
.A2(n_703),
.B(n_941),
.Y(n_1063)
);

AO32x2_ASAP7_75t_L g1064 ( 
.A1(n_888),
.A2(n_864),
.A3(n_897),
.B1(n_953),
.B2(n_623),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_859),
.B(n_976),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_888),
.A2(n_699),
.B1(n_878),
.B2(n_865),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_861),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_SL g1068 ( 
.A1(n_888),
.A2(n_699),
.B(n_864),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_878),
.B(n_328),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_867),
.A2(n_934),
.B(n_873),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_861),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_R g1072 ( 
.A(n_866),
.B(n_458),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_878),
.B(n_328),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_909),
.A2(n_699),
.B(n_589),
.C(n_574),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_973),
.A2(n_977),
.B(n_857),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_940),
.A2(n_872),
.A3(n_699),
.B(n_888),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_973),
.A2(n_977),
.B(n_857),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_921),
.B(n_922),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_859),
.B(n_921),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_973),
.A2(n_977),
.B(n_857),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_912),
.A2(n_589),
.B1(n_574),
.B2(n_598),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_898),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_859),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_912),
.B(n_787),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_SL g1085 ( 
.A(n_897),
.B(n_488),
.C(n_422),
.Y(n_1085)
);

AO31x2_ASAP7_75t_L g1086 ( 
.A1(n_940),
.A2(n_872),
.A3(n_699),
.B(n_888),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_861),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_R g1088 ( 
.A(n_907),
.B(n_451),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_861),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_867),
.A2(n_934),
.B(n_873),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_861),
.Y(n_1091)
);

OA22x2_ASAP7_75t_L g1092 ( 
.A1(n_897),
.A2(n_810),
.B1(n_933),
.B2(n_478),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_861),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_888),
.A2(n_699),
.B1(n_878),
.B2(n_865),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_861),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_859),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_888),
.A2(n_699),
.B(n_589),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_924),
.Y(n_1098)
);

O2A1O1Ixp5_ASAP7_75t_L g1099 ( 
.A1(n_888),
.A2(n_699),
.B(n_574),
.C(n_589),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_929),
.Y(n_1100)
);

OAI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1081),
.A2(n_1092),
.B1(n_1025),
.B2(n_1097),
.Y(n_1101)
);

INVxp67_ASAP7_75t_SL g1102 ( 
.A(n_1060),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1099),
.A2(n_1074),
.B(n_1054),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_982),
.A2(n_1073),
.B1(n_1069),
.B2(n_1061),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_990),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_981),
.Y(n_1106)
);

OA21x2_ASAP7_75t_L g1107 ( 
.A1(n_985),
.A2(n_989),
.B(n_1019),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1015),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1083),
.B(n_1058),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_1004),
.A2(n_1017),
.A3(n_1090),
.B(n_1070),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_1083),
.B(n_1058),
.Y(n_1111)
);

AOI21x1_ASAP7_75t_L g1112 ( 
.A1(n_992),
.A2(n_995),
.B(n_1044),
.Y(n_1112)
);

NAND2x1p5_ASAP7_75t_L g1113 ( 
.A(n_1058),
.B(n_1096),
.Y(n_1113)
);

OAI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1010),
.A2(n_1008),
.B1(n_1062),
.B2(n_1057),
.Y(n_1114)
);

AO21x1_ASAP7_75t_L g1115 ( 
.A1(n_1066),
.A2(n_1094),
.B(n_1037),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_1007),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1079),
.B(n_1011),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1009),
.A2(n_987),
.B(n_1021),
.Y(n_1118)
);

INVx8_ASAP7_75t_L g1119 ( 
.A(n_1015),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1039),
.A2(n_997),
.B(n_1063),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1068),
.A2(n_1001),
.B(n_994),
.Y(n_1121)
);

CKINVDCx11_ASAP7_75t_R g1122 ( 
.A(n_1059),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1030),
.A2(n_1034),
.B(n_1055),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_993),
.A2(n_983),
.B(n_1031),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_986),
.B(n_999),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1038),
.A2(n_988),
.B(n_1028),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1078),
.B(n_1056),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_984),
.A2(n_1023),
.B(n_1022),
.Y(n_1128)
);

AO21x1_ASAP7_75t_L g1129 ( 
.A1(n_1042),
.A2(n_1040),
.B(n_1041),
.Y(n_1129)
);

BUFx5_ASAP7_75t_L g1130 ( 
.A(n_1040),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1016),
.B(n_1084),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1085),
.A2(n_1067),
.B1(n_1071),
.B2(n_1093),
.C(n_1087),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1029),
.A2(n_1035),
.B(n_1045),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1088),
.Y(n_1134)
);

AOI221xp5_ASAP7_75t_L g1135 ( 
.A1(n_1095),
.A2(n_1013),
.B1(n_1082),
.B2(n_1091),
.C(n_1089),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1032),
.A2(n_1072),
.B1(n_1036),
.B2(n_1027),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1002),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1035),
.A2(n_996),
.B(n_1048),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_1018),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1027),
.A2(n_1005),
.B1(n_1011),
.B2(n_1033),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1053),
.B(n_1076),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1064),
.A2(n_1026),
.B(n_1046),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1064),
.A2(n_1065),
.B(n_1051),
.Y(n_1143)
);

BUFx8_ASAP7_75t_SL g1144 ( 
.A(n_1100),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1064),
.A2(n_1050),
.B(n_1047),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1024),
.A2(n_991),
.B(n_1098),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1098),
.A2(n_1049),
.B(n_1047),
.Y(n_1147)
);

AOI211xp5_ASAP7_75t_L g1148 ( 
.A1(n_1003),
.A2(n_1043),
.B(n_1012),
.C(n_1096),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1012),
.A2(n_1002),
.B1(n_1096),
.B2(n_998),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1052),
.A2(n_998),
.B1(n_1006),
.B2(n_1053),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1020),
.B(n_1076),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1014),
.A2(n_1054),
.A3(n_1074),
.B(n_1004),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1020),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1020),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1086),
.A2(n_1077),
.B(n_1075),
.Y(n_1155)
);

OAI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1086),
.A2(n_1081),
.B1(n_1092),
.B2(n_1025),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1086),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_1068),
.B(n_948),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_990),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1058),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1083),
.Y(n_1161)
);

OAI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1081),
.A2(n_1092),
.B1(n_1025),
.B2(n_933),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1000),
.B(n_1010),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_981),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1075),
.A2(n_1080),
.B(n_1077),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1058),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_986),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1075),
.A2(n_1080),
.B(n_1077),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_985),
.A2(n_989),
.B(n_1019),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1025),
.A2(n_1081),
.B1(n_1010),
.B2(n_649),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_1015),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_990),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1000),
.B(n_1010),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1081),
.A2(n_574),
.B1(n_589),
.B2(n_598),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1088),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1054),
.A2(n_699),
.B(n_1074),
.C(n_1097),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_1100),
.Y(n_1177)
);

INVx6_ASAP7_75t_L g1178 ( 
.A(n_1015),
.Y(n_1178)
);

OA21x2_ASAP7_75t_L g1179 ( 
.A1(n_985),
.A2(n_989),
.B(n_1019),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1020),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1081),
.A2(n_574),
.B1(n_589),
.B2(n_598),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1000),
.B(n_1010),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1007),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_981),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1054),
.A2(n_699),
.B(n_1074),
.C(n_1097),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1020),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1055),
.A2(n_1090),
.B(n_1070),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1025),
.A2(n_1081),
.B1(n_1010),
.B2(n_649),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1099),
.A2(n_699),
.B(n_1054),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1054),
.A2(n_699),
.B(n_1074),
.C(n_1097),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_981),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1099),
.A2(n_699),
.B(n_1054),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_985),
.A2(n_989),
.B(n_1019),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_986),
.B(n_999),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_981),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1083),
.B(n_976),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1163),
.B(n_1173),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1174),
.A2(n_1181),
.B(n_1190),
.C(n_1185),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1187),
.A2(n_1185),
.B(n_1176),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1187),
.A2(n_1190),
.B(n_1176),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1194),
.B(n_1167),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1163),
.B(n_1173),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1105),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1180),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1159),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1182),
.B(n_1114),
.Y(n_1206)
);

O2A1O1Ixp5_ASAP7_75t_L g1207 ( 
.A1(n_1103),
.A2(n_1192),
.B(n_1189),
.C(n_1121),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1106),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1170),
.B(n_1188),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1170),
.B(n_1188),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1122),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1101),
.B(n_1162),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1102),
.B(n_1167),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1156),
.A2(n_1189),
.B1(n_1103),
.B2(n_1104),
.C(n_1115),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1116),
.B(n_1183),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1144),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1116),
.B(n_1183),
.Y(n_1217)
);

NOR2xp67_ASAP7_75t_L g1218 ( 
.A(n_1171),
.B(n_1108),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1136),
.A2(n_1140),
.B1(n_1135),
.B2(n_1149),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1135),
.B(n_1131),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1142),
.A2(n_1143),
.B(n_1121),
.C(n_1132),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1119),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1160),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_SL g1224 ( 
.A1(n_1186),
.A2(n_1129),
.B(n_1152),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1148),
.A2(n_1134),
.B1(n_1158),
.B2(n_1175),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1139),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_SL g1227 ( 
.A1(n_1150),
.A2(n_1158),
.B(n_1196),
.Y(n_1227)
);

OA21x2_ASAP7_75t_L g1228 ( 
.A1(n_1118),
.A2(n_1155),
.B(n_1120),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1172),
.Y(n_1229)
);

AOI211xp5_ASAP7_75t_L g1230 ( 
.A1(n_1150),
.A2(n_1142),
.B(n_1145),
.C(n_1143),
.Y(n_1230)
);

O2A1O1Ixp5_ASAP7_75t_L g1231 ( 
.A1(n_1112),
.A2(n_1124),
.B(n_1151),
.C(n_1153),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1160),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1147),
.B(n_1161),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1178),
.A2(n_1171),
.B1(n_1113),
.B2(n_1109),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1177),
.Y(n_1235)
);

AOI211xp5_ASAP7_75t_L g1236 ( 
.A1(n_1145),
.A2(n_1195),
.B(n_1191),
.C(n_1184),
.Y(n_1236)
);

O2A1O1Ixp5_ASAP7_75t_L g1237 ( 
.A1(n_1123),
.A2(n_1154),
.B(n_1157),
.C(n_1164),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1111),
.A2(n_1119),
.B1(n_1166),
.B2(n_1193),
.Y(n_1238)
);

AOI211xp5_ASAP7_75t_L g1239 ( 
.A1(n_1166),
.A2(n_1128),
.B(n_1138),
.C(n_1133),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1146),
.B(n_1126),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1107),
.A2(n_1179),
.B(n_1169),
.C(n_1110),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1130),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1130),
.B(n_1110),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1130),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1165),
.B(n_1168),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1174),
.A2(n_699),
.B(n_1074),
.C(n_1054),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1174),
.A2(n_888),
.B(n_1097),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1117),
.B(n_1137),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1117),
.B(n_1137),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1174),
.A2(n_1181),
.B1(n_1081),
.B2(n_1032),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1122),
.Y(n_1251)
);

O2A1O1Ixp5_ASAP7_75t_L g1252 ( 
.A1(n_1103),
.A2(n_1097),
.B(n_1099),
.C(n_1074),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1121),
.A2(n_997),
.B(n_1187),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1117),
.B(n_1137),
.Y(n_1254)
);

AOI21x1_ASAP7_75t_SL g1255 ( 
.A1(n_1141),
.A2(n_1042),
.B(n_1037),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1174),
.A2(n_1181),
.B1(n_1081),
.B2(n_1032),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1105),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1117),
.B(n_1137),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1127),
.B(n_1013),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1102),
.Y(n_1260)
);

AOI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1141),
.A2(n_1042),
.B(n_1037),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1163),
.B(n_1173),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1163),
.B(n_1173),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1122),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1174),
.A2(n_1097),
.B(n_1181),
.C(n_1081),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1125),
.B(n_1194),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1174),
.A2(n_888),
.B(n_1097),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1199),
.B(n_1200),
.Y(n_1268)
);

INVx5_ASAP7_75t_L g1269 ( 
.A(n_1240),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1265),
.A2(n_1267),
.B(n_1247),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1231),
.A2(n_1207),
.B(n_1221),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1209),
.B(n_1210),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1243),
.B(n_1230),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1237),
.Y(n_1274)
);

AO21x2_ASAP7_75t_L g1275 ( 
.A1(n_1221),
.A2(n_1241),
.B(n_1265),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1240),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1204),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1208),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1250),
.A2(n_1256),
.B1(n_1212),
.B2(n_1214),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1253),
.B(n_1231),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1198),
.A2(n_1246),
.B(n_1245),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1244),
.B(n_1207),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1246),
.A2(n_1212),
.B(n_1225),
.Y(n_1283)
);

AO21x2_ASAP7_75t_L g1284 ( 
.A1(n_1242),
.A2(n_1204),
.B(n_1244),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1227),
.B(n_1233),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1260),
.B(n_1206),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1228),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1228),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1213),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1197),
.B(n_1262),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1239),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1236),
.B(n_1252),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1201),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1252),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1220),
.A2(n_1224),
.B(n_1238),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1266),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1219),
.A2(n_1202),
.B(n_1263),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1215),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1255),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1259),
.B(n_1217),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1255),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1278),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1279),
.A2(n_1270),
.B1(n_1297),
.B2(n_1275),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1282),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1282),
.B(n_1254),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1284),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1282),
.B(n_1248),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1287),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_SL g1309 ( 
.A(n_1270),
.B(n_1234),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1289),
.B(n_1232),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1277),
.B(n_1223),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1278),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1269),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1284),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1269),
.Y(n_1315)
);

NOR2x1_ASAP7_75t_L g1316 ( 
.A(n_1291),
.B(n_1222),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1276),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1273),
.B(n_1249),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1277),
.Y(n_1319)
);

OR2x6_ASAP7_75t_L g1320 ( 
.A(n_1285),
.B(n_1258),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1269),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1274),
.B(n_1229),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1288),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1288),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1280),
.B(n_1261),
.Y(n_1325)
);

AOI221xp5_ASAP7_75t_L g1326 ( 
.A1(n_1303),
.A2(n_1279),
.B1(n_1283),
.B2(n_1292),
.C(n_1297),
.Y(n_1326)
);

OAI33xp33_ASAP7_75t_L g1327 ( 
.A1(n_1322),
.A2(n_1289),
.A3(n_1298),
.B1(n_1286),
.B2(n_1291),
.B3(n_1290),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1313),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1302),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1303),
.A2(n_1275),
.B1(n_1268),
.B2(n_1281),
.Y(n_1330)
);

AOI33xp33_ASAP7_75t_L g1331 ( 
.A1(n_1325),
.A2(n_1292),
.A3(n_1294),
.B1(n_1291),
.B2(n_1300),
.B3(n_1280),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1316),
.A2(n_1268),
.B1(n_1271),
.B2(n_1285),
.Y(n_1332)
);

AOI33xp33_ASAP7_75t_L g1333 ( 
.A1(n_1325),
.A2(n_1292),
.A3(n_1294),
.B1(n_1300),
.B2(n_1280),
.B3(n_1274),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1304),
.B(n_1293),
.Y(n_1334)
);

NOR5xp2_ASAP7_75t_SL g1335 ( 
.A(n_1309),
.B(n_1275),
.C(n_1295),
.D(n_1271),
.E(n_1281),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1308),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1313),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1309),
.A2(n_1268),
.B1(n_1285),
.B2(n_1272),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1302),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1318),
.A2(n_1275),
.B1(n_1268),
.B2(n_1281),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1302),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1313),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1308),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1316),
.A2(n_1268),
.B(n_1286),
.Y(n_1344)
);

NAND4xp25_ASAP7_75t_SL g1345 ( 
.A(n_1304),
.B(n_1272),
.C(n_1290),
.D(n_1294),
.Y(n_1345)
);

NOR4xp25_ASAP7_75t_SL g1346 ( 
.A(n_1317),
.B(n_1211),
.C(n_1264),
.D(n_1251),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1313),
.B(n_1269),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1308),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1322),
.Y(n_1349)
);

OAI221xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1325),
.A2(n_1268),
.B1(n_1272),
.B2(n_1298),
.C(n_1285),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1315),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1319),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1312),
.Y(n_1353)
);

OAI31xp33_ASAP7_75t_L g1354 ( 
.A1(n_1322),
.A2(n_1301),
.A3(n_1299),
.B(n_1296),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1311),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1318),
.A2(n_1275),
.B1(n_1268),
.B2(n_1281),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1315),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1320),
.Y(n_1358)
);

NOR2x1_ASAP7_75t_L g1359 ( 
.A(n_1345),
.B(n_1315),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1334),
.B(n_1319),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1332),
.B(n_1285),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1349),
.Y(n_1362)
);

INVx4_ASAP7_75t_SL g1363 ( 
.A(n_1332),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1344),
.A2(n_1306),
.B(n_1314),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1329),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1349),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1349),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1329),
.Y(n_1368)
);

NOR2x1p5_ASAP7_75t_L g1369 ( 
.A(n_1358),
.B(n_1315),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1334),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1347),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_SL g1372 ( 
.A(n_1335),
.B(n_1346),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1331),
.B(n_1296),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1339),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1337),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1337),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1336),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1339),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1358),
.B(n_1321),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1341),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1341),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_1355),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1337),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1355),
.B(n_1310),
.Y(n_1384)
);

INVx5_ASAP7_75t_L g1385 ( 
.A(n_1337),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1336),
.A2(n_1348),
.B(n_1343),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1333),
.B(n_1305),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1343),
.A2(n_1324),
.B(n_1323),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1327),
.B(n_1235),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1369),
.B(n_1337),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1369),
.B(n_1337),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1385),
.B(n_1351),
.Y(n_1392)
);

AND2x2_ASAP7_75t_SL g1393 ( 
.A(n_1389),
.B(n_1326),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1366),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1365),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1365),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1385),
.B(n_1351),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1373),
.B(n_1353),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1385),
.B(n_1351),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1385),
.B(n_1351),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1387),
.B(n_1352),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1368),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1385),
.B(n_1351),
.Y(n_1403)
);

NAND4xp25_ASAP7_75t_SL g1404 ( 
.A(n_1359),
.B(n_1330),
.C(n_1356),
.D(n_1340),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1366),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1370),
.B(n_1353),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1362),
.B(n_1384),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1368),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1385),
.B(n_1358),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1374),
.Y(n_1410)
);

NAND2x1_ASAP7_75t_L g1411 ( 
.A(n_1359),
.B(n_1383),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1374),
.Y(n_1412)
);

INVxp67_ASAP7_75t_SL g1413 ( 
.A(n_1367),
.Y(n_1413)
);

NAND4xp25_ASAP7_75t_L g1414 ( 
.A(n_1383),
.B(n_1354),
.C(n_1350),
.D(n_1310),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1371),
.B(n_1351),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_L g1416 ( 
.A(n_1383),
.B(n_1338),
.C(n_1358),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1371),
.B(n_1328),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1362),
.B(n_1352),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1371),
.B(n_1342),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1388),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_1376),
.Y(n_1421)
);

AOI211xp5_ASAP7_75t_L g1422 ( 
.A1(n_1372),
.A2(n_1354),
.B(n_1335),
.C(n_1226),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1384),
.B(n_1307),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1388),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1388),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1383),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1371),
.B(n_1342),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1378),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1360),
.B(n_1307),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1388),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1386),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1363),
.B(n_1347),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1422),
.B(n_1363),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1395),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1401),
.B(n_1360),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1395),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1390),
.B(n_1376),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1393),
.B(n_1382),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1396),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1411),
.B(n_1361),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1390),
.B(n_1363),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1401),
.B(n_1378),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1426),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1411),
.A2(n_1361),
.B1(n_1268),
.B2(n_1364),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1392),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1426),
.Y(n_1446)
);

NOR3x1_ASAP7_75t_L g1447 ( 
.A(n_1432),
.B(n_1414),
.C(n_1413),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1394),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1393),
.B(n_1375),
.Y(n_1449)
);

NAND2x1p5_ASAP7_75t_L g1450 ( 
.A(n_1392),
.B(n_1375),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1393),
.B(n_1293),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1391),
.B(n_1363),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1396),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1391),
.B(n_1415),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1415),
.B(n_1363),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1405),
.B(n_1346),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1398),
.B(n_1307),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1431),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1422),
.A2(n_1361),
.B1(n_1320),
.B2(n_1285),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1402),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1416),
.B(n_1379),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1398),
.B(n_1407),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1402),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1407),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1397),
.B(n_1379),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1408),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1431),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1449),
.B(n_1404),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1466),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1466),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1448),
.B(n_1421),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1433),
.A2(n_1361),
.B1(n_1421),
.B2(n_1409),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1443),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1450),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1454),
.B(n_1397),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1438),
.A2(n_1414),
.B(n_1364),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1459),
.A2(n_1361),
.B1(n_1409),
.B2(n_1403),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1450),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1441),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1454),
.B(n_1399),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1461),
.B(n_1216),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1450),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1451),
.B(n_1418),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1464),
.B(n_1418),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1443),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1441),
.B(n_1399),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1447),
.B(n_1423),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1434),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1445),
.B(n_1400),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1436),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1439),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1453),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1486),
.B(n_1452),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1476),
.A2(n_1456),
.B(n_1440),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_SL g1495 ( 
.A1(n_1468),
.A2(n_1445),
.B(n_1446),
.C(n_1444),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1468),
.B(n_1456),
.C(n_1446),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1474),
.Y(n_1497)
);

AOI222xp33_ASAP7_75t_L g1498 ( 
.A1(n_1487),
.A2(n_1452),
.B1(n_1455),
.B2(n_1437),
.C1(n_1465),
.C2(n_1460),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1481),
.B(n_1435),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1479),
.A2(n_1455),
.B1(n_1440),
.B2(n_1465),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1477),
.A2(n_1440),
.B1(n_1435),
.B2(n_1462),
.Y(n_1501)
);

OAI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1472),
.A2(n_1440),
.B1(n_1462),
.B2(n_1437),
.C(n_1442),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1480),
.A2(n_1457),
.B1(n_1409),
.B2(n_1442),
.Y(n_1503)
);

OAI221xp5_ASAP7_75t_L g1504 ( 
.A1(n_1484),
.A2(n_1471),
.B1(n_1481),
.B2(n_1483),
.C(n_1474),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_SL g1505 ( 
.A(n_1484),
.B(n_1403),
.C(n_1400),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1473),
.A2(n_1463),
.B(n_1467),
.C(n_1458),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1473),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1485),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1480),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1485),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1480),
.A2(n_1409),
.B1(n_1379),
.B2(n_1364),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1496),
.A2(n_1475),
.B1(n_1489),
.B2(n_1364),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1508),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1508),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1509),
.B(n_1489),
.Y(n_1515)
);

NAND2x1_ASAP7_75t_L g1516 ( 
.A(n_1493),
.B(n_1478),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1505),
.B(n_1499),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1504),
.B(n_1478),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1502),
.B(n_1482),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1507),
.B(n_1488),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1510),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1500),
.B(n_1482),
.Y(n_1522)
);

AND4x1_ASAP7_75t_L g1523 ( 
.A(n_1518),
.B(n_1498),
.C(n_1494),
.D(n_1506),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1513),
.B(n_1497),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_SL g1525 ( 
.A1(n_1519),
.A2(n_1501),
.B(n_1503),
.C(n_1511),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1517),
.A2(n_1495),
.B(n_1491),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1514),
.Y(n_1527)
);

NOR3xp33_ASAP7_75t_L g1528 ( 
.A(n_1522),
.B(n_1492),
.C(n_1490),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1512),
.B(n_1379),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1521),
.B(n_1469),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1515),
.B(n_1470),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1516),
.A2(n_1281),
.B1(n_1271),
.B2(n_1458),
.Y(n_1532)
);

OAI21xp33_ASAP7_75t_L g1533 ( 
.A1(n_1520),
.A2(n_1419),
.B(n_1417),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1526),
.A2(n_1467),
.B1(n_1431),
.B2(n_1419),
.C(n_1417),
.Y(n_1534)
);

AOI21xp33_ASAP7_75t_L g1535 ( 
.A1(n_1525),
.A2(n_1427),
.B(n_1408),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1528),
.A2(n_1271),
.B1(n_1427),
.B2(n_1295),
.Y(n_1536)
);

OAI21xp33_ASAP7_75t_L g1537 ( 
.A1(n_1533),
.A2(n_1428),
.B(n_1410),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1529),
.A2(n_1410),
.B1(n_1412),
.B2(n_1428),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1537),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1538),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1535),
.B(n_1524),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1534),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1536),
.B(n_1527),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1535),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1544),
.B(n_1523),
.Y(n_1545)
);

NOR3x1_ASAP7_75t_L g1546 ( 
.A(n_1541),
.B(n_1530),
.C(n_1531),
.Y(n_1546)
);

AOI211xp5_ASAP7_75t_L g1547 ( 
.A1(n_1544),
.A2(n_1218),
.B(n_1205),
.C(n_1203),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1542),
.B(n_1532),
.Y(n_1548)
);

OAI221xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1539),
.A2(n_1430),
.B1(n_1425),
.B2(n_1424),
.C(n_1420),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1546),
.B(n_1540),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1545),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1548),
.B(n_1543),
.Y(n_1552)
);

NOR2x1_ASAP7_75t_L g1553 ( 
.A(n_1550),
.B(n_1257),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1553),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1554),
.A2(n_1547),
.B1(n_1552),
.B2(n_1551),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1555),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_L g1557 ( 
.A(n_1556),
.B(n_1549),
.C(n_1412),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1557),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1557),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1558),
.A2(n_1559),
.B(n_1430),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1558),
.B(n_1406),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_R g1562 ( 
.A1(n_1560),
.A2(n_1561),
.B1(n_1430),
.B2(n_1420),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1562),
.A2(n_1425),
.B(n_1424),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1563),
.A2(n_1372),
.B1(n_1377),
.B2(n_1380),
.C(n_1381),
.Y(n_1564)
);

AOI211xp5_ASAP7_75t_L g1565 ( 
.A1(n_1564),
.A2(n_1429),
.B(n_1357),
.C(n_1377),
.Y(n_1565)
);


endmodule