module fake_aes_11993_n_28 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
NAND2xp5_ASAP7_75t_L g13 ( .A(n_1), .B(n_11), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_7), .A2(n_6), .B(n_3), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_8), .Y(n_15) );
INVx6_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_5), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_18), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
NOR2xp33_ASAP7_75t_SL g23 ( .A(n_22), .B(n_17), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_0), .Y(n_25) );
CKINVDCx6p67_ASAP7_75t_R g26 ( .A(n_25), .Y(n_26) );
OAI222xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_18), .B1(n_15), .B2(n_13), .C1(n_14), .C2(n_16), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_10), .B1(n_2), .B2(n_4), .Y(n_28) );
endmodule