module fake_netlist_5_1613_n_1945 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1945);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1945;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_43),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_61),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_133),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_81),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_23),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_35),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_101),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_0),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_165),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_102),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_83),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_13),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_117),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_60),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_147),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_124),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_169),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_9),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_19),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

INVx4_ASAP7_75t_R g231 ( 
.A(n_176),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_24),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_130),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_38),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_108),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_120),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_70),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_173),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_23),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_40),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_87),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_92),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_172),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_24),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_116),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_17),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_34),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_42),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_145),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_84),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_78),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_180),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_8),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_32),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_107),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_98),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_16),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_36),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_3),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_13),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_22),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_112),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_76),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_154),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_86),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_189),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_106),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_156),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_51),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_64),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_136),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_90),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_46),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_31),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_29),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_44),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_161),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_77),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_44),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_65),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_2),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_5),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_75),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_174),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_170),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_96),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_16),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_60),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_140),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_159),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_155),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_146),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_41),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_9),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_192),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_148),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_141),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_190),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_95),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_18),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_21),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_62),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_162),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_144),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_183),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_91),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_182),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_7),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_33),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_137),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_185),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_37),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_71),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_62),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_43),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_68),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_82),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_34),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_51),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_171),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_55),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_47),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_25),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_73),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_50),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_14),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_168),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_160),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_127),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_166),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_50),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_157),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_30),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_45),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_63),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_15),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_111),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_123),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_47),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_69),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_94),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_21),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_167),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_20),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_61),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_163),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_29),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_55),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_20),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_26),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_104),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_5),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_39),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_132),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_115),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_109),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_8),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_66),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_135),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_178),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_125),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_31),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_67),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_179),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_72),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_110),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_122),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_138),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_18),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_114),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_74),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_15),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_59),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_88),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_12),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_80),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_32),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_26),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_121),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_181),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_150),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_6),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_58),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_1),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_177),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_184),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_199),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_387),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_232),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_199),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_297),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_200),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_284),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_199),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_199),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_235),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_199),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_258),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_239),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_394),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_258),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_258),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_258),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_244),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_240),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_258),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_287),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_254),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_255),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_287),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_302),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_287),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_287),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_256),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_287),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_368),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_213),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_368),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_257),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_262),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_238),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_368),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_197),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g439 ( 
.A(n_195),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_197),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_268),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_268),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_310),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_310),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_195),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_201),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_269),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_282),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_271),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_273),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_276),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_282),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_333),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_280),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_333),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_305),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_356),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_206),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_285),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_356),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_323),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_353),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_247),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_212),
.B(n_0),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_226),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_324),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_385),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_353),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g469 ( 
.A(n_207),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_324),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_292),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_234),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_243),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_201),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_241),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_249),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_263),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_251),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_265),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_248),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_283),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_303),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_294),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_302),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_295),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_304),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_296),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_299),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_211),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_311),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_300),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_301),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_315),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_319),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_322),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_325),
.Y(n_497)
);

BUFx2_ASAP7_75t_SL g498 ( 
.A(n_212),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_336),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_211),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_419),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_419),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_398),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_400),
.B(n_216),
.Y(n_506)
);

BUFx8_ASAP7_75t_L g507 ( 
.A(n_424),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_405),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_404),
.A2(n_415),
.B1(n_411),
.B2(n_399),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_405),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_406),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_407),
.B(n_216),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_422),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_410),
.B(n_272),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_409),
.B(n_202),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_412),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_416),
.B(n_272),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_498),
.B(n_308),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_412),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_445),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_414),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_418),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_423),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_423),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_498),
.B(n_308),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_420),
.B(n_348),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_446),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g538 ( 
.A1(n_425),
.A2(n_229),
.B(n_198),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_481),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_428),
.B(n_348),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_494),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_421),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_427),
.B(n_365),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_433),
.B(n_365),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_429),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_429),
.B(n_370),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_431),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_435),
.B(n_370),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_403),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_430),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_475),
.A2(n_359),
.B1(n_252),
.B2(n_395),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_434),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_478),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_437),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_474),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_473),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_490),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_464),
.B(n_202),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_447),
.B(n_198),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_449),
.B(n_229),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_473),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_450),
.B(n_250),
.Y(n_574)
);

CKINVDCx11_ASAP7_75t_R g575 ( 
.A(n_456),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_461),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_451),
.B(n_454),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_462),
.B(n_278),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_471),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_484),
.B(n_486),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_476),
.B(n_202),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_467),
.Y(n_582)
);

AO22x2_ASAP7_75t_L g583 ( 
.A1(n_511),
.A2(n_278),
.B1(n_286),
.B2(n_279),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_505),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_502),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_505),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_556),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_532),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_493),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_524),
.B(n_488),
.Y(n_591)
);

AO21x2_ASAP7_75t_L g592 ( 
.A1(n_571),
.A2(n_203),
.B(n_196),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_502),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_506),
.B(n_489),
.Y(n_594)
);

INVxp33_ASAP7_75t_SL g595 ( 
.A(n_562),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_532),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_567),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_504),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_535),
.B(n_492),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_544),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_504),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_528),
.A2(n_331),
.B1(n_380),
.B2(n_236),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_559),
.B(n_328),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_L g604 ( 
.A(n_537),
.B(n_463),
.C(n_436),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_570),
.A2(n_465),
.B1(n_439),
.B2(n_373),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_L g607 ( 
.A(n_570),
.B(n_202),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_509),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_574),
.B(n_424),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_508),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_532),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_504),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_512),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_512),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_501),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_504),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_501),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_501),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_513),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_578),
.B(n_462),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_515),
.B(n_459),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_520),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_513),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_517),
.Y(n_624)
);

AND3x2_ASAP7_75t_L g625 ( 
.A(n_555),
.B(n_286),
.C(n_279),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_572),
.B(n_485),
.Y(n_626)
);

AND3x2_ASAP7_75t_L g627 ( 
.A(n_569),
.B(n_313),
.C(n_293),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_570),
.A2(n_383),
.B1(n_393),
.B2(n_345),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_518),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_504),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_577),
.B(n_443),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_545),
.B(n_485),
.Y(n_632)
);

XOR2x2_ASAP7_75t_L g633 ( 
.A(n_541),
.B(n_500),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_514),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_580),
.A2(n_417),
.B1(n_466),
.B2(n_470),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_578),
.B(n_468),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_514),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_519),
.B(n_293),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_557),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_518),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_523),
.B(n_458),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_514),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_564),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_536),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_546),
.B(n_547),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_545),
.B(n_302),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_564),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_514),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_516),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_514),
.Y(n_651)
);

INVx8_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_521),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_540),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_521),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_570),
.B(n_202),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_579),
.B(n_340),
.Y(n_657)
);

AND3x2_ASAP7_75t_L g658 ( 
.A(n_541),
.B(n_367),
.C(n_313),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_544),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_525),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_570),
.B(n_306),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_578),
.B(n_468),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_525),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_522),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_579),
.B(n_340),
.Y(n_665)
);

INVx8_ASAP7_75t_L g666 ( 
.A(n_570),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_527),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_507),
.B(n_444),
.C(n_578),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_565),
.B(n_469),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_522),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_565),
.B(n_482),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_527),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_526),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_507),
.B(n_253),
.C(n_245),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_529),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_549),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_549),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_540),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_526),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_552),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_543),
.B(n_438),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_552),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_503),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_543),
.B(n_317),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_507),
.B(n_340),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_575),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_543),
.B(n_344),
.Y(n_688)
);

NAND3xp33_ASAP7_75t_SL g689 ( 
.A(n_576),
.B(n_388),
.C(n_218),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_543),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_540),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_568),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_550),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_550),
.B(n_440),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_550),
.B(n_320),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_507),
.B(n_204),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_550),
.B(n_530),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_530),
.B(n_338),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_568),
.B(n_204),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_540),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_503),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_540),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_548),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_503),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_573),
.B(n_205),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_539),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_573),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_548),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_581),
.B(n_205),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_581),
.B(n_208),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_531),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_548),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_531),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_520),
.B(n_306),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_533),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_533),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_534),
.B(n_339),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_539),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_534),
.B(n_208),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_581),
.B(n_209),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_548),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_542),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_542),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_520),
.B(n_306),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_551),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

NOR2x1p5_ASAP7_75t_L g728 ( 
.A(n_566),
.B(n_215),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_553),
.B(n_264),
.C(n_260),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_553),
.A2(n_222),
.B1(n_397),
.B2(n_396),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_566),
.B(n_476),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_548),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_560),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_566),
.B(n_209),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_560),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_584),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_585),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_690),
.B(n_510),
.Y(n_738)
);

BUFx6f_ASAP7_75t_SL g739 ( 
.A(n_597),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_639),
.A2(n_538),
.B1(n_367),
.B2(n_306),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_690),
.B(n_510),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_723),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_585),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_639),
.B(n_306),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

O2A1O1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_734),
.A2(n_477),
.B(n_479),
.C(n_480),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_642),
.B(n_510),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_624),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_589),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_645),
.B(n_214),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_594),
.B(n_510),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_693),
.B(n_554),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_646),
.A2(n_357),
.B1(n_354),
.B2(n_351),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_693),
.B(n_554),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_593),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_591),
.B(n_554),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_646),
.A2(n_346),
.B1(n_343),
.B2(n_341),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_589),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_596),
.B(n_214),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_599),
.B(n_554),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_669),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_626),
.B(n_217),
.Y(n_762)
);

INVx8_ASAP7_75t_L g763 ( 
.A(n_631),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_609),
.B(n_217),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_593),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_586),
.B(n_558),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_646),
.A2(n_369),
.B1(n_222),
.B2(n_221),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_588),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_644),
.B(n_558),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_651),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_646),
.B(n_220),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_595),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_631),
.B(n_220),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_648),
.B(n_692),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_684),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_583),
.A2(n_538),
.B1(n_334),
.B2(n_330),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_707),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_731),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_712),
.B(n_558),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_731),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_714),
.B(n_558),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_221),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_731),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_716),
.B(n_558),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_596),
.B(n_611),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_638),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_717),
.B(n_561),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_622),
.B(n_538),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_596),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_728),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_635),
.B(n_362),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_596),
.B(n_210),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_583),
.A2(n_592),
.B1(n_628),
.B2(n_682),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_596),
.B(n_223),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_638),
.B(n_561),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_671),
.B(n_267),
.C(n_266),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_631),
.B(n_362),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_650),
.B(n_561),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_583),
.A2(n_538),
.B1(n_327),
.B2(n_326),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_650),
.B(n_561),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_597),
.B(n_358),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_624),
.B(n_358),
.Y(n_802)
);

AO221x1_ASAP7_75t_L g803 ( 
.A1(n_583),
.A2(n_230),
.B1(n_366),
.B2(n_225),
.C(n_352),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_653),
.B(n_561),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_653),
.B(n_563),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_686),
.B(n_477),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_655),
.B(n_563),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_655),
.B(n_563),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_701),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_651),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_699),
.B(n_281),
.C(n_270),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_620),
.B(n_358),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_664),
.B(n_563),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_664),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_611),
.B(n_227),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_670),
.B(n_673),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_611),
.B(n_233),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_670),
.B(n_563),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_620),
.B(n_479),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_673),
.B(n_237),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_647),
.B(n_369),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_657),
.B(n_371),
.Y(n_822)
);

NOR3xp33_ASAP7_75t_L g823 ( 
.A(n_689),
.B(n_480),
.C(n_499),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_595),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_680),
.B(n_242),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_680),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_723),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_735),
.B(n_246),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_735),
.B(n_259),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_724),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_611),
.Y(n_831)
);

NOR2x1p5_ASAP7_75t_L g832 ( 
.A(n_674),
.B(n_215),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_615),
.B(n_261),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_611),
.B(n_371),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_636),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_701),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_636),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_640),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_615),
.B(n_274),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_662),
.B(n_483),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_662),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_617),
.B(n_275),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_682),
.Y(n_843)
);

CKINVDCx11_ASAP7_75t_R g844 ( 
.A(n_640),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_697),
.B(n_288),
.Y(n_845)
);

NAND2x1_ASAP7_75t_L g846 ( 
.A(n_601),
.B(n_520),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_617),
.B(n_307),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_SL g848 ( 
.A(n_600),
.B(n_582),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_704),
.Y(n_849)
);

INVx5_ASAP7_75t_L g850 ( 
.A(n_652),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_592),
.A2(n_321),
.B1(n_349),
.B2(n_316),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_618),
.B(n_592),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_704),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_706),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_694),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_618),
.B(n_698),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_658),
.Y(n_857)
);

INVxp33_ASAP7_75t_L g858 ( 
.A(n_633),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_606),
.B(n_309),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_706),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_708),
.B(n_314),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_708),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_694),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_665),
.B(n_372),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_610),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_718),
.B(n_381),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_705),
.B(n_382),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_724),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_652),
.B(n_372),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_719),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_719),
.B(n_374),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_720),
.B(n_520),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_621),
.B(n_520),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_726),
.B(n_520),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_652),
.B(n_374),
.Y(n_875)
);

BUFx8_ASAP7_75t_L g876 ( 
.A(n_687),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_633),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_632),
.B(n_375),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_668),
.B(n_483),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_688),
.A2(n_607),
.B1(n_656),
.B2(n_661),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_605),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_726),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_729),
.B(n_730),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_605),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_608),
.Y(n_885)
);

BUFx6f_ASAP7_75t_SL g886 ( 
.A(n_687),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_727),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_622),
.B(n_727),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_733),
.B(n_375),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_SL g890 ( 
.A(n_696),
.B(n_218),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_685),
.B(n_376),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_695),
.B(n_376),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_651),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_733),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_608),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_602),
.B(n_499),
.C(n_497),
.Y(n_896)
);

NAND2xp33_ASAP7_75t_L g897 ( 
.A(n_652),
.B(n_377),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_613),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_625),
.B(n_487),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_613),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_598),
.B(n_377),
.Y(n_901)
);

BUFx6f_ASAP7_75t_SL g902 ( 
.A(n_587),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_SL g903 ( 
.A1(n_603),
.A2(n_219),
.B1(n_224),
.B2(n_228),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_598),
.B(n_378),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_622),
.B(n_378),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_688),
.B(n_379),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_598),
.B(n_379),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_856),
.B(n_614),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_761),
.B(n_614),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_747),
.B(n_619),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_850),
.A2(n_666),
.B(n_616),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_742),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_838),
.B(n_600),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_744),
.A2(n_710),
.B1(n_711),
.B2(n_721),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_748),
.Y(n_915)
);

AND2x6_ASAP7_75t_SL g916 ( 
.A(n_821),
.B(n_603),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_SL g917 ( 
.A(n_858),
.B(n_659),
.C(n_821),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_742),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_898),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_816),
.B(n_619),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_883),
.B(n_659),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_898),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_827),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_750),
.B(n_590),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_827),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_786),
.B(n_623),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_830),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_893),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_814),
.B(n_826),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_SL g930 ( 
.A1(n_740),
.A2(n_666),
.B(n_491),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_R g931 ( 
.A(n_865),
.B(n_627),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_843),
.A2(n_604),
.B1(n_722),
.B2(n_630),
.Y(n_932)
);

OAI221xp5_ASAP7_75t_L g933 ( 
.A1(n_906),
.A2(n_590),
.B1(n_312),
.B2(n_298),
.C(n_291),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_789),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_801),
.B(n_487),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_778),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_772),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_780),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_762),
.B(n_612),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_783),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_868),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_772),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_855),
.A2(n_863),
.B1(n_837),
.B2(n_841),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_750),
.B(n_491),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_762),
.B(n_612),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_867),
.B(n_612),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_891),
.B(n_630),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_850),
.B(n_622),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_882),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_751),
.B(n_623),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_891),
.B(n_892),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_892),
.B(n_630),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_789),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_849),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_835),
.B(n_495),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_852),
.B(n_629),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_777),
.B(n_740),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_774),
.B(n_634),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_824),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_845),
.A2(n_722),
.B1(n_637),
.B2(n_732),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_802),
.B(n_495),
.Y(n_961)
);

AND2x2_ASAP7_75t_SL g962 ( 
.A(n_848),
.B(n_607),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_840),
.B(n_634),
.Y(n_963)
);

INVx6_ASAP7_75t_L g964 ( 
.A(n_876),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_824),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_736),
.B(n_634),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_745),
.B(n_637),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_789),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_877),
.B(n_496),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_849),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_749),
.B(n_637),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_SL g972 ( 
.A1(n_903),
.A2(n_666),
.B1(n_656),
.B2(n_661),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_887),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_850),
.B(n_622),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_758),
.B(n_643),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_859),
.A2(n_672),
.B(n_663),
.C(n_667),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_775),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_763),
.B(n_790),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_819),
.Y(n_979)
);

BUFx4f_ASAP7_75t_SL g980 ( 
.A(n_876),
.Y(n_980)
);

NAND2xp33_ASAP7_75t_SL g981 ( 
.A(n_739),
.B(n_390),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_894),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_756),
.B(n_760),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_SL g984 ( 
.A(n_858),
.B(n_219),
.C(n_224),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_866),
.B(n_629),
.Y(n_985)
);

AND2x6_ASAP7_75t_L g986 ( 
.A(n_812),
.B(n_641),
.Y(n_986)
);

OR2x4_ASAP7_75t_L g987 ( 
.A(n_773),
.B(n_496),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_819),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_768),
.B(n_497),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_895),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_859),
.A2(n_676),
.B(n_660),
.C(n_663),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_850),
.B(n_666),
.Y(n_992)
);

INVx5_ASAP7_75t_L g993 ( 
.A(n_893),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_793),
.B(n_641),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_789),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_744),
.A2(n_675),
.B1(n_660),
.B2(n_667),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_878),
.B(n_764),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_809),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_793),
.B(n_836),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_853),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_854),
.B(n_672),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_851),
.A2(n_803),
.B1(n_906),
.B2(n_845),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_860),
.B(n_675),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_822),
.B(n_440),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_739),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_862),
.Y(n_1006)
);

AND2x6_ASAP7_75t_SL g1007 ( 
.A(n_822),
.B(n_441),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_870),
.B(n_676),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_878),
.B(n_390),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_857),
.B(n_879),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_737),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_851),
.B(n_677),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_844),
.B(n_902),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_890),
.B(n_389),
.C(n_386),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_743),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_881),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_773),
.B(n_601),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_785),
.A2(n_616),
.B(n_601),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_755),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_776),
.B(n_799),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_771),
.A2(n_732),
.B1(n_643),
.B2(n_649),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_785),
.A2(n_616),
.B(n_702),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_765),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_771),
.Y(n_1024)
);

NOR2x2_ASAP7_75t_L g1025 ( 
.A(n_806),
.B(n_228),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_864),
.B(n_782),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_764),
.B(n_782),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_776),
.B(n_677),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_902),
.Y(n_1029)
);

AND3x2_ASAP7_75t_SL g1030 ( 
.A(n_864),
.B(n_832),
.C(n_767),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_799),
.B(n_678),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_884),
.B(n_678),
.Y(n_1032)
);

NOR2x1_ASAP7_75t_L g1033 ( 
.A(n_806),
.B(n_796),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_885),
.Y(n_1034)
);

BUFx5_ASAP7_75t_L g1035 ( 
.A(n_788),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_797),
.A2(n_681),
.B(n_683),
.C(n_649),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_900),
.B(n_820),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_795),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_797),
.A2(n_732),
.B1(n_643),
.B2(n_649),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_825),
.B(n_681),
.Y(n_1040)
);

NOR2x1p5_ASAP7_75t_L g1041 ( 
.A(n_899),
.B(n_364),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_831),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_798),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_886),
.B(n_391),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_871),
.B(n_364),
.Y(n_1045)
);

INVx6_ASAP7_75t_L g1046 ( 
.A(n_899),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_828),
.B(n_683),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_879),
.B(n_654),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_871),
.A2(n_703),
.B1(n_654),
.B2(n_679),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_831),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_879),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_752),
.A2(n_702),
.B(n_651),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_SL g1053 ( 
.A(n_811),
.B(n_389),
.C(n_386),
.Y(n_1053)
);

CKINVDCx8_ASAP7_75t_R g1054 ( 
.A(n_763),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_SL g1055 ( 
.A(n_880),
.B(n_391),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_753),
.B(n_392),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_800),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_804),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_805),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_831),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_757),
.B(n_392),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_766),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_807),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_893),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_808),
.Y(n_1065)
);

CKINVDCx11_ASAP7_75t_R g1066 ( 
.A(n_763),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_806),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_813),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_833),
.A2(n_839),
.B1(n_842),
.B2(n_847),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_886),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_R g1071 ( 
.A(n_889),
.B(n_384),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_791),
.B(n_396),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_L g1073 ( 
.A(n_893),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_829),
.B(n_654),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_873),
.A2(n_703),
.B1(n_679),
.B2(n_702),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_823),
.B(n_679),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_818),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_901),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_880),
.B(n_904),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_907),
.B(n_397),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_788),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_754),
.A2(n_651),
.B(n_691),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_769),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_738),
.B(n_289),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_896),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_861),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_846),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_861),
.A2(n_703),
.B1(n_713),
.B2(n_709),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_779),
.Y(n_1089)
);

INVx5_ASAP7_75t_L g1090 ( 
.A(n_770),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_741),
.B(n_691),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_792),
.A2(n_713),
.B1(n_709),
.B2(n_700),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_810),
.B(n_691),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_888),
.B(n_441),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_874),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_SL g1096 ( 
.A1(n_872),
.A2(n_384),
.B1(n_355),
.B2(n_318),
.Y(n_1096)
);

AOI21xp33_ASAP7_75t_L g1097 ( 
.A1(n_781),
.A2(n_725),
.B(n_715),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_784),
.B(n_691),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1026),
.B(n_787),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_928),
.Y(n_1100)
);

NOR2x1_ASAP7_75t_L g1101 ( 
.A(n_997),
.B(n_905),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_951),
.B(n_905),
.Y(n_1102)
);

O2A1O1Ixp5_ASAP7_75t_L g1103 ( 
.A1(n_1027),
.A2(n_815),
.B(n_792),
.C(n_794),
.Y(n_1103)
);

AO31x2_ASAP7_75t_L g1104 ( 
.A1(n_1036),
.A2(n_455),
.A3(n_457),
.B(n_460),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_915),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_912),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_919),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1024),
.B(n_746),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_913),
.Y(n_1109)
);

CKINVDCx8_ASAP7_75t_R g1110 ( 
.A(n_1007),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_924),
.B(n_888),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1020),
.A2(n_794),
.B1(n_815),
.B2(n_817),
.Y(n_1112)
);

CKINVDCx16_ASAP7_75t_R g1113 ( 
.A(n_1013),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1020),
.A2(n_817),
.B1(n_290),
.B2(n_329),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_L g1115 ( 
.A1(n_1079),
.A2(n_448),
.B(n_457),
.C(n_455),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_961),
.B(n_442),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_933),
.B(n_759),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_957),
.A2(n_1002),
.B1(n_994),
.B2(n_1028),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_922),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_942),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1073),
.A2(n_897),
.B(n_875),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1073),
.A2(n_869),
.B(n_834),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_935),
.B(n_442),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_SL g1124 ( 
.A(n_917),
.B(n_350),
.C(n_332),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_930),
.A2(n_725),
.B(n_715),
.C(n_335),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_983),
.A2(n_448),
.B(n_452),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_944),
.B(n_691),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_928),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_962),
.B(n_700),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_993),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_909),
.B(n_700),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_994),
.A2(n_361),
.B1(n_337),
.B2(n_342),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_928),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_918),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1009),
.A2(n_452),
.B(n_453),
.C(n_460),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_983),
.A2(n_993),
.B(n_950),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_937),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_923),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1028),
.A2(n_360),
.B1(n_347),
.B2(n_453),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1055),
.A2(n_713),
.B(n_709),
.C(n_700),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_959),
.B(n_713),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_925),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_SL g1143 ( 
.A1(n_1017),
.A2(n_231),
.B(n_709),
.C(n_700),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_927),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1031),
.A2(n_709),
.B1(n_6),
.B2(n_7),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_1066),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_993),
.A2(n_194),
.B(n_164),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1012),
.A2(n_158),
.B(n_149),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_969),
.B(n_4),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1029),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_965),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_993),
.A2(n_142),
.B(n_139),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_926),
.Y(n_1153)
);

OR2x2_ASAP7_75t_L g1154 ( 
.A(n_1045),
.B(n_4),
.Y(n_1154)
);

AOI222xp33_ASAP7_75t_L g1155 ( 
.A1(n_984),
.A2(n_1096),
.B1(n_1051),
.B2(n_1085),
.C1(n_1004),
.C2(n_955),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_936),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_938),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1093),
.A2(n_129),
.B(n_128),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1010),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_908),
.B(n_126),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1010),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_987),
.B(n_10),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_987),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_908),
.B(n_119),
.Y(n_1164)
);

BUFx8_ASAP7_75t_L g1165 ( 
.A(n_1067),
.Y(n_1165)
);

XOR2x2_ASAP7_75t_L g1166 ( 
.A(n_921),
.B(n_11),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_910),
.A2(n_118),
.B(n_103),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_SL g1168 ( 
.A(n_1054),
.B(n_100),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1070),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1056),
.A2(n_11),
.B(n_12),
.C(n_19),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1061),
.A2(n_22),
.B(n_25),
.C(n_27),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1046),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1046),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1084),
.A2(n_27),
.B(n_28),
.C(n_30),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_1005),
.B(n_932),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_1064),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1038),
.B(n_1043),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1091),
.A2(n_920),
.B(n_947),
.Y(n_1178)
);

OAI22x1_ASAP7_75t_L g1179 ( 
.A1(n_943),
.A2(n_28),
.B1(n_33),
.B2(n_35),
.Y(n_1179)
);

BUFx2_ASAP7_75t_SL g1180 ( 
.A(n_979),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_952),
.A2(n_59),
.B(n_39),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_1071),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_926),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1057),
.B(n_37),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_988),
.B(n_40),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_939),
.A2(n_41),
.B(n_45),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_978),
.B(n_1048),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_SL g1188 ( 
.A(n_1090),
.B(n_964),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1031),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1189)
);

NOR2x1_ASAP7_75t_L g1190 ( 
.A(n_1033),
.B(n_978),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_955),
.B(n_49),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_929),
.B(n_52),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1089),
.B(n_52),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_986),
.A2(n_58),
.B1(n_54),
.B2(n_56),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_940),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_914),
.A2(n_53),
.B(n_54),
.C(n_56),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1076),
.B(n_53),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_999),
.A2(n_57),
.B1(n_1012),
.B2(n_972),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1048),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_911),
.A2(n_57),
.B(n_963),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_945),
.A2(n_985),
.B(n_1098),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_L g1202 ( 
.A1(n_1080),
.A2(n_946),
.B(n_985),
.C(n_1082),
.Y(n_1202)
);

OR2x6_ASAP7_75t_L g1203 ( 
.A(n_964),
.B(n_978),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1076),
.B(n_989),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_989),
.B(n_1086),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_986),
.A2(n_1094),
.B1(n_1083),
.B2(n_1068),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_980),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1044),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1098),
.A2(n_1074),
.B(n_992),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_990),
.Y(n_1211)
);

NAND2xp33_ASAP7_75t_SL g1212 ( 
.A(n_1053),
.B(n_1014),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1011),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_931),
.A2(n_999),
.B1(n_973),
.B2(n_941),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1072),
.A2(n_982),
.B(n_949),
.C(n_1037),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_L g1216 ( 
.A1(n_1069),
.A2(n_1063),
.B(n_1037),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1041),
.B(n_1094),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1042),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_976),
.A2(n_991),
.B(n_1077),
.C(n_1065),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1074),
.A2(n_1052),
.B(n_958),
.Y(n_1220)
);

CKINVDCx14_ASAP7_75t_R g1221 ( 
.A(n_981),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_916),
.B(n_1062),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1015),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_977),
.B(n_1000),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_998),
.Y(n_1225)
);

OA21x2_ASAP7_75t_L g1226 ( 
.A1(n_1040),
.A2(n_1047),
.B(n_996),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1050),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1019),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1040),
.B(n_1047),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1018),
.A2(n_1022),
.B(n_934),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_948),
.A2(n_974),
.B(n_1090),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_953),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_986),
.A2(n_1006),
.B1(n_1016),
.B2(n_1034),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1081),
.A2(n_1088),
.B1(n_1039),
.B2(n_1092),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_R g1235 ( 
.A(n_953),
.B(n_968),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1023),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_968),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1001),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1025),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_954),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1001),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1095),
.A2(n_1097),
.B(n_1021),
.C(n_966),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_SL g1243 ( 
.A(n_1030),
.B(n_1049),
.C(n_960),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1081),
.A2(n_1032),
.B(n_1087),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1003),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1095),
.B(n_970),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1097),
.A2(n_995),
.B(n_1087),
.C(n_1075),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1003),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1201),
.A2(n_956),
.B(n_1008),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1111),
.B(n_1035),
.Y(n_1250)
);

AOI211x1_ASAP7_75t_L g1251 ( 
.A1(n_1189),
.A2(n_967),
.B(n_971),
.C(n_975),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1230),
.A2(n_1008),
.B(n_1032),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1178),
.A2(n_956),
.B(n_986),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1211),
.Y(n_1254)
);

BUFx2_ASAP7_75t_R g1255 ( 
.A(n_1208),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1244),
.A2(n_1220),
.B(n_1210),
.Y(n_1256)
);

OAI22x1_ASAP7_75t_L g1257 ( 
.A1(n_1197),
.A2(n_1030),
.B1(n_1060),
.B2(n_995),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1128),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1128),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1229),
.A2(n_1035),
.B(n_956),
.Y(n_1260)
);

NAND3x1_ASAP7_75t_L g1261 ( 
.A(n_1222),
.B(n_956),
.C(n_1035),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1106),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1116),
.B(n_1177),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1134),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1177),
.B(n_1207),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1100),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1118),
.A2(n_1102),
.B(n_1202),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_R g1268 ( 
.A(n_1109),
.B(n_1150),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1198),
.A2(n_1207),
.B1(n_1229),
.B2(n_1153),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1200),
.A2(n_1121),
.B(n_1231),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1205),
.B(n_1120),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1117),
.A2(n_1216),
.B(n_1215),
.C(n_1198),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1156),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1105),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1128),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1165),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1148),
.A2(n_1118),
.B(n_1234),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1163),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1123),
.B(n_1183),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1137),
.B(n_1151),
.Y(n_1280)
);

NAND3x1_ASAP7_75t_L g1281 ( 
.A(n_1190),
.B(n_1162),
.C(n_1194),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1206),
.A2(n_1233),
.B1(n_1127),
.B2(n_1204),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1238),
.B(n_1241),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1245),
.B(n_1248),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1112),
.A2(n_1234),
.A3(n_1219),
.B(n_1145),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1199),
.B(n_1159),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1148),
.A2(n_1101),
.B(n_1103),
.C(n_1171),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1160),
.A2(n_1164),
.B(n_1099),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1122),
.A2(n_1164),
.B(n_1160),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1247),
.A2(n_1143),
.B(n_1112),
.Y(n_1290)
);

CKINVDCx6p67_ASAP7_75t_R g1291 ( 
.A(n_1146),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1145),
.A2(n_1125),
.A3(n_1196),
.B(n_1189),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1226),
.A2(n_1130),
.B(n_1131),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1157),
.B(n_1195),
.Y(n_1294)
);

BUFx2_ASAP7_75t_R g1295 ( 
.A(n_1169),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1144),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1138),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1113),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1130),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1243),
.A2(n_1214),
.B(n_1126),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1142),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1226),
.A2(n_1129),
.B(n_1108),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1187),
.B(n_1217),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_L g1304 ( 
.A(n_1174),
.B(n_1155),
.C(n_1170),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1184),
.B(n_1132),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1161),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1107),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1181),
.A2(n_1175),
.B(n_1246),
.C(n_1212),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1192),
.A2(n_1185),
.B(n_1193),
.C(n_1155),
.Y(n_1309)
);

NOR2x1_ASAP7_75t_L g1310 ( 
.A(n_1176),
.B(n_1237),
.Y(n_1310)
);

AND3x4_ASAP7_75t_L g1311 ( 
.A(n_1217),
.B(n_1187),
.C(n_1124),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1132),
.B(n_1139),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1119),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1158),
.A2(n_1115),
.B(n_1167),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1139),
.B(n_1225),
.Y(n_1315)
);

AOI221x1_ASAP7_75t_L g1316 ( 
.A1(n_1179),
.A2(n_1114),
.B1(n_1152),
.B2(n_1147),
.C(n_1141),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1191),
.B(n_1154),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1209),
.Y(n_1318)
);

AOI221x1_ASAP7_75t_L g1319 ( 
.A1(n_1114),
.A2(n_1224),
.B1(n_1240),
.B2(n_1227),
.C(n_1218),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1213),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1186),
.A2(n_1228),
.B(n_1236),
.Y(n_1321)
);

NOR2x1_ASAP7_75t_SL g1322 ( 
.A(n_1100),
.B(n_1237),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1100),
.B(n_1232),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1224),
.A2(n_1168),
.B(n_1223),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1135),
.Y(n_1325)
);

AO32x2_ASAP7_75t_L g1326 ( 
.A1(n_1104),
.A2(n_1176),
.A3(n_1166),
.B1(n_1149),
.B2(n_1221),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1168),
.A2(n_1218),
.B(n_1227),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1172),
.B(n_1110),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1203),
.B(n_1173),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1104),
.A2(n_1239),
.A3(n_1235),
.B(n_1227),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1165),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1133),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1133),
.A2(n_1180),
.B(n_1182),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1156),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1111),
.B(n_761),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1111),
.B(n_761),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1120),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1111),
.B(n_595),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1211),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1230),
.A2(n_1244),
.B(n_1220),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1230),
.A2(n_1244),
.B(n_1220),
.Y(n_1341)
);

AOI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1198),
.A2(n_924),
.B1(n_602),
.B2(n_933),
.C(n_559),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1155),
.A2(n_924),
.B(n_603),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1140),
.A2(n_1118),
.A3(n_1198),
.B(n_1242),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1178),
.A2(n_850),
.B(n_1201),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1111),
.A2(n_951),
.B1(n_997),
.B2(n_1026),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_L g1347 ( 
.A(n_1100),
.B(n_1078),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1211),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1230),
.A2(n_1244),
.B(n_1220),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1230),
.A2(n_1244),
.B(n_1220),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1111),
.B(n_595),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1178),
.A2(n_850),
.B(n_1201),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1230),
.A2(n_1244),
.B(n_1220),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1111),
.B(n_761),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1205),
.B(n_761),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1205),
.B(n_761),
.Y(n_1356)
);

NAND2xp33_ASAP7_75t_L g1357 ( 
.A(n_1190),
.B(n_951),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1111),
.B(n_761),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1140),
.A2(n_1118),
.A3(n_1198),
.B(n_1242),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1140),
.A2(n_1118),
.A3(n_1198),
.B(n_1242),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1111),
.B(n_761),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1211),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1117),
.B(n_951),
.C(n_924),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1210),
.A2(n_1136),
.B(n_1201),
.Y(n_1364)
);

INVx5_ASAP7_75t_L g1365 ( 
.A(n_1130),
.Y(n_1365)
);

O2A1O1Ixp5_ASAP7_75t_L g1366 ( 
.A1(n_1198),
.A2(n_951),
.B(n_997),
.C(n_1027),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1198),
.A2(n_951),
.B1(n_1020),
.B2(n_740),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1111),
.B(n_595),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1130),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1111),
.A2(n_924),
.B1(n_951),
.B2(n_1026),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1210),
.A2(n_1136),
.B(n_1201),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1205),
.B(n_761),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1211),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1111),
.B(n_761),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1178),
.A2(n_850),
.B(n_1201),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1178),
.A2(n_850),
.B(n_1201),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_SL g1377 ( 
.A1(n_1196),
.A2(n_951),
.B(n_997),
.C(n_1027),
.Y(n_1377)
);

AO22x2_ASAP7_75t_L g1378 ( 
.A1(n_1198),
.A2(n_1145),
.B1(n_1189),
.B2(n_1243),
.Y(n_1378)
);

OAI22x1_ASAP7_75t_L g1379 ( 
.A1(n_1197),
.A2(n_924),
.B1(n_603),
.B2(n_590),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1102),
.A2(n_951),
.B(n_924),
.C(n_1026),
.Y(n_1380)
);

AO31x2_ASAP7_75t_L g1381 ( 
.A1(n_1140),
.A2(n_1118),
.A3(n_1198),
.B(n_1242),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1111),
.B(n_761),
.Y(n_1382)
);

O2A1O1Ixp5_ASAP7_75t_SL g1383 ( 
.A1(n_1145),
.A2(n_997),
.B(n_1189),
.C(n_1027),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1211),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1111),
.B(n_761),
.Y(n_1385)
);

AOI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1210),
.A2(n_1136),
.B(n_1201),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1178),
.A2(n_850),
.B(n_1201),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1111),
.B(n_761),
.Y(n_1388)
);

NOR2x1_ASAP7_75t_SL g1389 ( 
.A(n_1130),
.B(n_1100),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1230),
.A2(n_1244),
.B(n_1220),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1120),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1102),
.A2(n_951),
.B(n_924),
.C(n_1026),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1117),
.B(n_951),
.C(n_924),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1146),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1111),
.B(n_761),
.Y(n_1395)
);

BUFx12f_ASAP7_75t_L g1396 ( 
.A(n_1146),
.Y(n_1396)
);

AO32x2_ASAP7_75t_L g1397 ( 
.A1(n_1198),
.A2(n_1145),
.A3(n_1118),
.B1(n_1189),
.B2(n_1139),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1363),
.A2(n_1393),
.B(n_1392),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1274),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1254),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1324),
.B(n_1327),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1365),
.B(n_1266),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1351),
.A2(n_1370),
.B1(n_1363),
.B2(n_1393),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1339),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1304),
.A2(n_1378),
.B1(n_1346),
.B2(n_1312),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1290),
.A2(n_1287),
.A3(n_1289),
.B(n_1293),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1349),
.A2(n_1353),
.B(n_1350),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1342),
.A2(n_1304),
.B1(n_1370),
.B2(n_1378),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1348),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1362),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1258),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1373),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1372),
.B(n_1317),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1380),
.A2(n_1343),
.B(n_1272),
.C(n_1338),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1343),
.A2(n_1368),
.B(n_1309),
.C(n_1308),
.Y(n_1416)
);

NOR2x1_ASAP7_75t_SL g1417 ( 
.A(n_1365),
.B(n_1250),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1267),
.A2(n_1300),
.B(n_1253),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1384),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1267),
.A2(n_1300),
.B(n_1390),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1354),
.B(n_1358),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1379),
.A2(n_1311),
.B1(n_1281),
.B2(n_1374),
.Y(n_1423)
);

BUFx8_ASAP7_75t_SL g1424 ( 
.A(n_1394),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1344),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1396),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1258),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1302),
.A2(n_1345),
.B(n_1387),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1303),
.B(n_1297),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1262),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1361),
.B(n_1382),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1264),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1256),
.A2(n_1270),
.B(n_1386),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1303),
.B(n_1301),
.Y(n_1434)
);

INVxp67_ASAP7_75t_L g1435 ( 
.A(n_1280),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1291),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1277),
.B(n_1261),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1271),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1263),
.B(n_1385),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1388),
.A2(n_1395),
.B1(n_1357),
.B2(n_1315),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1296),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1329),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1305),
.A2(n_1367),
.B1(n_1269),
.B2(n_1265),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1249),
.A2(n_1319),
.B(n_1253),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1329),
.Y(n_1445)
);

NAND2x1p5_ASAP7_75t_L g1446 ( 
.A(n_1365),
.B(n_1323),
.Y(n_1446)
);

NAND2x1p5_ASAP7_75t_L g1447 ( 
.A(n_1323),
.B(n_1299),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1367),
.A2(n_1269),
.B1(n_1279),
.B2(n_1257),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1283),
.B(n_1284),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1294),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1259),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1273),
.B(n_1334),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1333),
.B(n_1282),
.Y(n_1453)
);

AO31x2_ASAP7_75t_L g1454 ( 
.A1(n_1260),
.A2(n_1352),
.A3(n_1376),
.B(n_1375),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1377),
.A2(n_1366),
.B(n_1328),
.C(n_1337),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1364),
.A2(n_1371),
.B(n_1314),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1326),
.B(n_1306),
.Y(n_1457)
);

OAI21xp33_ASAP7_75t_L g1458 ( 
.A1(n_1383),
.A2(n_1325),
.B(n_1286),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1397),
.A2(n_1331),
.B1(n_1276),
.B2(n_1285),
.Y(n_1459)
);

AOI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1288),
.A2(n_1316),
.B(n_1321),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1326),
.B(n_1278),
.Y(n_1461)
);

AOI21xp33_ASAP7_75t_L g1462 ( 
.A1(n_1307),
.A2(n_1313),
.B(n_1320),
.Y(n_1462)
);

AO21x1_ASAP7_75t_L g1463 ( 
.A1(n_1397),
.A2(n_1251),
.B(n_1326),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1251),
.A2(n_1285),
.B(n_1359),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1322),
.A2(n_1389),
.B(n_1347),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1330),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1391),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1369),
.A2(n_1310),
.B(n_1332),
.Y(n_1468)
);

CKINVDCx8_ASAP7_75t_R g1469 ( 
.A(n_1318),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1330),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1330),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1259),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1275),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1359),
.A2(n_1360),
.B(n_1381),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1292),
.A2(n_1298),
.B(n_1275),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1275),
.A2(n_1255),
.B(n_1268),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1344),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1363),
.A2(n_951),
.B(n_1393),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1254),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1363),
.A2(n_951),
.B(n_1393),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1363),
.A2(n_951),
.B(n_1393),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1363),
.A2(n_951),
.B(n_1393),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1254),
.Y(n_1484)
);

BUFx12f_ASAP7_75t_L g1485 ( 
.A(n_1394),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1254),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1254),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1295),
.Y(n_1491)
);

AND2x2_ASAP7_75t_SL g1492 ( 
.A(n_1312),
.B(n_951),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1258),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1254),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1365),
.B(n_1188),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1254),
.Y(n_1496)
);

AO31x2_ASAP7_75t_L g1497 ( 
.A1(n_1290),
.A2(n_1287),
.A3(n_1289),
.B(n_1293),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1254),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_SL g1499 ( 
.A(n_1295),
.B(n_595),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1271),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1254),
.Y(n_1501)
);

AND2x2_ASAP7_75t_SL g1502 ( 
.A(n_1312),
.B(n_951),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1380),
.A2(n_1392),
.B(n_951),
.C(n_924),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1504)
);

CKINVDCx16_ASAP7_75t_R g1505 ( 
.A(n_1268),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1351),
.A2(n_924),
.B1(n_1370),
.B2(n_1363),
.Y(n_1506)
);

AOI221x1_ASAP7_75t_L g1507 ( 
.A1(n_1304),
.A2(n_1378),
.B1(n_1277),
.B2(n_1198),
.C(n_1363),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1508)
);

NAND2x1p5_ASAP7_75t_L g1509 ( 
.A(n_1365),
.B(n_1188),
.Y(n_1509)
);

BUFx2_ASAP7_75t_SL g1510 ( 
.A(n_1274),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1355),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1394),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1363),
.A2(n_951),
.B(n_1393),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1271),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1290),
.A2(n_1293),
.B(n_1302),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1521)
);

BUFx2_ASAP7_75t_SL g1522 ( 
.A(n_1274),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1344),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1344),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1274),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1254),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1355),
.B(n_1356),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1274),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1335),
.B(n_1336),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1363),
.A2(n_951),
.B(n_1393),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1344),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1254),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1252),
.A2(n_1341),
.B(n_1340),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1414),
.B(n_1407),
.Y(n_1535)
);

CKINVDCx6p67_ASAP7_75t_R g1536 ( 
.A(n_1426),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1409),
.A2(n_1423),
.B1(n_1431),
.B2(n_1421),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1489),
.B(n_1527),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1426),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1507),
.A2(n_1456),
.B(n_1433),
.Y(n_1540)
);

NOR2xp67_ASAP7_75t_L g1541 ( 
.A(n_1435),
.B(n_1511),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1495),
.A2(n_1509),
.B(n_1449),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1495),
.A2(n_1509),
.B(n_1416),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1500),
.B(n_1517),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1409),
.A2(n_1421),
.B1(n_1431),
.B2(n_1440),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1399),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1475),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1399),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1491),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1506),
.A2(n_1481),
.B1(n_1529),
.B2(n_1515),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1455),
.A2(n_1415),
.B(n_1417),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1403),
.A2(n_1483),
.B(n_1478),
.C(n_1480),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1482),
.A2(n_1531),
.B(n_1513),
.C(n_1398),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1422),
.B(n_1439),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1512),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1475),
.Y(n_1556)
);

AND2x6_ASAP7_75t_L g1557 ( 
.A(n_1466),
.B(n_1470),
.Y(n_1557)
);

O2A1O1Ixp5_ASAP7_75t_L g1558 ( 
.A1(n_1463),
.A2(n_1460),
.B(n_1520),
.C(n_1471),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1458),
.A2(n_1435),
.B(n_1511),
.C(n_1453),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1492),
.B(n_1502),
.Y(n_1560)
);

CKINVDCx16_ASAP7_75t_R g1561 ( 
.A(n_1499),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1486),
.A2(n_1534),
.B(n_1530),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1453),
.A2(n_1443),
.B(n_1467),
.C(n_1438),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1479),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1486),
.A2(n_1534),
.B(n_1530),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1488),
.A2(n_1504),
.B(n_1508),
.Y(n_1566)
);

O2A1O1Ixp5_ASAP7_75t_L g1567 ( 
.A1(n_1428),
.A2(n_1465),
.B(n_1462),
.C(n_1434),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1492),
.B(n_1502),
.Y(n_1568)
);

INVxp67_ASAP7_75t_SL g1569 ( 
.A(n_1487),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1475),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1457),
.B(n_1461),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1450),
.B(n_1405),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1405),
.B(n_1429),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1525),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1459),
.A2(n_1443),
.B1(n_1448),
.B2(n_1453),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1434),
.B(n_1452),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1488),
.A2(n_1504),
.B(n_1508),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1448),
.A2(n_1459),
.B(n_1425),
.C(n_1477),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1490),
.B(n_1494),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1437),
.A2(n_1445),
.B1(n_1442),
.B2(n_1491),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1525),
.Y(n_1581)
);

O2A1O1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1401),
.A2(n_1533),
.B(n_1400),
.C(n_1498),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1401),
.A2(n_1432),
.B(n_1441),
.C(n_1496),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1419),
.B(n_1430),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1518),
.A2(n_1521),
.B(n_1519),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1484),
.B(n_1501),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1526),
.B(n_1473),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1437),
.A2(n_1444),
.B(n_1446),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1425),
.A2(n_1532),
.B(n_1524),
.C(n_1523),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1418),
.B(n_1472),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1476),
.B(n_1412),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1512),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1510),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1518),
.A2(n_1519),
.B(n_1521),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1437),
.A2(n_1528),
.B1(n_1522),
.B2(n_1505),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1474),
.B(n_1464),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1474),
.B(n_1528),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1464),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1406),
.Y(n_1600)
);

AOI221x1_ASAP7_75t_SL g1601 ( 
.A1(n_1424),
.A2(n_1485),
.B1(n_1436),
.B2(n_1497),
.C(n_1406),
.Y(n_1601)
);

NOR2xp67_ASAP7_75t_L g1602 ( 
.A(n_1485),
.B(n_1451),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1447),
.A2(n_1446),
.B1(n_1402),
.B2(n_1469),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1412),
.A2(n_1493),
.B1(n_1427),
.B2(n_1420),
.C(n_1447),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1412),
.B(n_1427),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1514),
.A2(n_1516),
.B(n_1408),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1451),
.B(n_1468),
.Y(n_1607)
);

OAI31xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1424),
.A2(n_1454),
.A3(n_1506),
.B(n_1393),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1454),
.A2(n_1290),
.B(n_1507),
.Y(n_1609)
);

AOI221x1_ASAP7_75t_SL g1610 ( 
.A1(n_1506),
.A2(n_1351),
.B1(n_924),
.B2(n_1393),
.C(n_1363),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1409),
.A2(n_924),
.B1(n_1351),
.B2(n_1370),
.Y(n_1611)
);

BUFx3_ASAP7_75t_L g1612 ( 
.A(n_1399),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1414),
.B(n_1407),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1421),
.B(n_1431),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1409),
.A2(n_924),
.B1(n_1351),
.B2(n_1370),
.Y(n_1615)
);

O2A1O1Ixp5_ASAP7_75t_L g1616 ( 
.A1(n_1398),
.A2(n_951),
.B(n_1300),
.C(n_997),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1414),
.B(n_1407),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1404),
.B(n_1413),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1415),
.A2(n_1503),
.B(n_1416),
.C(n_951),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1414),
.B(n_1407),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1414),
.B(n_1407),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1557),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1611),
.A2(n_1615),
.B1(n_1545),
.B2(n_1537),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1600),
.B(n_1599),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1582),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1550),
.B(n_1569),
.Y(n_1626)
);

OR2x6_ASAP7_75t_L g1627 ( 
.A(n_1589),
.B(n_1583),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1591),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1609),
.B(n_1571),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1562),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1609),
.B(n_1597),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1598),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1547),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1589),
.B(n_1551),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1551),
.B(n_1543),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1547),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1614),
.A2(n_1578),
.B1(n_1619),
.B2(n_1575),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1557),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1556),
.B(n_1570),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1557),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1570),
.B(n_1590),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1557),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1553),
.B(n_1552),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1558),
.A2(n_1567),
.B(n_1578),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1557),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1540),
.B(n_1560),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1543),
.B(n_1542),
.Y(n_1647)
);

AO21x1_ASAP7_75t_SL g1648 ( 
.A1(n_1568),
.A2(n_1572),
.B(n_1573),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1616),
.A2(n_1604),
.B(n_1619),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1559),
.A2(n_1563),
.B(n_1607),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1562),
.A2(n_1586),
.B(n_1577),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1618),
.B(n_1564),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1592),
.B(n_1579),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1585),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1584),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1565),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1610),
.B(n_1554),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1587),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1588),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1601),
.B(n_1608),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1656),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1638),
.B(n_1605),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1624),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1541),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1646),
.B(n_1586),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1623),
.A2(n_1538),
.B1(n_1621),
.B2(n_1535),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1629),
.B(n_1595),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1624),
.Y(n_1669)
);

NAND4xp25_ASAP7_75t_L g1670 ( 
.A(n_1643),
.B(n_1544),
.C(n_1617),
.D(n_1613),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1631),
.B(n_1577),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1622),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1632),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1646),
.B(n_1566),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1631),
.B(n_1577),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1643),
.B(n_1596),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1636),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1630),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1631),
.B(n_1606),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1628),
.B(n_1620),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1630),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1632),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1633),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1637),
.B(n_1603),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1636),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1623),
.A2(n_1536),
.B1(n_1561),
.B2(n_1576),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1633),
.Y(n_1687)
);

AOI31xp33_ASAP7_75t_L g1688 ( 
.A1(n_1684),
.A2(n_1637),
.A3(n_1660),
.B(n_1625),
.Y(n_1688)
);

OAI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1684),
.A2(n_1660),
.B(n_1625),
.C(n_1657),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1676),
.A2(n_1657),
.B1(n_1635),
.B2(n_1649),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1677),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1677),
.Y(n_1692)
);

NOR2x1p5_ASAP7_75t_L g1693 ( 
.A(n_1670),
.B(n_1536),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1676),
.A2(n_1635),
.B1(n_1648),
.B2(n_1634),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1687),
.Y(n_1695)
);

OR2x6_ASAP7_75t_L g1696 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1672),
.B(n_1640),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1683),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1661),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1672),
.B(n_1640),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1685),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1634),
.Y(n_1703)
);

NAND2xp33_ASAP7_75t_R g1704 ( 
.A(n_1664),
.B(n_1549),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1705)
);

OAI33xp33_ASAP7_75t_L g1706 ( 
.A1(n_1670),
.A2(n_1664),
.A3(n_1680),
.B1(n_1626),
.B2(n_1655),
.B3(n_1674),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1686),
.A2(n_1635),
.B1(n_1634),
.B2(n_1593),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1686),
.B(n_1644),
.C(n_1626),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1668),
.B(n_1669),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1683),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1666),
.A2(n_1635),
.B1(n_1648),
.B2(n_1634),
.Y(n_1712)
);

OAI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1666),
.A2(n_1635),
.B1(n_1634),
.B2(n_1647),
.C(n_1627),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1687),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1685),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1662),
.A2(n_1635),
.B1(n_1648),
.B2(n_1650),
.Y(n_1716)
);

NAND2xp33_ASAP7_75t_SL g1717 ( 
.A(n_1672),
.B(n_1593),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1673),
.A2(n_1644),
.B(n_1649),
.C(n_1641),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1662),
.A2(n_1650),
.B1(n_1647),
.B2(n_1644),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1673),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1682),
.A2(n_1649),
.B1(n_1644),
.B2(n_1650),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1682),
.A2(n_1627),
.B1(n_1641),
.B2(n_1647),
.C(n_1594),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1683),
.B(n_1639),
.Y(n_1723)
);

OAI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1665),
.A2(n_1644),
.B(n_1649),
.C(n_1652),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1679),
.A2(n_1658),
.B1(n_1654),
.B2(n_1652),
.C(n_1659),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1668),
.B(n_1645),
.Y(n_1726)
);

INVxp33_ASAP7_75t_L g1727 ( 
.A(n_1662),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1700),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1698),
.Y(n_1729)
);

OA21x2_ASAP7_75t_L g1730 ( 
.A1(n_1721),
.A2(n_1651),
.B(n_1678),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1698),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1710),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1695),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1714),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1700),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_SL g1736 ( 
.A1(n_1688),
.A2(n_1645),
.B(n_1580),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1710),
.Y(n_1737)
);

INVx4_ASAP7_75t_SL g1738 ( 
.A(n_1707),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1691),
.Y(n_1739)
);

CKINVDCx20_ASAP7_75t_R g1740 ( 
.A(n_1720),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1698),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1698),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1711),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1691),
.B(n_1692),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1692),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1709),
.A2(n_1649),
.B(n_1627),
.Y(n_1746)
);

INVx4_ASAP7_75t_SL g1747 ( 
.A(n_1707),
.Y(n_1747)
);

NAND2x1_ASAP7_75t_L g1748 ( 
.A(n_1711),
.B(n_1627),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1702),
.B(n_1671),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1702),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1715),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1701),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1715),
.Y(n_1753)
);

OA21x2_ASAP7_75t_L g1754 ( 
.A1(n_1718),
.A2(n_1681),
.B(n_1678),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1699),
.Y(n_1755)
);

INVx4_ASAP7_75t_SL g1756 ( 
.A(n_1696),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1694),
.B(n_1653),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1723),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1725),
.B(n_1671),
.Y(n_1759)
);

INVx4_ASAP7_75t_SL g1760 ( 
.A(n_1696),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1733),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1728),
.Y(n_1762)
);

NAND2x1p5_ASAP7_75t_L g1763 ( 
.A(n_1748),
.B(n_1690),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1729),
.B(n_1727),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1759),
.B(n_1671),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1756),
.B(n_1696),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1759),
.B(n_1675),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1739),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1745),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_SL g1770 ( 
.A(n_1736),
.B(n_1709),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1729),
.B(n_1697),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1731),
.B(n_1697),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1731),
.B(n_1705),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1745),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1750),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1751),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1741),
.B(n_1705),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1758),
.B(n_1723),
.Y(n_1778)
);

NAND5xp2_ASAP7_75t_SL g1779 ( 
.A(n_1736),
.B(n_1689),
.C(n_1746),
.D(n_1724),
.E(n_1720),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1741),
.B(n_1708),
.Y(n_1780)
);

OAI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1746),
.A2(n_1690),
.B1(n_1713),
.B2(n_1704),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1742),
.B(n_1708),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1742),
.B(n_1726),
.Y(n_1783)
);

AND2x4_ASAP7_75t_SL g1784 ( 
.A(n_1740),
.B(n_1647),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1753),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1752),
.B(n_1726),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1752),
.B(n_1696),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1734),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1758),
.B(n_1665),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1728),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1728),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_L g1792 ( 
.A(n_1754),
.B(n_1719),
.C(n_1716),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1756),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1735),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1756),
.B(n_1696),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1753),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1756),
.B(n_1703),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1756),
.B(n_1703),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1744),
.B(n_1667),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1760),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1738),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1744),
.B(n_1693),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1801),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1761),
.B(n_1743),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1788),
.B(n_1749),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1768),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1768),
.Y(n_1807)
);

NAND2x1_ASAP7_75t_L g1808 ( 
.A(n_1793),
.B(n_1800),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1793),
.B(n_1738),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1770),
.B(n_1757),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1769),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1800),
.B(n_1795),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1770),
.B(n_1732),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1774),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1781),
.B(n_1732),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1802),
.B(n_1801),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1774),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1801),
.B(n_1737),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1762),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1795),
.B(n_1738),
.Y(n_1821)
);

INVxp67_ASAP7_75t_SL g1822 ( 
.A(n_1763),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1801),
.B(n_1737),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1775),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1765),
.B(n_1755),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1775),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1778),
.B(n_1754),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1776),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1762),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1766),
.B(n_1738),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1776),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1765),
.B(n_1693),
.Y(n_1832)
);

AND3x1_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1747),
.C(n_1738),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1785),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1767),
.B(n_1747),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1767),
.B(n_1747),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1771),
.B(n_1747),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1785),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1762),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1807),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1811),
.A2(n_1779),
.B(n_1792),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1804),
.B(n_1778),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1807),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1810),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1833),
.A2(n_1792),
.B1(n_1779),
.B2(n_1722),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1810),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1812),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1816),
.B(n_1799),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1813),
.B(n_1796),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1808),
.B(n_1539),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1821),
.B(n_1797),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1812),
.Y(n_1852)
);

INVx3_ASAP7_75t_SL g1853 ( 
.A(n_1803),
.Y(n_1853)
);

INVx3_ASAP7_75t_SL g1854 ( 
.A(n_1803),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1813),
.B(n_1747),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1808),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1821),
.B(n_1787),
.Y(n_1857)
);

INVxp67_ASAP7_75t_L g1858 ( 
.A(n_1803),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1830),
.A2(n_1798),
.B1(n_1766),
.B2(n_1763),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1834),
.Y(n_1860)
);

AND2x4_ASAP7_75t_SL g1861 ( 
.A(n_1830),
.B(n_1766),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1834),
.Y(n_1862)
);

AO21x2_ASAP7_75t_L g1863 ( 
.A1(n_1822),
.A2(n_1796),
.B(n_1791),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1806),
.B(n_1771),
.Y(n_1864)
);

CKINVDCx16_ASAP7_75t_R g1865 ( 
.A(n_1809),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1809),
.B(n_1787),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1845),
.A2(n_1830),
.B1(n_1837),
.B2(n_1836),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1865),
.B(n_1817),
.Y(n_1868)
);

OAI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1841),
.A2(n_1763),
.B1(n_1835),
.B2(n_1814),
.C(n_1832),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1863),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1845),
.A2(n_1798),
.B1(n_1766),
.B2(n_1717),
.Y(n_1871)
);

O2A1O1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1841),
.A2(n_1823),
.B(n_1819),
.C(n_1827),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1855),
.B(n_1798),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1849),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1856),
.A2(n_1848),
.B1(n_1850),
.B2(n_1854),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1861),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1851),
.B(n_1772),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_SL g1878 ( 
.A1(n_1850),
.A2(n_1555),
.B1(n_1539),
.B2(n_1549),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1866),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1857),
.B(n_1815),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1859),
.A2(n_1798),
.B(n_1825),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1858),
.B(n_1818),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_L g1883 ( 
.A(n_1850),
.B(n_1826),
.C(n_1824),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1855),
.A2(n_1784),
.B1(n_1706),
.B2(n_1748),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1849),
.Y(n_1885)
);

OAI31xp33_ASAP7_75t_L g1886 ( 
.A1(n_1856),
.A2(n_1784),
.A3(n_1827),
.B(n_1805),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1842),
.B(n_1805),
.Y(n_1887)
);

OAI221xp5_ASAP7_75t_SL g1888 ( 
.A1(n_1858),
.A2(n_1831),
.B1(n_1828),
.B2(n_1838),
.C(n_1712),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1870),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1876),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1878),
.B(n_1555),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1868),
.B(n_1853),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1879),
.B(n_1864),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1870),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_SL g1895 ( 
.A1(n_1869),
.A2(n_1883),
.B1(n_1881),
.B2(n_1874),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1887),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1877),
.B(n_1853),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1882),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1873),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1880),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1895),
.A2(n_1872),
.B(n_1875),
.Y(n_1901)
);

AOI221x1_ASAP7_75t_L g1902 ( 
.A1(n_1894),
.A2(n_1885),
.B1(n_1843),
.B2(n_1840),
.C(n_1844),
.Y(n_1902)
);

OAI21xp33_ASAP7_75t_L g1903 ( 
.A1(n_1895),
.A2(n_1867),
.B(n_1871),
.Y(n_1903)
);

AOI211x1_ASAP7_75t_SL g1904 ( 
.A1(n_1899),
.A2(n_1864),
.B(n_1886),
.C(n_1829),
.Y(n_1904)
);

AOI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1890),
.A2(n_1888),
.B1(n_1884),
.B2(n_1847),
.C(n_1846),
.Y(n_1905)
);

OAI21xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1896),
.A2(n_1889),
.B(n_1897),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1891),
.A2(n_1888),
.B(n_1889),
.Y(n_1907)
);

AOI211xp5_ASAP7_75t_L g1908 ( 
.A1(n_1892),
.A2(n_1852),
.B(n_1862),
.C(n_1860),
.Y(n_1908)
);

NAND4xp25_ASAP7_75t_SL g1909 ( 
.A(n_1893),
.B(n_1764),
.C(n_1772),
.D(n_1773),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1900),
.B(n_1773),
.Y(n_1910)
);

OAI21xp33_ASAP7_75t_SL g1911 ( 
.A1(n_1901),
.A2(n_1898),
.B(n_1829),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1903),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1904),
.A2(n_1784),
.B(n_1764),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1906),
.A2(n_1839),
.B(n_1820),
.Y(n_1914)
);

AOI211xp5_ASAP7_75t_L g1915 ( 
.A1(n_1907),
.A2(n_1602),
.B(n_1839),
.C(n_1820),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1910),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1916),
.B(n_1908),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1913),
.B(n_1909),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1914),
.Y(n_1919)
);

NAND3xp33_ASAP7_75t_L g1920 ( 
.A(n_1915),
.B(n_1905),
.C(n_1902),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1911),
.B(n_1863),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1912),
.B(n_1777),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1916),
.B(n_1546),
.Y(n_1923)
);

NAND2xp33_ASAP7_75t_R g1924 ( 
.A(n_1919),
.B(n_1754),
.Y(n_1924)
);

NAND2xp33_ASAP7_75t_L g1925 ( 
.A(n_1923),
.B(n_1777),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1920),
.A2(n_1760),
.B1(n_1794),
.B2(n_1791),
.Y(n_1926)
);

AOI211x1_ASAP7_75t_L g1927 ( 
.A1(n_1917),
.A2(n_1780),
.B(n_1786),
.C(n_1782),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1922),
.B(n_1780),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1928),
.B(n_1918),
.Y(n_1929)
);

NAND4xp75_ASAP7_75t_L g1930 ( 
.A(n_1927),
.B(n_1921),
.C(n_1754),
.D(n_1730),
.Y(n_1930)
);

OAI221xp5_ASAP7_75t_L g1931 ( 
.A1(n_1926),
.A2(n_1925),
.B1(n_1924),
.B2(n_1791),
.C(n_1790),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1930),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1932),
.Y(n_1933)
);

NOR2x1p5_ASAP7_75t_L g1934 ( 
.A(n_1933),
.B(n_1929),
.Y(n_1934)
);

HB1xp67_ASAP7_75t_L g1935 ( 
.A(n_1933),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1935),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1934),
.B(n_1931),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1936),
.B(n_1790),
.Y(n_1938)
);

CKINVDCx20_ASAP7_75t_R g1939 ( 
.A(n_1937),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1939),
.A2(n_1790),
.B1(n_1794),
.B2(n_1789),
.Y(n_1940)
);

OA21x2_ASAP7_75t_L g1941 ( 
.A1(n_1940),
.A2(n_1938),
.B(n_1794),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1941),
.A2(n_1786),
.B1(n_1783),
.B2(n_1782),
.Y(n_1942)
);

XOR2xp5_ASAP7_75t_L g1943 ( 
.A(n_1942),
.B(n_1546),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_SL g1944 ( 
.A1(n_1943),
.A2(n_1548),
.B1(n_1574),
.B2(n_1612),
.Y(n_1944)
);

AOI211xp5_ASAP7_75t_L g1945 ( 
.A1(n_1944),
.A2(n_1581),
.B(n_1612),
.C(n_1574),
.Y(n_1945)
);


endmodule