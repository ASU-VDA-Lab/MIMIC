module fake_jpeg_16419_n_113 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_11),
.B(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_17),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_12),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_14),
.B(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_27),
.B1(n_26),
.B2(n_14),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_12),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_51),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_22),
.B(n_15),
.C(n_11),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_47),
.B(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_44),
.B1(n_33),
.B2(n_30),
.Y(n_60)
);

OAI22x1_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_13),
.B1(n_37),
.B2(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_13),
.C(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_20),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_22),
.CON(n_47),
.SN(n_47)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_35),
.B(n_21),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_32),
.B1(n_14),
.B2(n_16),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_39),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_18),
.C(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_66),
.B1(n_21),
.B2(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_30),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_36),
.B1(n_18),
.B2(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_74),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_58),
.B(n_54),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_62),
.A2(n_50),
.B(n_2),
.C(n_3),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_9),
.C(n_2),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_59),
.C(n_57),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_9),
.B1(n_2),
.B2(n_4),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_66),
.B1(n_63),
.B2(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_83),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_88),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_64),
.C(n_65),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_77),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_77),
.B1(n_72),
.B2(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_83),
.C(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_72),
.C(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_1),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_104),
.Y(n_107)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_89),
.A3(n_90),
.B1(n_96),
.B2(n_93),
.C1(n_72),
.C2(n_8),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_105),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_SL g109 ( 
.A(n_106),
.B(n_5),
.C(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_109),
.B(n_8),
.Y(n_112)
);

OAI321xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_107),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C(n_5),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.Y(n_113)
);


endmodule