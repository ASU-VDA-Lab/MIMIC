module fake_jpeg_6754_n_214 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_214);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_35),
.B(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_14),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_49),
.Y(n_52)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_41),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_4),
.B(n_5),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_23),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_14),
.B(n_4),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_51),
.Y(n_87)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_107)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_59),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_20),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_33),
.A2(n_26),
.B1(n_22),
.B2(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_84),
.B1(n_86),
.B2(n_9),
.Y(n_111)
);

OAI221xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.C(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_63),
.Y(n_110)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_71),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_51),
.B1(n_68),
.B2(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_34),
.A2(n_28),
.B1(n_27),
.B2(n_30),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_16),
.B1(n_25),
.B2(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_38),
.B(n_15),
.Y(n_71)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_34),
.B(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_15),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_6),
.Y(n_103)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_22),
.B1(n_24),
.B2(n_16),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_16),
.C(n_22),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_90),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_89),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_95),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_25),
.C(n_13),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_103),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_107),
.B1(n_66),
.B2(n_85),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_5),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_69),
.B(n_52),
.C(n_66),
.D(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_52),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_8),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_75),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_74),
.B(n_77),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_120),
.C(n_104),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_69),
.B1(n_68),
.B2(n_53),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_118),
.B(n_135),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_122),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_57),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_59),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_57),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_56),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_92),
.B1(n_94),
.B2(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_63),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_97),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_136),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_78),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_133),
.A2(n_126),
.B(n_127),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_153),
.B(n_113),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_132),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_150),
.C(n_151),
.Y(n_158)
);

NAND4xp25_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_72),
.C(n_94),
.D(n_50),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_142),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_96),
.B1(n_107),
.B2(n_88),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_124),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_118),
.C(n_116),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_103),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_114),
.B1(n_115),
.B2(n_112),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_98),
.Y(n_153)
);

OAI211xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_148),
.B(n_156),
.C(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_109),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_167),
.B(n_145),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_171),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_114),
.B1(n_112),
.B2(n_120),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_151),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_170),
.B1(n_145),
.B2(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_137),
.B1(n_149),
.B2(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_153),
.B1(n_143),
.B2(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_141),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_150),
.C(n_156),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_139),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_183),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_161),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_171),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_176),
.C(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_172),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_189),
.B(n_193),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_163),
.B(n_166),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_181),
.B(n_175),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_125),
.B(n_122),
.C(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_123),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_138),
.Y(n_193)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_197),
.A2(n_198),
.B(n_189),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_182),
.B(n_178),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_203),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_160),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_201),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_192),
.A3(n_185),
.B1(n_179),
.B2(n_121),
.C1(n_129),
.C2(n_142),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_203),
.Y(n_211)
);

AOI211xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_192),
.B(n_135),
.C(n_12),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_135),
.B(n_92),
.Y(n_209)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_209),
.B(n_211),
.CI(n_210),
.CON(n_212),
.SN(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_211),
.A2(n_205),
.B(n_12),
.C(n_11),
.Y(n_213)
);


endmodule