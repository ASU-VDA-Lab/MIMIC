module fake_jpeg_13240_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_13),
.B(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_26),
.B(n_31),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

INVx8_ASAP7_75t_SL g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_21),
.C(n_47),
.Y(n_82)
);

BUFx2_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_64),
.Y(n_95)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_91),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_55),
.B1(n_74),
.B2(n_53),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_99),
.B1(n_76),
.B2(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_75),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_61),
.B(n_52),
.C(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_0),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_68),
.B1(n_54),
.B2(n_66),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_61),
.C(n_70),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_24),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_116),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_75),
.B(n_73),
.C(n_65),
.Y(n_107)
);

AO21x1_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_109),
.B(n_16),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_0),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_108),
.B(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_1),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_76),
.B(n_72),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_14),
.B(n_45),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_114)
);

OR2x2_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_15),
.Y(n_140)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_22),
.C(n_46),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_51),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_125),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_6),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_132),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_8),
.C(n_9),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_112),
.C(n_20),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_101),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_141),
.B1(n_44),
.B2(n_40),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_12),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_12),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_138),
.A2(n_17),
.B1(n_28),
.B2(n_35),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_14),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_138),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_121),
.B(n_123),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_146),
.C(n_149),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_37),
.C(n_38),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_154),
.B(n_156),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_39),
.C(n_41),
.Y(n_149)
);

XOR2x2_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_42),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_133),
.C(n_126),
.Y(n_155)
);

AND2x4_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_141),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_156),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_159),
.B(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_150),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_165),
.B(n_151),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_163),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_161),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_170),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_158),
.C(n_144),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_151),
.Y(n_173)
);


endmodule