module fake_jpeg_28733_n_69 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_36),
.B1(n_5),
.B2(n_6),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_10),
.B1(n_24),
.B2(n_23),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_25),
.B1(n_21),
.B2(n_20),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_26),
.B1(n_2),
.B2(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_9),
.B1(n_19),
.B2(n_47),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_29),
.B(n_31),
.Y(n_42)
);

XNOR2x2_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_50),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_7),
.B(n_8),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_9),
.C(n_43),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_58),
.B(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_34),
.B1(n_14),
.B2(n_17),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_57),
.B1(n_55),
.B2(n_54),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_18),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_63),
.Y(n_65)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_53),
.Y(n_67)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_51),
.B(n_60),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.B1(n_61),
.B2(n_52),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_65),
.C(n_59),
.Y(n_69)
);


endmodule