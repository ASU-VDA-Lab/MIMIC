module real_jpeg_31939_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_620;
wire n_578;
wire n_328;
wire n_456;
wire n_366;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_0),
.Y(n_209)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_0),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_0),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_1),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_1),
.A2(n_262),
.B1(n_346),
.B2(n_351),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_1),
.A2(n_119),
.B1(n_262),
.B2(n_537),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_1),
.A2(n_262),
.B1(n_590),
.B2(n_591),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_2),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_2),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_2),
.A2(n_287),
.B1(n_397),
.B2(n_400),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_2),
.A2(n_287),
.B1(n_537),
.B2(n_571),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_2),
.A2(n_287),
.B1(n_579),
.B2(n_580),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_4),
.A2(n_289),
.B1(n_292),
.B2(n_296),
.Y(n_288)
);

INVx2_ASAP7_75t_R g296 ( 
.A(n_4),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_4),
.A2(n_296),
.B1(n_431),
.B2(n_435),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_4),
.A2(n_296),
.B1(n_489),
.B2(n_492),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_4),
.A2(n_296),
.B1(n_554),
.B2(n_558),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

AOI21x1_ASAP7_75t_L g266 ( 
.A1(n_5),
.A2(n_267),
.B(n_271),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_5),
.A2(n_65),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_5),
.A2(n_65),
.B1(n_422),
.B2(n_426),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_6),
.A2(n_251),
.B(n_255),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_6),
.B(n_364),
.Y(n_363)
);

OAI32xp33_ASAP7_75t_L g497 ( 
.A1(n_6),
.A2(n_126),
.A3(n_498),
.B1(n_501),
.B2(n_507),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_6),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_6),
.B(n_157),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_6),
.A2(n_412),
.B1(n_589),
.B2(n_597),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_6),
.A2(n_508),
.B1(n_615),
.B2(n_620),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_7),
.A2(n_30),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx2_ASAP7_75t_R g236 ( 
.A(n_7),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_7),
.A2(n_236),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_7),
.A2(n_186),
.B1(n_236),
.B2(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_7),
.A2(n_236),
.B1(n_515),
.B2(n_519),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_9),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_10),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_10),
.Y(n_522)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_12),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_12),
.A2(n_117),
.B1(n_160),
.B2(n_164),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_12),
.A2(n_117),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_13),
.A2(n_33),
.B1(n_162),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_13),
.A2(n_33),
.B1(n_319),
.B2(n_322),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_13),
.A2(n_33),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

CKINVDCx11_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_15),
.A2(n_146),
.B1(n_152),
.B2(n_155),
.Y(n_145)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_15),
.A2(n_155),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_15),
.A2(n_155),
.B1(n_220),
.B2(n_371),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_16),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_16),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_16),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_17),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_17),
.Y(n_138)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_19),
.A2(n_79),
.B1(n_85),
.B2(n_86),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_19),
.A2(n_86),
.B1(n_162),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_19),
.A2(n_86),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_19),
.A2(n_86),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_241),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_239),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_176),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_25),
.B(n_176),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_169),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_73),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_27),
.B(n_168),
.C(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_27),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_27),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_646)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B(n_53),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_28),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_37),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_37),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_38),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_39),
.A2(n_54),
.B1(n_395),
.B2(n_402),
.Y(n_394)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_41),
.Y(n_258)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_44),
.Y(n_428)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_45),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_45),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_45),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_45),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_48),
.Y(n_303)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_48),
.Y(n_312)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_50),
.Y(n_291)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NAND2x1p5_ASAP7_75t_L g234 ( 
.A(n_54),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_64),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_65),
.B(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_68),
.A2(n_299),
.A3(n_304),
.B1(n_308),
.B2(n_316),
.Y(n_298)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_72),
.Y(n_257)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_72),
.Y(n_401)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_72),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_87),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_75),
.A2(n_250),
.B1(n_258),
.B2(n_259),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_75),
.A2(n_76),
.B1(n_430),
.B2(n_436),
.Y(n_429)
);

OAI22x1_ASAP7_75t_L g446 ( 
.A1(n_75),
.A2(n_258),
.B1(n_396),
.B2(n_430),
.Y(n_446)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_82),
.Y(n_238)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_83),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_123),
.B1(n_124),
.B2(n_168),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_88),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_88),
.A2(n_168),
.B1(n_170),
.B2(n_181),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_100),
.B(n_113),
.Y(n_88)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_89),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_89),
.A2(n_100),
.B1(n_195),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_89),
.A2(n_100),
.B1(n_266),
.B2(n_273),
.Y(n_265)
);

OAI22x1_ASAP7_75t_SL g375 ( 
.A1(n_89),
.A2(n_100),
.B1(n_266),
.B2(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_89),
.A2(n_100),
.B1(n_225),
.B2(n_376),
.Y(n_417)
);

OAI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_89),
.A2(n_100),
.B1(n_273),
.B2(n_487),
.Y(n_486)
);

OAI22x1_ASAP7_75t_L g568 ( 
.A1(n_89),
.A2(n_100),
.B1(n_569),
.B2(n_570),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_89),
.B(n_508),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AO21x2_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_101),
.B(n_108),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_91),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_91)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_92),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_93),
.Y(n_223)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_93),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_93),
.Y(n_557)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_93),
.Y(n_561)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_96),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_97),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_107),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_107),
.Y(n_494)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_107),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_121),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_122),
.Y(n_276)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_145),
.B1(n_156),
.B2(n_159),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_125),
.A2(n_145),
.B1(n_156),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_125),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_125),
.A2(n_156),
.B1(n_288),
.B2(n_388),
.Y(n_387)
);

OAI22x1_ASAP7_75t_L g444 ( 
.A1(n_125),
.A2(n_156),
.B1(n_388),
.B2(n_421),
.Y(n_444)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_132),
.B(n_139),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_127),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_128),
.Y(n_315)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_138),
.Y(n_286)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_139)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_141),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_142),
.Y(n_226)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_151),
.Y(n_295)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_156),
.A2(n_281),
.B1(n_283),
.B2(n_288),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_156),
.A2(n_283),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_172),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_157),
.A2(n_185),
.B1(n_282),
.B2(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_158),
.A2(n_281),
.B1(n_345),
.B2(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_163),
.Y(n_351)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_175),
.Y(n_307)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_175),
.Y(n_393)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_175),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.C(n_203),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_179),
.A2(n_180),
.B1(n_646),
.B2(n_647),
.Y(n_645)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_183),
.B(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_184),
.B(n_189),
.Y(n_454)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_188),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B1(n_201),
.B2(n_202),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_190),
.A2(n_530),
.B1(n_535),
.B2(n_536),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_190),
.A2(n_202),
.B1(n_488),
.B2(n_624),
.Y(n_623)
);

OA21x2_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B(n_193),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g539 ( 
.A1(n_192),
.A2(n_540),
.B(n_543),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_193),
.Y(n_535)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_203),
.B(n_645),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_206),
.B(n_231),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g455 ( 
.A(n_205),
.B(n_456),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_224),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_206),
.B(n_224),
.Y(n_440)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_206),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_210),
.B(n_217),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_209),
.Y(n_374)
);

INVx4_ASAP7_75t_SL g597 ( 
.A(n_209),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_210),
.A2(n_318),
.B1(n_327),
.B2(n_329),
.Y(n_317)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_210),
.Y(n_412)
);

AO22x1_ASAP7_75t_L g513 ( 
.A1(n_210),
.A2(n_327),
.B1(n_358),
.B2(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_211),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_211),
.A2(n_330),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_211),
.A2(n_578),
.B1(n_589),
.B2(n_592),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_215),
.Y(n_416)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_216),
.Y(n_321)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_216),
.Y(n_359)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_218),
.A2(n_370),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_230),
.Y(n_571)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_232),
.B(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_235),
.Y(n_436)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_640),
.B(n_648),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_478),
.B(n_635),
.Y(n_243)
);

NAND4xp25_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_406),
.C(n_458),
.D(n_471),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_365),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_246),
.B(n_365),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_297),
.C(n_342),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_247),
.B(n_481),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_264),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_249),
.B(n_265),
.C(n_280),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_257),
.Y(n_435)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_258),
.Y(n_364)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_259),
.Y(n_402)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_280),
.Y(n_264)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_295),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_297),
.B(n_342),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_317),
.B1(n_335),
.B2(n_341),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_298),
.B(n_341),
.Y(n_405)
);

OAI32xp33_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_304),
.A3(n_308),
.B1(n_316),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

AO22x1_ASAP7_75t_SL g352 ( 
.A1(n_318),
.A2(n_353),
.B1(n_357),
.B2(n_358),
.Y(n_352)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_325),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_326),
.Y(n_542)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_326),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_326),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_352),
.C(n_362),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_343),
.B(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_352),
.B(n_363),
.Y(n_484)
);

INVx3_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_356),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_356),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_356),
.Y(n_601)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_357),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_357),
.A2(n_373),
.B1(n_577),
.B2(n_584),
.Y(n_576)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_384),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_382),
.B2(n_383),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_375),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_369),
.B(n_375),
.Y(n_447)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

BUFx4f_ASAP7_75t_SL g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_380),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_383),
.B(n_385),
.C(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_405),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_394),
.B1(n_403),
.B2(n_404),
.Y(n_386)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_387),
.Y(n_403)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_394),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

A2O1A1O1Ixp25_ASAP7_75t_L g635 ( 
.A1(n_406),
.A2(n_458),
.B(n_636),
.C(n_638),
.D(n_639),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_448),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_407),
.B(n_448),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_439),
.C(n_441),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_418),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_438),
.C(n_450),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_411),
.B(n_417),
.Y(n_468)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

OAI22xp33_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_429),
.B1(n_437),
.B2(n_438),
.Y(n_418)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_429),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_442),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.C(n_447),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_443),
.A2(n_444),
.B1(n_446),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_451),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_449),
.B(n_642),
.C(n_643),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_453),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g642 ( 
.A(n_455),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_469),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_459),
.B(n_469),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_464),
.C(n_468),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.C(n_467),
.Y(n_464)
);

MAJx2_ASAP7_75t_L g475 ( 
.A(n_465),
.B(n_466),
.C(n_467),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_474),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_472),
.B(n_474),
.C(n_637),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

AOI21x1_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_523),
.B(n_634),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_482),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_SL g634 ( 
.A(n_480),
.B(n_482),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_485),
.C(n_495),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g629 ( 
.A(n_483),
.B(n_630),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_485),
.A2(n_496),
.B(n_631),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_486),
.B(n_496),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_494),
.Y(n_532)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_513),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g611 ( 
.A(n_497),
.B(n_513),
.Y(n_611)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_504),
.Y(n_534)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_505),
.Y(n_537)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_509),
.Y(n_507)
);

OAI21xp33_ASAP7_75t_SL g530 ( 
.A1(n_508),
.A2(n_531),
.B(n_533),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_534),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_508),
.B(n_600),
.Y(n_599)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_514),
.Y(n_565)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_522),
.Y(n_546)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_522),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_524),
.A2(n_628),
.B(n_633),
.Y(n_523)
);

AOI21x1_ASAP7_75t_L g524 ( 
.A1(n_525),
.A2(n_608),
.B(n_627),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_574),
.B(n_607),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_550),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_527),
.B(n_550),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_528),
.B(n_538),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_528),
.A2(n_529),
.B1(n_538),
.B2(n_539),
.Y(n_585)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_533),
.A2(n_544),
.B(n_547),
.Y(n_543)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_536),
.Y(n_569)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_545),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_551),
.B(n_566),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_551),
.B(n_568),
.C(n_572),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_552),
.A2(n_553),
.B1(n_562),
.B2(n_565),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_553),
.Y(n_584)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_556),
.Y(n_579)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_567),
.A2(n_568),
.B1(n_572),
.B2(n_573),
.Y(n_566)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_567),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_568),
.Y(n_573)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_575),
.A2(n_586),
.B(n_606),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_585),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_576),
.B(n_585),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_579),
.Y(n_591)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_587),
.A2(n_595),
.B(n_605),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_594),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_588),
.B(n_594),
.Y(n_605)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_596),
.B(n_598),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g598 ( 
.A(n_599),
.B(n_602),
.Y(n_598)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_609),
.B(n_610),
.Y(n_608)
);

NOR2x1_ASAP7_75t_SL g627 ( 
.A(n_609),
.B(n_610),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_611),
.B(n_612),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_611),
.B(n_623),
.C(n_626),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_613),
.A2(n_623),
.B1(n_625),
.B2(n_626),
.Y(n_612)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_613),
.Y(n_626)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_623),
.Y(n_625)
);

NOR2x1_ASAP7_75t_SL g628 ( 
.A(n_629),
.B(n_632),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_629),
.B(n_632),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_SL g640 ( 
.A(n_641),
.B(n_644),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_641),
.B(n_644),
.Y(n_649)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_646),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);


endmodule