module fake_jpeg_12937_n_607 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_607);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_607;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_0),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_64),
.Y(n_124)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_62),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_67),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_76),
.Y(n_128)
);

INVx5_ASAP7_75t_SL g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_69),
.Y(n_143)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_73),
.Y(n_197)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_87),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_42),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_84),
.A2(n_23),
.B1(n_55),
.B2(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_14),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_89),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_21),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_96),
.B(n_103),
.Y(n_178)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_100),
.Y(n_201)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_21),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_20),
.B(n_14),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_104),
.B(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_106),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_21),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_20),
.B(n_14),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_112),
.B(n_115),
.Y(n_191)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_45),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_8),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_42),
.Y(n_121)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_125),
.B(n_136),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_33),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_132),
.B(n_158),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_41),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_133),
.B(n_169),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_63),
.B(n_33),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_93),
.B(n_49),
.CON(n_139),
.SN(n_139)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_120),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_84),
.A2(n_49),
.B(n_37),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_142),
.B(n_186),
.Y(n_205)
);

BUFx4f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_24),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_67),
.A2(n_42),
.B1(n_58),
.B2(n_51),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_16),
.B1(n_46),
.B2(n_48),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

BUFx16f_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_82),
.B(n_53),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_168),
.B(n_172),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_63),
.B(n_53),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_62),
.A2(n_49),
.B1(n_45),
.B2(n_26),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_32),
.B1(n_55),
.B2(n_50),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_54),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_91),
.B(n_54),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_188),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_121),
.B(n_49),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_72),
.B(n_57),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_187),
.B(n_17),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_92),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_32),
.B1(n_55),
.B2(n_23),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_81),
.B(n_26),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_22),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_70),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_91),
.B(n_57),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_37),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_94),
.A2(n_58),
.B1(n_16),
.B2(n_51),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_46),
.C(n_48),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_206),
.Y(n_315)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_207),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_133),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_208),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_122),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_209),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_212),
.B(n_248),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_213),
.B(n_220),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_214),
.A2(n_216),
.B1(n_265),
.B2(n_268),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_153),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_215),
.B(n_219),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_139),
.A2(n_142),
.B1(n_167),
.B2(n_98),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_217),
.A2(n_230),
.B1(n_236),
.B2(n_271),
.Y(n_287)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_218),
.Y(n_325)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_222),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_223),
.Y(n_314)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_191),
.A2(n_41),
.B(n_38),
.C(n_26),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_225),
.B(n_243),
.Y(n_301)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_227),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx3_ASAP7_75t_SL g330 ( 
.A(n_228),
.Y(n_330)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_229),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_160),
.A2(n_73),
.B1(n_65),
.B2(n_66),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_191),
.A2(n_95),
.B1(n_75),
.B2(n_89),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_231),
.A2(n_233),
.B1(n_245),
.B2(n_171),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_153),
.A2(n_71),
.B1(n_110),
.B2(n_106),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_128),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_238),
.B(n_257),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_135),
.Y(n_239)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_127),
.Y(n_240)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_157),
.Y(n_242)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_194),
.B1(n_200),
.B2(n_178),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_128),
.B(n_186),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_246),
.B(n_258),
.Y(n_333)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_127),
.Y(n_247)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_124),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_150),
.Y(n_249)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_154),
.Y(n_254)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_254),
.Y(n_322)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_259),
.Y(n_300)
);

INVx11_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_256),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_196),
.A2(n_22),
.B(n_38),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_124),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_201),
.B(n_17),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_260),
.B(n_261),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_203),
.B(n_52),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_199),
.Y(n_262)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_146),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_264),
.Y(n_302)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_148),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_179),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_166),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_269),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_143),
.B(n_52),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_267),
.B(n_273),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_197),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_174),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_270),
.A2(n_272),
.B1(n_195),
.B2(n_163),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_151),
.A2(n_119),
.B1(n_117),
.B2(n_111),
.Y(n_271)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_163),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_184),
.B(n_41),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_129),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_275),
.Y(n_319)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_282),
.A2(n_289),
.B1(n_304),
.B2(n_312),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_205),
.C(n_215),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_285),
.B(n_327),
.C(n_270),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_216),
.A2(n_189),
.B1(n_126),
.B2(n_195),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_208),
.A2(n_147),
.B1(n_138),
.B2(n_167),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_226),
.B(n_126),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_306),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_225),
.B(n_175),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_205),
.A2(n_161),
.B1(n_155),
.B2(n_181),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_307),
.A2(n_145),
.B1(n_272),
.B2(n_229),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_256),
.A2(n_213),
.B(n_206),
.C(n_258),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_310),
.A2(n_28),
.B(n_223),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_230),
.A2(n_183),
.B1(n_175),
.B2(n_140),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_209),
.B(n_251),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_329),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_244),
.B(n_185),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_320),
.B(n_192),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_211),
.A2(n_144),
.B1(n_164),
.B2(n_149),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_326),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_232),
.B(n_137),
.C(n_183),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_235),
.B(n_50),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_236),
.B(n_50),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_331),
.B(n_332),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_222),
.B(n_32),
.Y(n_332)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_227),
.C(n_249),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_357),
.C(n_361),
.Y(n_395)
);

AND2x4_ASAP7_75t_SL g335 ( 
.A(n_306),
.B(n_211),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_335),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_218),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_336),
.B(n_338),
.Y(n_400)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_221),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_324),
.A2(n_217),
.B1(n_214),
.B2(n_271),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_363),
.B1(n_283),
.B2(n_312),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_342),
.A2(n_369),
.B1(n_330),
.B2(n_289),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_247),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_281),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_345),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_152),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_348),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_165),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_325),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_349),
.B(n_353),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_279),
.A2(n_262),
.B1(n_252),
.B2(n_240),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_350),
.A2(n_330),
.B1(n_325),
.B2(n_280),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_317),
.Y(n_353)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_303),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_354),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_324),
.A2(n_38),
.B(n_22),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_356),
.A2(n_294),
.B(n_332),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_313),
.B(n_263),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_288),
.Y(n_358)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_28),
.B(n_23),
.C(n_210),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_362),
.Y(n_398)
);

INVx13_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_360),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_319),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_293),
.A2(n_268),
.B1(n_265),
.B2(n_241),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_301),
.B(n_264),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_370),
.Y(n_414)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_305),
.B(n_192),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_368),
.A2(n_372),
.B(n_373),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_301),
.B(n_210),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_297),
.Y(n_371)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_277),
.B(n_210),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_277),
.B(n_239),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_284),
.Y(n_374)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_300),
.B(n_237),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_375),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_318),
.B(n_321),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_294),
.B(n_327),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_380),
.A2(n_390),
.B1(n_391),
.B2(n_407),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_381),
.B(n_377),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_323),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_343),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_341),
.A2(n_315),
.B1(n_287),
.B2(n_331),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_385),
.A2(n_388),
.B1(n_405),
.B2(n_411),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_341),
.A2(n_315),
.B1(n_287),
.B2(n_323),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_397),
.A2(n_368),
.B(n_335),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_295),
.C(n_284),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_334),
.C(n_397),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_355),
.A2(n_330),
.B1(n_311),
.B2(n_228),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_340),
.A2(n_280),
.B1(n_309),
.B2(n_296),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_409),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_355),
.A2(n_311),
.B1(n_309),
.B2(n_296),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_337),
.Y(n_412)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_412),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_376),
.C(n_372),
.Y(n_416)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_420),
.C(n_427),
.Y(n_453)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_410),
.Y(n_417)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_395),
.B(n_357),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_418),
.B(n_425),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_419),
.A2(n_444),
.B(n_383),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_362),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_348),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_423),
.B(n_446),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_346),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_353),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_351),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_428),
.B(n_430),
.Y(n_461)
);

NOR2x1_ASAP7_75t_L g479 ( 
.A(n_429),
.B(n_394),
.Y(n_479)
);

A2O1A1O1Ixp25_ASAP7_75t_L g430 ( 
.A1(n_398),
.A2(n_351),
.B(n_346),
.C(n_365),
.D(n_343),
.Y(n_430)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_388),
.A2(n_352),
.B1(n_364),
.B2(n_368),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_439),
.B1(n_441),
.B2(n_450),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_334),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_437),
.C(n_447),
.Y(n_456)
);

INVx13_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_436),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_404),
.B(n_338),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_445),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_391),
.A2(n_373),
.B1(n_336),
.B2(n_370),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_390),
.A2(n_359),
.B1(n_347),
.B2(n_335),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_403),
.Y(n_442)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_442),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_410),
.Y(n_443)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_398),
.B(n_369),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_386),
.B(n_335),
.C(n_322),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_379),
.B(n_360),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_392),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_400),
.B(n_302),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_393),
.C(n_400),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_411),
.A2(n_363),
.B1(n_342),
.B2(n_366),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_436),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_451),
.B(n_455),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_447),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_457),
.A2(n_358),
.B(n_349),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_414),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_459),
.B(n_463),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_431),
.A2(n_414),
.B1(n_407),
.B2(n_415),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_432),
.B1(n_422),
.B2(n_446),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_429),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_421),
.A2(n_405),
.B1(n_415),
.B2(n_393),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_465),
.A2(n_476),
.B1(n_480),
.B2(n_424),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_384),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_418),
.B(n_381),
.C(n_384),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_426),
.C(n_424),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_413),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_473),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_425),
.B(n_413),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_450),
.A2(n_383),
.B1(n_387),
.B2(n_392),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_475),
.A2(n_432),
.B1(n_442),
.B2(n_440),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_412),
.B1(n_378),
.B2(n_389),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_477),
.A2(n_479),
.B(n_422),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_437),
.B(n_444),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_322),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_448),
.A2(n_378),
.B1(n_389),
.B2(n_394),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_430),
.B(n_401),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_481),
.B(n_408),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_453),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_482),
.B(n_490),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_483),
.A2(n_492),
.B1(n_496),
.B2(n_474),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_485),
.A2(n_497),
.B1(n_461),
.B2(n_462),
.Y(n_520)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_486),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_489),
.Y(n_527)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_488),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_477),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_472),
.A2(n_423),
.B(n_426),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_491),
.A2(n_504),
.B(n_479),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_456),
.B(n_402),
.C(n_409),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_493),
.B(n_495),
.C(n_457),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_502),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_402),
.C(n_401),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_465),
.A2(n_433),
.B1(n_417),
.B2(n_443),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_460),
.A2(n_454),
.B1(n_468),
.B2(n_466),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_382),
.Y(n_498)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_498),
.Y(n_526)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_464),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_503),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_458),
.Y(n_501)
);

CKINVDCx14_ASAP7_75t_R g511 ( 
.A(n_501),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_339),
.Y(n_502)
);

INVx13_ASAP7_75t_L g503 ( 
.A(n_471),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_478),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_476),
.B(n_410),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_508),
.Y(n_528)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_474),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_480),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_509),
.A2(n_467),
.B1(n_452),
.B2(n_469),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_513),
.A2(n_519),
.B1(n_522),
.B2(n_532),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_517),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_515),
.A2(n_491),
.B(n_482),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_516),
.B(n_531),
.C(n_502),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_484),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_470),
.C(n_452),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_530),
.Y(n_540)
);

OAI22x1_ASAP7_75t_L g519 ( 
.A1(n_485),
.A2(n_472),
.B1(n_481),
.B2(n_462),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_520),
.A2(n_496),
.B1(n_507),
.B2(n_505),
.Y(n_534)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_521),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_492),
.A2(n_469),
.B1(n_345),
.B2(n_314),
.Y(n_522)
);

NAND2xp67_ASAP7_75t_SL g529 ( 
.A(n_486),
.B(n_490),
.Y(n_529)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_529),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_495),
.B(n_276),
.C(n_308),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_489),
.B(n_276),
.C(n_308),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_509),
.A2(n_314),
.B1(n_281),
.B2(n_290),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_533),
.A2(n_536),
.B(n_530),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_534),
.A2(n_538),
.B1(n_539),
.B2(n_543),
.Y(n_554)
);

OAI321xp33_ASAP7_75t_L g535 ( 
.A1(n_523),
.A2(n_506),
.A3(n_499),
.B1(n_488),
.B2(n_500),
.C(n_508),
.Y(n_535)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_535),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_512),
.A2(n_523),
.B(n_515),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_520),
.A2(n_497),
.B1(n_494),
.B2(n_484),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_526),
.A2(n_498),
.B1(n_504),
.B2(n_503),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_546),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_528),
.A2(n_314),
.B1(n_290),
.B2(n_328),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_528),
.A2(n_328),
.B1(n_325),
.B2(n_291),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_544),
.B(n_548),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_291),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_527),
.B(n_516),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_518),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_529),
.A2(n_360),
.B1(n_354),
.B2(n_316),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_511),
.B(n_298),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_549),
.B(n_278),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_517),
.B(n_316),
.C(n_278),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_551),
.B(n_513),
.C(n_514),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_537),
.A2(n_525),
.B1(n_524),
.B2(n_531),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_552),
.A2(n_558),
.B1(n_559),
.B2(n_544),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_550),
.A2(n_519),
.B(n_524),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_555),
.A2(n_562),
.B(n_563),
.Y(n_570)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_556),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_560),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_522),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_541),
.B(n_510),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_546),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_547),
.B(n_532),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_542),
.B(n_510),
.C(n_298),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_541),
.B(n_354),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_543),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_540),
.B(n_9),
.Y(n_566)
);

AOI221xp5_ASAP7_75t_L g575 ( 
.A1(n_566),
.A2(n_11),
.B1(n_13),
.B2(n_10),
.C(n_7),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_567),
.A2(n_555),
.B(n_557),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_569),
.A2(n_571),
.B(n_565),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_563),
.A2(n_538),
.B(n_539),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_554),
.B(n_545),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_573),
.B(n_578),
.C(n_561),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_577),
.Y(n_587)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_575),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_534),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_576),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_553),
.B(n_551),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_579),
.B(n_10),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_568),
.A2(n_559),
.B(n_564),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_582),
.A2(n_13),
.B(n_3),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_583),
.B(n_586),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_584),
.B(n_585),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_572),
.B(n_560),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_572),
.B(n_21),
.C(n_3),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_588),
.B(n_589),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_576),
.B(n_13),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_581),
.A2(n_570),
.B(n_573),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_590),
.B(n_594),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_587),
.B(n_578),
.Y(n_591)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_591),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_581),
.B(n_574),
.C(n_579),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_2),
.C(n_4),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_SL g597 ( 
.A1(n_592),
.A2(n_580),
.B(n_588),
.C(n_6),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_597),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_600),
.B(n_2),
.Y(n_602)
);

A2O1A1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_602),
.A2(n_598),
.B(n_599),
.C(n_6),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_603),
.B(n_601),
.C(n_4),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_604),
.B(n_595),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_605),
.A2(n_593),
.B1(n_21),
.B2(n_4),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_606),
.A2(n_2),
.B(n_4),
.Y(n_607)
);


endmodule