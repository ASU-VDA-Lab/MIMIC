module fake_aes_11908_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_7), .B(n_8), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_2), .B(n_9), .Y(n_12) );
OAI22xp5_ASAP7_75t_L g13 ( .A1(n_4), .A2(n_8), .B1(n_5), .B2(n_0), .Y(n_13) );
AND2x6_ASAP7_75t_L g14 ( .A(n_7), .B(n_10), .Y(n_14) );
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
NAND2x1_ASAP7_75t_L g17 ( .A(n_1), .B(n_2), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_15), .B(n_0), .Y(n_18) );
AOI22xp33_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_12), .B(n_1), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_12), .B1(n_14), .B2(n_17), .Y(n_22) );
AO21x2_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_11), .B(n_18), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_18), .B(n_17), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_24), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_22), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_13), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_19), .B1(n_12), .B2(n_14), .Y(n_31) );
NAND2xp33_ASAP7_75t_L g32 ( .A(n_29), .B(n_14), .Y(n_32) );
AOI21xp5_ASAP7_75t_L g33 ( .A1(n_29), .A2(n_20), .B(n_19), .Y(n_33) );
AOI222xp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_14), .B1(n_3), .B2(n_5), .C1(n_6), .C2(n_9), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
OAI211xp5_ASAP7_75t_SL g36 ( .A1(n_31), .A2(n_14), .B(n_6), .C(n_10), .Y(n_36) );
AO21x2_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_14), .B(n_4), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
AOI22xp5_ASAP7_75t_SL g39 ( .A1(n_38), .A2(n_34), .B1(n_36), .B2(n_37), .Y(n_39) );
AOI21xp33_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_37), .B(n_38), .Y(n_40) );
endmodule