module fake_netlist_5_996_n_1937 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1937);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1937;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1735;
wire n_1697;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_41),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_75),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_132),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_104),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_97),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_37),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_118),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_26),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_4),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_24),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_4),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_62),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_35),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_13),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_90),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_88),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_30),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_113),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_122),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_36),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_82),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_102),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_73),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_16),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_49),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_92),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_81),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_108),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_41),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_154),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_14),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_18),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_49),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_101),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

INVxp33_ASAP7_75t_R g224 ( 
.A(n_91),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_66),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_110),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_71),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_151),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_72),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_17),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_125),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_14),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_15),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_17),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_20),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_109),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_69),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_42),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_83),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_140),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_145),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_147),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_127),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_149),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_148),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_169),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_85),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_172),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_70),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_131),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_146),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_123),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_124),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_116),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_51),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_67),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_164),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_107),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_58),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_139),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_42),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_120),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_141),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_143),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_100),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_5),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_19),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_133),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_115),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_43),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_161),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_78),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_155),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_29),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_111),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_52),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_157),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_21),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_8),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_34),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_30),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_129),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_60),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_152),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_15),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_23),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_128),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_32),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_52),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_45),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_74),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_1),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_59),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_117),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_98),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_94),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_99),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_22),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_34),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_79),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_22),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_6),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_16),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_44),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_137),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_126),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_40),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_171),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_39),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_93),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_27),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_11),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_44),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_6),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_114),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_28),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_138),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_54),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_46),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_9),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_33),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_55),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_153),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_54),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_130),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_76),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_20),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_80),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_19),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_32),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_37),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_50),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_64),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_204),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_241),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_179),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_207),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_176),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_182),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_300),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_267),
.B(n_0),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_208),
.Y(n_358)
);

INVxp33_ASAP7_75t_SL g359 ( 
.A(n_181),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_241),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_177),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_241),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_178),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_297),
.B(n_0),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_241),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_185),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_180),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_186),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_190),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_267),
.B(n_1),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_297),
.B(n_2),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_242),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_329),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_300),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_289),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_191),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_184),
.B(n_2),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_293),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_298),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_228),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_194),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_293),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_195),
.Y(n_389)
);

BUFx2_ASAP7_75t_SL g390 ( 
.A(n_231),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_187),
.B(n_3),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_298),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_197),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_251),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_199),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_297),
.B(n_7),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_259),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_262),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_269),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_192),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_232),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_285),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_184),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_234),
.B(n_7),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_189),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_189),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_187),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_232),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_210),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_312),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_210),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_216),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_200),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_216),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_201),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_183),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_212),
.B(n_9),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_302),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_237),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_237),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_256),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_205),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_272),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_193),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_256),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_206),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_211),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_268),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_232),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_390),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_349),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_349),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_365),
.B(n_212),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_376),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_349),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_375),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_357),
.B(n_217),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_365),
.B(n_290),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_351),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_360),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_385),
.B(n_214),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_356),
.A2(n_209),
.B1(n_317),
.B2(n_175),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_405),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_188),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_417),
.B(n_215),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_360),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_362),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_188),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_362),
.Y(n_465)
);

OR2x6_ASAP7_75t_L g466 ( 
.A(n_373),
.B(n_290),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_366),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_348),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_367),
.Y(n_470)
);

CKINVDCx6p67_ASAP7_75t_R g471 ( 
.A(n_430),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_402),
.B(n_384),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_367),
.Y(n_473)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_377),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_378),
.B(n_222),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_378),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_379),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_373),
.B(n_311),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_408),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_382),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_402),
.B(n_198),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_372),
.B(n_272),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_R g492 ( 
.A(n_359),
.B(n_368),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_396),
.B(n_198),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_391),
.B(n_226),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_396),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_397),
.B(n_311),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_404),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_423),
.B(n_227),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_407),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_202),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_356),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_383),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_202),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_416),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_441),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_441),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_441),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_440),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_441),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_472),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_440),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_441),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_446),
.B(n_431),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_440),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_451),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_449),
.B(n_430),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_511),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_469),
.B(n_374),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_449),
.A2(n_266),
.B1(n_425),
.B2(n_305),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_472),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_479),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_452),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_471),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_469),
.B(n_416),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_505),
.A2(n_496),
.B1(n_511),
.B2(n_445),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_472),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_479),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_479),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_505),
.A2(n_411),
.B1(n_383),
.B2(n_234),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_446),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_505),
.B(n_225),
.C(n_218),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_477),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_511),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_438),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_453),
.B(n_354),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_438),
.B(n_361),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_477),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_479),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_513),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_446),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_465),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_465),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_441),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_511),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_441),
.Y(n_561)
);

BUFx4f_ASAP7_75t_L g562 ( 
.A(n_496),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_513),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_437),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_454),
.B(n_352),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_441),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_453),
.B(n_364),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_465),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_489),
.B(n_369),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_489),
.B(n_370),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_468),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_496),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_455),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_437),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_468),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_437),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_509),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_442),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_442),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_455),
.Y(n_585)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_511),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_442),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_448),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_496),
.B(n_204),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_464),
.B(n_371),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_511),
.A2(n_420),
.B1(n_422),
.B2(n_433),
.Y(n_592)
);

AND2x2_ASAP7_75t_SL g593 ( 
.A(n_496),
.B(n_204),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_457),
.B(n_381),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_509),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_457),
.B(n_387),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_455),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_505),
.B(n_225),
.C(n_218),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_463),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_444),
.Y(n_602)
);

INVxp33_ASAP7_75t_SL g603 ( 
.A(n_454),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_444),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_463),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_482),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_496),
.B(n_204),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_448),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_482),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_505),
.A2(n_274),
.B1(n_292),
.B2(n_303),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_462),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_444),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_458),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_494),
.B(n_389),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_458),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_494),
.B(n_393),
.Y(n_617)
);

AND2x6_ASAP7_75t_L g618 ( 
.A(n_505),
.B(n_204),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_463),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_458),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_461),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_473),
.Y(n_622)
);

AO21x2_ASAP7_75t_L g623 ( 
.A1(n_502),
.A2(n_238),
.B(n_233),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_445),
.A2(n_450),
.B1(n_466),
.B2(n_456),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_464),
.B(n_395),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_462),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_473),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_502),
.B(n_469),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_487),
.B(n_429),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_480),
.B(n_238),
.C(n_233),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_471),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_456),
.B(n_434),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_460),
.A2(n_299),
.B1(n_275),
.B2(n_263),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_448),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_461),
.Y(n_636)
);

AO22x2_ASAP7_75t_L g637 ( 
.A1(n_445),
.A2(n_303),
.B1(n_287),
.B2(n_292),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_456),
.B(n_353),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_467),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_473),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_467),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_460),
.A2(n_314),
.B1(n_283),
.B2(n_413),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_467),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_470),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_487),
.B(n_276),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_471),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_487),
.B(n_230),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_470),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_475),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_475),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_475),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g653 ( 
.A1(n_445),
.A2(n_244),
.B(n_240),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_481),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_460),
.B(n_436),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_448),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_445),
.B(n_223),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_481),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_507),
.B(n_390),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_448),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_493),
.B(n_418),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_473),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_481),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_450),
.B(n_272),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_484),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_547),
.B(n_450),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_555),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_562),
.B(n_624),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_555),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_562),
.B(n_450),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_520),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_549),
.Y(n_672)
);

AND2x6_ASAP7_75t_SL g673 ( 
.A(n_572),
.B(n_268),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_565),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_612),
.B(n_355),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_553),
.B(n_450),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_556),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_520),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_562),
.A2(n_466),
.B(n_450),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_593),
.A2(n_466),
.B1(n_480),
.B2(n_512),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_586),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_565),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_566),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_520),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_523),
.B(n_512),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_523),
.B(n_599),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_617),
.B(n_507),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_618),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_539),
.B(n_223),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_628),
.B(n_507),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_576),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_545),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_593),
.A2(n_615),
.B1(n_586),
.B2(n_529),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_612),
.B(n_626),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_541),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_541),
.B(n_507),
.Y(n_696)
);

OAI21xp33_ASAP7_75t_L g697 ( 
.A1(n_533),
.A2(n_274),
.B(n_271),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_541),
.B(n_507),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_593),
.B(n_507),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_529),
.A2(n_512),
.B(n_466),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_534),
.B(n_510),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_534),
.B(n_510),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_576),
.B(n_223),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_566),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_545),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_526),
.B(n_358),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_551),
.B(n_363),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_570),
.B(n_510),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_576),
.B(n_548),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_626),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_576),
.B(n_223),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_623),
.A2(n_466),
.B1(n_512),
.B2(n_510),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_601),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_595),
.B(n_510),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_548),
.B(n_223),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_598),
.B(n_510),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_645),
.A2(n_633),
.B(n_630),
.C(n_531),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_620),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_560),
.B(n_512),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_620),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_R g721 ( 
.A(n_537),
.B(n_492),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_560),
.B(n_577),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_577),
.B(n_512),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_577),
.B(n_243),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_531),
.B(n_386),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_601),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_601),
.B(n_466),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_605),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_655),
.B(n_394),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_605),
.B(n_466),
.Y(n_730)
);

INVx8_ASAP7_75t_L g731 ( 
.A(n_618),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_659),
.B(n_245),
.Y(n_732)
);

INVxp33_ASAP7_75t_L g733 ( 
.A(n_578),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_605),
.B(n_466),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_619),
.B(n_490),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_538),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_619),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_552),
.B(n_590),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_621),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_619),
.B(n_246),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_538),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_573),
.A2(n_492),
.B1(n_399),
.B2(n_398),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_532),
.B(n_248),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_661),
.B(n_490),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_621),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_623),
.A2(n_296),
.B1(n_244),
.B2(n_247),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_537),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_592),
.B(n_493),
.C(n_203),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_625),
.B(n_638),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_589),
.B(n_240),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_525),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_578),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_586),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_586),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_544),
.A2(n_401),
.B1(n_406),
.B2(n_288),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_532),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_525),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_585),
.B(n_224),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_585),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_661),
.B(n_493),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_642),
.B(n_219),
.C(n_196),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_533),
.B(n_220),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_532),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_611),
.B(n_229),
.C(n_221),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_527),
.B(n_530),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_582),
.B(n_342),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_629),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_629),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_644),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_527),
.B(n_490),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_530),
.B(n_490),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_532),
.B(n_250),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_532),
.B(n_253),
.Y(n_773)
);

AOI22x1_ASAP7_75t_L g774 ( 
.A1(n_543),
.A2(n_348),
.B1(n_264),
.B2(n_260),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_664),
.B(n_235),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_543),
.B(n_490),
.Y(n_776)
);

NAND2x1_ASAP7_75t_L g777 ( 
.A(n_515),
.B(n_514),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_567),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_634),
.B(n_418),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_648),
.B(n_490),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_567),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_644),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_597),
.B(n_236),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_632),
.B(n_342),
.Y(n_784)
);

NAND3xp33_ASAP7_75t_L g785 ( 
.A(n_631),
.B(n_252),
.C(n_239),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_579),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_579),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_516),
.B(n_499),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_535),
.B(n_257),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_652),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_535),
.B(n_258),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_535),
.B(n_261),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_623),
.B(n_270),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_535),
.B(n_278),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_632),
.Y(n_795)
);

AND3x1_ASAP7_75t_L g796 ( 
.A(n_603),
.B(n_280),
.C(n_271),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_581),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_535),
.B(n_265),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_542),
.B(n_279),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_516),
.B(n_499),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_542),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_542),
.B(n_291),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_524),
.B(n_499),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_342),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_542),
.B(n_294),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_637),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_542),
.B(n_295),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_524),
.B(n_499),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_569),
.A2(n_459),
.B(n_447),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_581),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_554),
.B(n_273),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_554),
.B(n_277),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_652),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_554),
.B(n_281),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_554),
.B(n_301),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_554),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_583),
.B(n_499),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_583),
.B(n_304),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_584),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_584),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_587),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_587),
.B(n_307),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_637),
.B(n_247),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_637),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_637),
.A2(n_338),
.B1(n_282),
.B2(n_284),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_647),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_602),
.B(n_508),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_602),
.B(n_313),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_561),
.B(n_308),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_604),
.B(n_316),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_631),
.A2(n_315),
.B1(n_343),
.B2(n_341),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_561),
.B(n_309),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_604),
.B(n_318),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_613),
.B(n_508),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_613),
.B(n_614),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_546),
.A2(n_327),
.B(n_280),
.C(n_287),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_762),
.A2(n_546),
.B(n_600),
.C(n_327),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_721),
.Y(n_838)
);

O2A1O1Ixp5_ASAP7_75t_L g839 ( 
.A1(n_703),
.A2(n_653),
.B(n_600),
.C(n_521),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_670),
.A2(n_515),
.B(n_518),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_SL g841 ( 
.A1(n_729),
.A2(n_568),
.B1(n_319),
.B2(n_337),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_670),
.A2(n_515),
.B(n_518),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_733),
.B(n_614),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_668),
.B(n_561),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_679),
.A2(n_515),
.B(n_521),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_666),
.B(n_676),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_668),
.B(n_561),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_728),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_722),
.A2(n_636),
.B(n_616),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_728),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_667),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_667),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_669),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_747),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_722),
.A2(n_723),
.B(n_719),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_754),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_669),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_793),
.A2(n_636),
.B(n_616),
.C(n_639),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_723),
.A2(n_640),
.B(n_622),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_836),
.A2(n_639),
.B(n_641),
.C(n_643),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_719),
.A2(n_640),
.B(n_622),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_795),
.B(n_310),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_674),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_736),
.B(n_419),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_760),
.B(n_641),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_741),
.B(n_419),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_671),
.B(n_643),
.Y(n_867)
);

NOR2x1p5_ASAP7_75t_SL g868 ( 
.A(n_718),
.B(n_653),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_678),
.B(n_646),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_693),
.A2(n_640),
.B(n_622),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_672),
.B(n_568),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_684),
.B(n_646),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_686),
.B(n_421),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_752),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_717),
.A2(n_346),
.B(n_328),
.C(n_324),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_677),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_780),
.A2(n_662),
.B(n_517),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_700),
.A2(n_662),
.B(n_517),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_738),
.A2(n_608),
.B1(n_589),
.B2(n_618),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_708),
.B(n_563),
.Y(n_880)
);

O2A1O1Ixp5_ASAP7_75t_L g881 ( 
.A1(n_703),
.A2(n_650),
.B(n_649),
.C(n_651),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_695),
.B(n_649),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_692),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_727),
.A2(n_662),
.B(n_517),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_755),
.A2(n_749),
.B(n_775),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_733),
.B(n_650),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_711),
.A2(n_654),
.B(n_651),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_714),
.B(n_563),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_730),
.A2(n_662),
.B(n_517),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_705),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_734),
.A2(n_519),
.B(n_514),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_766),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_694),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_682),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_682),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_689),
.A2(n_618),
.B1(n_589),
.B2(n_608),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_687),
.A2(n_654),
.B1(n_663),
.B2(n_658),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_709),
.A2(n_519),
.B(n_514),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_683),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_710),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_699),
.A2(n_663),
.B(n_658),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_707),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_713),
.B(n_514),
.Y(n_903)
);

OAI21xp33_ASAP7_75t_L g904 ( 
.A1(n_697),
.A2(n_326),
.B(n_322),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_709),
.A2(n_559),
.B(n_519),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_683),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_704),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_725),
.B(n_421),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_716),
.B(n_563),
.Y(n_909)
);

AOI21x1_ASAP7_75t_L g910 ( 
.A1(n_711),
.A2(n_536),
.B(n_528),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_675),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_826),
.Y(n_912)
);

O2A1O1Ixp5_ASAP7_75t_L g913 ( 
.A1(n_732),
.A2(n_635),
.B(n_660),
.C(n_609),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_748),
.A2(n_589),
.B1(n_608),
.B2(n_618),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_754),
.B(n_426),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_704),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_690),
.A2(n_559),
.B(n_519),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_836),
.A2(n_249),
.B(n_254),
.C(n_340),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_696),
.A2(n_698),
.B(n_744),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_735),
.A2(n_559),
.B(n_563),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_726),
.B(n_559),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_737),
.B(n_589),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_701),
.A2(n_563),
.B(n_660),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_702),
.A2(n_594),
.B(n_660),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_680),
.B(n_588),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_759),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_806),
.A2(n_324),
.B(n_328),
.C(n_346),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_756),
.A2(n_594),
.B(n_660),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_824),
.A2(n_689),
.B(n_685),
.C(n_779),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_756),
.A2(n_594),
.B(n_588),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_770),
.A2(n_665),
.B(n_557),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_691),
.B(n_588),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_756),
.A2(n_594),
.B(n_588),
.Y(n_933)
);

INVx5_ASAP7_75t_L g934 ( 
.A(n_688),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_778),
.B(n_589),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_781),
.A2(n_340),
.B(n_254),
.C(n_255),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_786),
.B(n_589),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_718),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_742),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_787),
.B(n_608),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_732),
.A2(n_288),
.B(n_286),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_777),
.A2(n_656),
.B(n_635),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_783),
.B(n_426),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_746),
.A2(n_249),
.B1(n_330),
.B2(n_306),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_823),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_784),
.B(n_427),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_797),
.B(n_608),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_691),
.A2(n_656),
.B(n_635),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_706),
.B(n_810),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_691),
.A2(n_656),
.B(n_635),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_819),
.A2(n_255),
.B(n_260),
.C(n_264),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_820),
.Y(n_952)
);

BUFx4f_ASAP7_75t_SL g953 ( 
.A(n_743),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_720),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_765),
.A2(n_656),
.B(n_609),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_821),
.B(n_608),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_804),
.B(n_427),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_835),
.A2(n_609),
.B(n_522),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_724),
.A2(n_609),
.B(n_522),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_724),
.A2(n_681),
.B(n_801),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_720),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_751),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_739),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_712),
.A2(n_757),
.B1(n_681),
.B2(n_825),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_771),
.A2(n_665),
.B(n_575),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_763),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_681),
.A2(n_522),
.B(n_459),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_818),
.B(n_822),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_758),
.Y(n_969)
);

NOR2xp67_ASAP7_75t_L g970 ( 
.A(n_785),
.B(n_428),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_801),
.A2(n_522),
.B(n_459),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_740),
.A2(n_608),
.B1(n_618),
.B2(n_657),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_776),
.A2(n_800),
.B(n_788),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_816),
.A2(n_522),
.B(n_459),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_739),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_828),
.B(n_618),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_673),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_763),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_830),
.B(n_596),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_816),
.A2(n_522),
.B(n_459),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_833),
.A2(n_296),
.B(n_286),
.C(n_306),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_794),
.B(n_596),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_803),
.A2(n_459),
.B(n_627),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_817),
.A2(n_550),
.B(n_528),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_753),
.B(n_428),
.Y(n_985)
);

OAI21xp33_ASAP7_75t_L g986 ( 
.A1(n_761),
.A2(n_333),
.B(n_334),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_808),
.A2(n_459),
.B(n_627),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_745),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_764),
.B(n_330),
.C(n_335),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_799),
.B(n_606),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_796),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_802),
.B(n_606),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_827),
.A2(n_574),
.B(n_536),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_L g994 ( 
.A(n_740),
.B(n_336),
.C(n_339),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_823),
.A2(n_558),
.B(n_540),
.C(n_550),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_763),
.Y(n_996)
);

NOR2xp67_ASAP7_75t_L g997 ( 
.A(n_831),
.B(n_432),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_823),
.A2(n_321),
.B1(n_323),
.B2(n_325),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_823),
.B(n_344),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_753),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_805),
.B(n_432),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_745),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_767),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_807),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_753),
.A2(n_320),
.B1(n_332),
.B2(n_574),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_815),
.B(n_607),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_774),
.A2(n_657),
.B1(n_610),
.B2(n_607),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_767),
.B(n_610),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_768),
.B(n_540),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_763),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_768),
.B(n_769),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_769),
.B(n_557),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_782),
.B(n_558),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_782),
.B(n_564),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_790),
.B(n_564),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_790),
.B(n_571),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_829),
.A2(n_627),
.B(n_571),
.Y(n_1017)
);

BUFx4f_ASAP7_75t_L g1018 ( 
.A(n_688),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_813),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_834),
.A2(n_591),
.B(n_580),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_829),
.A2(n_627),
.B(n_575),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_813),
.B(n_580),
.Y(n_1022)
);

OAI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_743),
.A2(n_435),
.B(n_814),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_772),
.A2(n_591),
.B(n_508),
.C(n_491),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_772),
.B(n_773),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_773),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_876),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_846),
.A2(n_731),
.B(n_688),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_874),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_848),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_996),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_982),
.A2(n_731),
.B(n_688),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_996),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_996),
.Y(n_1034)
);

AO21x1_ASAP7_75t_L g1035 ( 
.A1(n_968),
.A2(n_832),
.B(n_814),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_885),
.A2(n_949),
.B(n_981),
.C(n_892),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_990),
.A2(n_731),
.B(n_832),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_949),
.A2(n_657),
.B1(n_750),
.B2(n_812),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_851),
.Y(n_1039)
);

OAI21xp33_ASAP7_75t_L g1040 ( 
.A1(n_943),
.A2(n_812),
.B(n_811),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1001),
.B(n_789),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_853),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_883),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_853),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_964),
.A2(n_657),
.B1(n_750),
.B2(n_798),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_996),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_992),
.A2(n_731),
.B(n_791),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_857),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_857),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1006),
.A2(n_811),
.B(n_789),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_981),
.A2(n_798),
.B(n_792),
.C(n_791),
.Y(n_1051)
);

BUFx2_ASAP7_75t_SL g1052 ( 
.A(n_890),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_890),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_850),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_1025),
.A2(n_929),
.B(n_855),
.C(n_1023),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_939),
.A2(n_1025),
.B1(n_865),
.B2(n_989),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_994),
.A2(n_792),
.B(n_715),
.C(n_809),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1004),
.B(n_715),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_902),
.B(n_12),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_854),
.B(n_657),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_966),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_848),
.A2(n_508),
.B1(n_491),
.B2(n_504),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_893),
.B(n_900),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_926),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_911),
.B(n_491),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_875),
.A2(n_941),
.A3(n_897),
.B(n_837),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_966),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_994),
.A2(n_657),
.B1(n_497),
.B2(n_504),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_858),
.A2(n_999),
.B(n_1026),
.C(n_843),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_SL g1070 ( 
.A(n_841),
.B(n_986),
.C(n_999),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_978),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_843),
.B(n_497),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_863),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_991),
.Y(n_1074)
);

INVx4_ASAP7_75t_L g1075 ( 
.A(n_850),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_953),
.B(n_497),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_989),
.A2(n_657),
.B1(n_501),
.B2(n_504),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_873),
.B(n_435),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_945),
.B(n_501),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_946),
.A2(n_501),
.B1(n_484),
.B2(n_506),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_969),
.B(n_12),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_886),
.B(n_483),
.Y(n_1082)
);

AO32x2_ASAP7_75t_L g1083 ( 
.A1(n_944),
.A2(n_13),
.A3(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_886),
.B(n_483),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_845),
.A2(n_439),
.B(n_443),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_908),
.B(n_957),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_952),
.B(n_483),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_927),
.A2(n_506),
.B(n_500),
.C(n_498),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_927),
.A2(n_506),
.B(n_500),
.C(n_498),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_925),
.A2(n_476),
.B1(n_506),
.B2(n_500),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_912),
.B(n_486),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_925),
.A2(n_476),
.B1(n_500),
.B2(n_498),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_862),
.B(n_25),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_978),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_838),
.B(n_96),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_852),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1018),
.A2(n_476),
.B1(n_498),
.B2(n_495),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_962),
.B(n_483),
.Y(n_1098)
);

INVxp67_ASAP7_75t_SL g1099 ( 
.A(n_856),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1018),
.A2(n_476),
.B1(n_495),
.B2(n_486),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_864),
.B(n_483),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_953),
.B(n_485),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_837),
.A2(n_495),
.B(n_486),
.C(n_485),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_864),
.B(n_483),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_875),
.A2(n_495),
.B(n_484),
.C(n_486),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_871),
.B(n_485),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_866),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_960),
.A2(n_439),
.B(n_443),
.Y(n_1108)
);

BUFx4f_ASAP7_75t_L g1109 ( 
.A(n_977),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_866),
.B(n_485),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_945),
.A2(n_503),
.B1(n_488),
.B2(n_484),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_878),
.A2(n_439),
.B(n_443),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_915),
.B(n_476),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1010),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_915),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_894),
.Y(n_1116)
);

OR2x6_ASAP7_75t_L g1117 ( 
.A(n_995),
.B(n_503),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_997),
.A2(n_476),
.B(n_443),
.C(n_447),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_985),
.A2(n_488),
.B1(n_503),
.B2(n_448),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_895),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_919),
.B(n_503),
.Y(n_1121)
);

AO32x1_ASAP7_75t_L g1122 ( 
.A1(n_907),
.A2(n_439),
.A3(n_447),
.B1(n_27),
.B2(n_29),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_976),
.A2(n_447),
.B(n_488),
.C(n_503),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_936),
.A2(n_25),
.B(n_26),
.C(n_31),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_SL g1125 ( 
.A(n_934),
.B(n_448),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_965),
.A2(n_448),
.B(n_134),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_859),
.A2(n_474),
.B(n_478),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_916),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_899),
.B(n_503),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_861),
.A2(n_474),
.B(n_478),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_844),
.A2(n_488),
.B1(n_503),
.B2(n_478),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_906),
.B(n_503),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_954),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_904),
.B(n_31),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_979),
.A2(n_503),
.B1(n_488),
.B2(n_478),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_985),
.B(n_867),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_856),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_934),
.B(n_488),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_934),
.B(n_488),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_840),
.A2(n_474),
.B(n_478),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_869),
.B(n_488),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1010),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_842),
.A2(n_474),
.B(n_478),
.Y(n_1143)
);

AOI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_998),
.A2(n_35),
.B(n_36),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_844),
.B(n_38),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_847),
.B(n_39),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_847),
.A2(n_488),
.B1(n_478),
.B2(n_473),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_970),
.B(n_478),
.C(n_473),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_872),
.B(n_882),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_954),
.B(n_473),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_961),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_938),
.A2(n_473),
.B1(n_474),
.B2(n_84),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_961),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_975),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_963),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_934),
.A2(n_474),
.B(n_473),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_879),
.A2(n_474),
.B1(n_77),
.B2(n_86),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_963),
.B(n_40),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1000),
.B(n_474),
.Y(n_1159)
);

AOI22x1_ASAP7_75t_L g1160 ( 
.A1(n_891),
.A2(n_65),
.B1(n_158),
.B2(n_144),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_SL g1161 ( 
.A(n_918),
.B(n_45),
.C(n_46),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_936),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1002),
.B(n_1003),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1000),
.B(n_988),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_988),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1019),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1019),
.A2(n_87),
.B1(n_142),
.B2(n_135),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_903),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_951),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1011),
.B(n_47),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1008),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_951),
.B(n_47),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1009),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_921),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_880),
.B(n_48),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_880),
.A2(n_162),
.B(n_121),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1013),
.B(n_48),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_888),
.A2(n_112),
.B(n_105),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_935),
.A2(n_103),
.B1(n_89),
.B2(n_53),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1012),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1015),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_860),
.A2(n_50),
.B(n_51),
.C(n_53),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_849),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1016),
.Y(n_1184)
);

NAND2x1p5_ASAP7_75t_L g1185 ( 
.A(n_932),
.B(n_55),
.Y(n_1185)
);

AO21x2_ASAP7_75t_L g1186 ( 
.A1(n_1055),
.A2(n_870),
.B(n_901),
.Y(n_1186)
);

AOI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1050),
.A2(n_888),
.B(n_909),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1056),
.A2(n_1005),
.B1(n_914),
.B2(n_972),
.Y(n_1188)
);

OAI22x1_ASAP7_75t_L g1189 ( 
.A1(n_1056),
.A2(n_887),
.B1(n_909),
.B2(n_932),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1115),
.B(n_868),
.Y(n_1190)
);

AO21x1_ASAP7_75t_L g1191 ( 
.A1(n_1036),
.A2(n_1024),
.B(n_889),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_SL g1192 ( 
.A1(n_1182),
.A2(n_940),
.B(n_947),
.C(n_937),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1086),
.A2(n_896),
.B1(n_956),
.B2(n_922),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_SL g1194 ( 
.A(n_1027),
.B(n_1022),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1029),
.B(n_1022),
.Y(n_1195)
);

NAND3x1_ASAP7_75t_L g1196 ( 
.A(n_1059),
.B(n_1093),
.C(n_1081),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1037),
.A2(n_877),
.B(n_884),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1035),
.A2(n_1014),
.A3(n_1013),
.B(n_1021),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1126),
.A2(n_910),
.B(n_905),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1078),
.B(n_1016),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1047),
.A2(n_923),
.B(n_913),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1064),
.B(n_898),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1069),
.A2(n_881),
.B(n_839),
.C(n_984),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1028),
.A2(n_920),
.B(n_917),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1149),
.B(n_1014),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1039),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1043),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1032),
.A2(n_955),
.B(n_950),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1041),
.A2(n_948),
.B(n_924),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1112),
.A2(n_973),
.B(n_928),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1136),
.B(n_1020),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1079),
.B(n_942),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1151),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1074),
.B(n_958),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1107),
.B(n_1076),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1108),
.A2(n_933),
.B(n_930),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1040),
.A2(n_959),
.B(n_993),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1053),
.Y(n_1218)
);

INVx3_ASAP7_75t_SL g1219 ( 
.A(n_1053),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1058),
.A2(n_896),
.B1(n_1007),
.B2(n_931),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1121),
.A2(n_1017),
.B(n_967),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1173),
.B(n_1007),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1052),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1123),
.A2(n_987),
.A3(n_983),
.B(n_974),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1106),
.B(n_56),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1057),
.A2(n_980),
.A3(n_971),
.B(n_58),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1183),
.A2(n_56),
.A3(n_57),
.B(n_1105),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1070),
.A2(n_57),
.B(n_1051),
.C(n_1134),
.Y(n_1228)
);

AO31x2_ASAP7_75t_L g1229 ( 
.A1(n_1175),
.A2(n_1146),
.A3(n_1145),
.B(n_1162),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1049),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1144),
.B(n_1179),
.C(n_1124),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1153),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1053),
.Y(n_1233)
);

AO21x1_ASAP7_75t_L g1234 ( 
.A1(n_1177),
.A2(n_1170),
.B(n_1158),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1045),
.A2(n_1038),
.B(n_1068),
.C(n_1077),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1045),
.A2(n_1038),
.B(n_1077),
.C(n_1169),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1082),
.A2(n_1084),
.B(n_1101),
.Y(n_1237)
);

INVx8_ASAP7_75t_L g1238 ( 
.A(n_1034),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1090),
.A2(n_1092),
.A3(n_1135),
.B(n_1062),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1141),
.A2(n_1117),
.B(n_1139),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1118),
.A2(n_1157),
.A3(n_1125),
.B(n_1100),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1030),
.A2(n_1154),
.B1(n_1099),
.B2(n_1174),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1073),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1054),
.Y(n_1244)
);

AOI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1168),
.A2(n_1104),
.B(n_1091),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1161),
.A2(n_1065),
.B(n_1102),
.C(n_1063),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1072),
.A2(n_1120),
.B1(n_1096),
.B2(n_1116),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1128),
.A2(n_1117),
.B1(n_1075),
.B2(n_1181),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1171),
.B(n_1180),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1117),
.A2(n_1138),
.B(n_1085),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1179),
.B(n_1167),
.C(n_1172),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1054),
.B(n_1075),
.Y(n_1252)
);

INVx5_ASAP7_75t_L g1253 ( 
.A(n_1034),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1097),
.A2(n_1127),
.A3(n_1130),
.B(n_1184),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1163),
.B(n_1079),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1110),
.A2(n_1079),
.B(n_1185),
.C(n_1113),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_1137),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1140),
.A2(n_1143),
.A3(n_1178),
.B(n_1176),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1133),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1060),
.A2(n_1150),
.B(n_1164),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1129),
.A2(n_1132),
.B(n_1156),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1054),
.A2(n_1164),
.B1(n_1137),
.B2(n_1048),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1095),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1103),
.A2(n_1098),
.B(n_1087),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1114),
.Y(n_1265)
);

OAI22x1_ASAP7_75t_L g1266 ( 
.A1(n_1160),
.A2(n_1167),
.B1(n_1044),
.B2(n_1042),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1061),
.A2(n_1067),
.B(n_1071),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1114),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1155),
.B(n_1166),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1165),
.A2(n_1122),
.A3(n_1066),
.B(n_1031),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1080),
.B(n_1094),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1114),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1061),
.A2(n_1094),
.B(n_1071),
.Y(n_1273)
);

BUFx4_ASAP7_75t_SL g1274 ( 
.A(n_1109),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1088),
.A2(n_1089),
.B(n_1147),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1142),
.B(n_1067),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1142),
.B(n_1031),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1159),
.A2(n_1152),
.B(n_1148),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1152),
.A2(n_1080),
.B(n_1122),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1147),
.A2(n_1131),
.B(n_1111),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1131),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1034),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1119),
.A2(n_1066),
.B(n_1033),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1083),
.B(n_1109),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1066),
.A2(n_1033),
.B(n_1122),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1046),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1046),
.B(n_1083),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1083),
.A2(n_1035),
.A3(n_875),
.B(n_1055),
.Y(n_1288)
);

NOR2x1_ASAP7_75t_R g1289 ( 
.A(n_1046),
.B(n_747),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1151),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1039),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1151),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_SL g1293 ( 
.A(n_1070),
.B(n_902),
.C(n_968),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1149),
.B(n_1086),
.Y(n_1294)
);

AO32x2_ASAP7_75t_L g1295 ( 
.A1(n_1090),
.A2(n_944),
.A3(n_964),
.B1(n_806),
.B2(n_824),
.Y(n_1295)
);

INVx5_ASAP7_75t_L g1296 ( 
.A(n_1034),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1055),
.A2(n_968),
.B(n_885),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1055),
.A2(n_846),
.B(n_562),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1096),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1096),
.Y(n_1300)
);

NOR2x1_ASAP7_75t_L g1301 ( 
.A(n_1075),
.B(n_876),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1035),
.A2(n_875),
.A3(n_1055),
.B(n_1123),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1096),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1035),
.A2(n_875),
.A3(n_1055),
.B(n_1123),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1086),
.B(n_725),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1035),
.A2(n_875),
.A3(n_1055),
.B(n_1123),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1086),
.B(n_725),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1054),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1036),
.A2(n_885),
.B(n_968),
.C(n_572),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1039),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1126),
.A2(n_965),
.B(n_1112),
.Y(n_1311)
);

INVxp67_ASAP7_75t_SL g1312 ( 
.A(n_1086),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1027),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1035),
.A2(n_875),
.A3(n_1055),
.B(n_1123),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1055),
.A2(n_846),
.B(n_562),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1055),
.A2(n_846),
.B(n_562),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1115),
.B(n_1079),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1027),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1055),
.A2(n_846),
.B(n_562),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1039),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1151),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1055),
.A2(n_846),
.B(n_562),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1059),
.A2(n_568),
.B(n_729),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1054),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1126),
.A2(n_965),
.B(n_1112),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1055),
.A2(n_846),
.B(n_562),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1151),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1070),
.B(n_721),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1036),
.A2(n_885),
.B(n_968),
.C(n_572),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1035),
.A2(n_875),
.A3(n_1055),
.B(n_1123),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1086),
.B(n_725),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1126),
.A2(n_965),
.B(n_1112),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1055),
.A2(n_875),
.B(n_1123),
.Y(n_1333)
);

AOI221x1_ASAP7_75t_L g1334 ( 
.A1(n_1182),
.A2(n_885),
.B1(n_968),
.B2(n_1144),
.C(n_875),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1055),
.A2(n_875),
.B(n_1123),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1027),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1134),
.A2(n_885),
.B1(n_968),
.B2(n_939),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_SL g1338 ( 
.A1(n_1055),
.A2(n_885),
.B(n_968),
.C(n_1182),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_SL g1339 ( 
.A1(n_1055),
.A2(n_885),
.B(n_968),
.C(n_1182),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1027),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1035),
.A2(n_875),
.A3(n_1055),
.B(n_1123),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1149),
.B(n_1086),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1053),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1027),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1039),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1086),
.B(n_725),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1126),
.A2(n_965),
.B(n_1112),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1055),
.A2(n_846),
.B(n_562),
.Y(n_1348)
);

INVxp67_ASAP7_75t_SL g1349 ( 
.A(n_1205),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1251),
.A2(n_1231),
.B1(n_1297),
.B2(n_1312),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1286),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1336),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1337),
.A2(n_1294),
.B1(n_1342),
.B2(n_1196),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1244),
.Y(n_1354)
);

INVx6_ASAP7_75t_L g1355 ( 
.A(n_1253),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1318),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1309),
.A2(n_1329),
.B1(n_1323),
.B2(n_1236),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1300),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1305),
.B(n_1307),
.Y(n_1359)
);

BUFx10_ASAP7_75t_L g1360 ( 
.A(n_1343),
.Y(n_1360)
);

INVx11_ASAP7_75t_L g1361 ( 
.A(n_1274),
.Y(n_1361)
);

INVx5_ASAP7_75t_L g1362 ( 
.A(n_1238),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1303),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1344),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1213),
.Y(n_1365)
);

BUFx4_ASAP7_75t_SL g1366 ( 
.A(n_1218),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1228),
.A2(n_1235),
.B1(n_1214),
.B2(n_1215),
.Y(n_1367)
);

CKINVDCx6p67_ASAP7_75t_R g1368 ( 
.A(n_1219),
.Y(n_1368)
);

OAI21xp33_ASAP7_75t_L g1369 ( 
.A1(n_1331),
.A2(n_1346),
.B(n_1293),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1213),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1313),
.A2(n_1340),
.B1(n_1255),
.B2(n_1223),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1200),
.A2(n_1207),
.B1(n_1248),
.B2(n_1262),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1233),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1232),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1225),
.B(n_1317),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1284),
.A2(n_1234),
.B1(n_1328),
.B2(n_1245),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1343),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1194),
.A2(n_1195),
.B1(n_1263),
.B2(n_1317),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1188),
.A2(n_1249),
.B1(n_1301),
.B2(n_1271),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1298),
.A2(n_1348),
.B1(n_1326),
.B2(n_1322),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1232),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1343),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1315),
.A2(n_1319),
.B1(n_1316),
.B2(n_1211),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1238),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1244),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1244),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1253),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1229),
.B(n_1272),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1229),
.B(n_1269),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1290),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1292),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1229),
.B(n_1206),
.Y(n_1392)
);

OAI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1334),
.A2(n_1222),
.B1(n_1247),
.B2(n_1281),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1308),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1321),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1186),
.A2(n_1281),
.B1(n_1333),
.B2(n_1335),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1268),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1253),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1308),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1252),
.A2(n_1324),
.B1(n_1242),
.B2(n_1265),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1296),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1321),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1327),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1327),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1324),
.A2(n_1289),
.B1(n_1282),
.B2(n_1190),
.Y(n_1405)
);

BUFx8_ASAP7_75t_L g1406 ( 
.A(n_1190),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1230),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1268),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1279),
.A2(n_1220),
.B1(n_1202),
.B2(n_1320),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1243),
.Y(n_1410)
);

BUFx2_ASAP7_75t_L g1411 ( 
.A(n_1296),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1296),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1333),
.A2(n_1335),
.B1(n_1191),
.B2(n_1237),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1259),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1246),
.B(n_1345),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1291),
.Y(n_1416)
);

CKINVDCx11_ASAP7_75t_R g1417 ( 
.A(n_1310),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1257),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1256),
.A2(n_1240),
.B1(n_1212),
.B2(n_1276),
.Y(n_1419)
);

CKINVDCx6p67_ASAP7_75t_R g1420 ( 
.A(n_1212),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_SL g1421 ( 
.A(n_1277),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1226),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1338),
.B(n_1339),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1287),
.A2(n_1189),
.B1(n_1193),
.B2(n_1266),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1270),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1227),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1278),
.A2(n_1280),
.B1(n_1217),
.B2(n_1209),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1227),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1227),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_SL g1430 ( 
.A(n_1295),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1267),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1270),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1288),
.B(n_1273),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_SL g1434 ( 
.A1(n_1283),
.A2(n_1260),
.B1(n_1250),
.B2(n_1275),
.Y(n_1434)
);

INVx6_ASAP7_75t_L g1435 ( 
.A(n_1226),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1264),
.A2(n_1285),
.B1(n_1201),
.B2(n_1197),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1221),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1203),
.A2(n_1187),
.B1(n_1208),
.B2(n_1204),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1192),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1288),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1295),
.A2(n_1288),
.B1(n_1341),
.B2(n_1330),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1295),
.A2(n_1302),
.B(n_1341),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1302),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1304),
.B(n_1306),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1261),
.A2(n_1216),
.B1(n_1210),
.B2(n_1199),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1304),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1241),
.A2(n_1314),
.B1(n_1341),
.B2(n_1330),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1311),
.A2(n_1347),
.B1(n_1332),
.B2(n_1325),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1241),
.A2(n_1314),
.B1(n_1239),
.B2(n_1198),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1314),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1198),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1254),
.B(n_1258),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1254),
.B(n_1258),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1239),
.A2(n_1241),
.B1(n_1254),
.B2(n_1224),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1224),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1239),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1323),
.A2(n_568),
.B(n_729),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1313),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1299),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1251),
.A2(n_729),
.B1(n_902),
.B2(n_762),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1299),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1337),
.A2(n_885),
.B1(n_968),
.B2(n_1251),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1253),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1337),
.A2(n_885),
.B1(n_968),
.B2(n_1251),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1337),
.A2(n_885),
.B1(n_968),
.B2(n_1251),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1337),
.A2(n_885),
.B1(n_968),
.B2(n_1251),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1337),
.A2(n_885),
.B1(n_968),
.B2(n_1251),
.Y(n_1467)
);

INVx8_ASAP7_75t_L g1468 ( 
.A(n_1238),
.Y(n_1468)
);

BUFx2_ASAP7_75t_SL g1469 ( 
.A(n_1286),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1318),
.Y(n_1470)
);

BUFx4f_ASAP7_75t_SL g1471 ( 
.A(n_1286),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1336),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1337),
.A2(n_885),
.B1(n_968),
.B2(n_1251),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1299),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1253),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1337),
.A2(n_968),
.B1(n_1342),
.B2(n_1294),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1244),
.Y(n_1477)
);

BUFx8_ASAP7_75t_SL g1478 ( 
.A(n_1286),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1205),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1299),
.Y(n_1480)
);

BUFx12f_ASAP7_75t_L g1481 ( 
.A(n_1318),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1299),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1294),
.A2(n_968),
.B1(n_1093),
.B2(n_489),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1337),
.A2(n_885),
.B1(n_968),
.B2(n_1251),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1337),
.A2(n_968),
.B1(n_1342),
.B2(n_1294),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_SL g1486 ( 
.A(n_1469),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1460),
.A2(n_1466),
.B1(n_1462),
.B2(n_1464),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1388),
.B(n_1440),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1448),
.A2(n_1445),
.B(n_1438),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1478),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1392),
.B(n_1365),
.Y(n_1491)
);

INVx5_ASAP7_75t_L g1492 ( 
.A(n_1439),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1406),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1365),
.B(n_1370),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1389),
.B(n_1444),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1364),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1428),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1375),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1458),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1370),
.B(n_1381),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1381),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1402),
.B(n_1374),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1406),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1418),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1357),
.A2(n_1367),
.B1(n_1353),
.B2(n_1483),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1425),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1456),
.B(n_1451),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1425),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1439),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1462),
.A2(n_1465),
.B(n_1484),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1442),
.A2(n_1436),
.B(n_1380),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1420),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1463),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1432),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1443),
.Y(n_1515)
);

AOI21xp33_ASAP7_75t_L g1516 ( 
.A1(n_1464),
.A2(n_1473),
.B(n_1466),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1476),
.A2(n_1485),
.B1(n_1349),
.B2(n_1479),
.Y(n_1517)
);

A2O1A1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1465),
.A2(n_1484),
.B(n_1473),
.C(n_1467),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_SL g1519 ( 
.A1(n_1423),
.A2(n_1415),
.B(n_1433),
.Y(n_1519)
);

BUFx2_ASAP7_75t_SL g1520 ( 
.A(n_1421),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1446),
.Y(n_1521)
);

NAND2x1_ASAP7_75t_L g1522 ( 
.A(n_1435),
.B(n_1383),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1450),
.B(n_1424),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1435),
.Y(n_1525)
);

INVx4_ASAP7_75t_SL g1526 ( 
.A(n_1435),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1405),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1455),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1409),
.A2(n_1453),
.B(n_1452),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1350),
.B(n_1467),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1395),
.B(n_1403),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1393),
.B(n_1376),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1355),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1372),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1404),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1355),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1450),
.B(n_1424),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1371),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1393),
.B(n_1376),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1358),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1449),
.B(n_1422),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1363),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1430),
.Y(n_1543)
);

BUFx4f_ASAP7_75t_SL g1544 ( 
.A(n_1351),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1419),
.Y(n_1545)
);

AO21x2_ASAP7_75t_L g1546 ( 
.A1(n_1409),
.A2(n_1441),
.B(n_1447),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1355),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1459),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1448),
.A2(n_1445),
.B(n_1436),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1441),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1461),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1380),
.A2(n_1427),
.B(n_1383),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1427),
.A2(n_1396),
.B(n_1454),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1396),
.B(n_1454),
.Y(n_1554)
);

AO21x2_ASAP7_75t_L g1555 ( 
.A1(n_1379),
.A2(n_1369),
.B(n_1480),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1359),
.B(n_1413),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1413),
.A2(n_1482),
.B(n_1474),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1457),
.A2(n_1378),
.B(n_1434),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1387),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1397),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1437),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1429),
.A2(n_1426),
.B1(n_1417),
.B2(n_1421),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1431),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1416),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1373),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1426),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1407),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1463),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1410),
.B(n_1414),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1398),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1356),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1382),
.B(n_1354),
.Y(n_1572)
);

CKINVDCx9p33_ASAP7_75t_R g1573 ( 
.A(n_1470),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1411),
.A2(n_1408),
.B(n_1386),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1400),
.A2(n_1398),
.B(n_1401),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1387),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1387),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1549),
.A2(n_1412),
.B(n_1475),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1505),
.A2(n_1481),
.B1(n_1368),
.B2(n_1471),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_L g1580 ( 
.A(n_1487),
.B(n_1394),
.C(n_1362),
.Y(n_1580)
);

BUFx4f_ASAP7_75t_L g1581 ( 
.A(n_1509),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1518),
.A2(n_1471),
.B1(n_1412),
.B2(n_1475),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1544),
.B(n_1481),
.Y(n_1583)
);

OA21x2_ASAP7_75t_L g1584 ( 
.A1(n_1549),
.A2(n_1475),
.B(n_1412),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1540),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1510),
.A2(n_1401),
.B(n_1477),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1495),
.B(n_1477),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1561),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1510),
.A2(n_1362),
.B(n_1468),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1498),
.B(n_1360),
.Y(n_1590)
);

AO22x2_ASAP7_75t_L g1591 ( 
.A1(n_1558),
.A2(n_1384),
.B1(n_1394),
.B2(n_1366),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1516),
.A2(n_1362),
.B(n_1399),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1491),
.B(n_1362),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1566),
.B(n_1360),
.Y(n_1594)
);

CKINVDCx14_ASAP7_75t_R g1595 ( 
.A(n_1490),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1542),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1543),
.B(n_1468),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1548),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1502),
.B(n_1377),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1522),
.A2(n_1468),
.B(n_1385),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1543),
.B(n_1352),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1516),
.A2(n_1472),
.B1(n_1399),
.B2(n_1377),
.C(n_1385),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1530),
.A2(n_1361),
.B(n_1517),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1491),
.B(n_1561),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1558),
.A2(n_1530),
.B(n_1545),
.C(n_1532),
.Y(n_1605)
);

AOI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1532),
.A2(n_1539),
.B(n_1534),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1535),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1563),
.B(n_1504),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1539),
.B(n_1538),
.C(n_1545),
.Y(n_1609)
);

AOI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1519),
.A2(n_1524),
.B1(n_1537),
.B2(n_1496),
.C(n_1550),
.Y(n_1610)
);

O2A1O1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1519),
.A2(n_1527),
.B(n_1565),
.C(n_1571),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1573),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1488),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1574),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1551),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1493),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1574),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1566),
.B(n_1572),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1560),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1572),
.B(n_1494),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1502),
.B(n_1526),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1486),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1556),
.B(n_1541),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1494),
.B(n_1500),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1499),
.B(n_1527),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1522),
.A2(n_1552),
.B(n_1563),
.Y(n_1626)
);

OR2x6_ASAP7_75t_L g1627 ( 
.A(n_1552),
.B(n_1520),
.Y(n_1627)
);

CKINVDCx6p67_ASAP7_75t_R g1628 ( 
.A(n_1493),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1524),
.A2(n_1537),
.B1(n_1550),
.B2(n_1562),
.C(n_1555),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1563),
.B(n_1501),
.Y(n_1630)
);

AOI22x1_ASAP7_75t_SL g1631 ( 
.A1(n_1576),
.A2(n_1577),
.B1(n_1567),
.B2(n_1513),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1527),
.A2(n_1520),
.B1(n_1555),
.B2(n_1563),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1493),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1541),
.B(n_1523),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1523),
.B(n_1531),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1523),
.Y(n_1636)
);

A2O1A1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1553),
.A2(n_1503),
.B(n_1512),
.C(n_1489),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1553),
.A2(n_1557),
.B(n_1489),
.Y(n_1638)
);

A2O1A1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1503),
.A2(n_1512),
.B(n_1554),
.C(n_1492),
.Y(n_1639)
);

INVx4_ASAP7_75t_L g1640 ( 
.A(n_1512),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1503),
.A2(n_1492),
.B1(n_1509),
.B2(n_1569),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1531),
.Y(n_1642)
);

NAND2x1_ASAP7_75t_L g1643 ( 
.A(n_1574),
.B(n_1570),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1526),
.B(n_1525),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1607),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1638),
.B(n_1511),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1638),
.B(n_1511),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1644),
.Y(n_1649)
);

OAI222xp33_ASAP7_75t_L g1650 ( 
.A1(n_1582),
.A2(n_1554),
.B1(n_1567),
.B2(n_1492),
.C1(n_1564),
.C2(n_1577),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1580),
.A2(n_1555),
.B1(n_1546),
.B2(n_1511),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1636),
.B(n_1546),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1642),
.B(n_1546),
.Y(n_1653)
);

BUFx2_ASAP7_75t_L g1654 ( 
.A(n_1614),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1578),
.B(n_1529),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1578),
.B(n_1529),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1584),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1623),
.B(n_1529),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1588),
.B(n_1604),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1617),
.B(n_1497),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1630),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1617),
.B(n_1528),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1608),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1624),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1508),
.Y(n_1665)
);

BUFx12f_ASAP7_75t_L g1666 ( 
.A(n_1622),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1608),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1585),
.B(n_1515),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1613),
.B(n_1634),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1605),
.A2(n_1492),
.B1(n_1509),
.B2(n_1574),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1626),
.B(n_1515),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1596),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1635),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1643),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1620),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1598),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1587),
.Y(n_1677)
);

AO21x2_ASAP7_75t_L g1678 ( 
.A1(n_1657),
.A2(n_1637),
.B(n_1589),
.Y(n_1678)
);

AOI211x1_ASAP7_75t_SL g1679 ( 
.A1(n_1670),
.A2(n_1582),
.B(n_1606),
.C(n_1603),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1673),
.B(n_1675),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1673),
.B(n_1618),
.Y(n_1681)
);

AOI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1670),
.A2(n_1639),
.B(n_1591),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1645),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1673),
.B(n_1619),
.Y(n_1684)
);

INVxp67_ASAP7_75t_SL g1685 ( 
.A(n_1663),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1670),
.A2(n_1606),
.B1(n_1629),
.B2(n_1610),
.C(n_1609),
.Y(n_1686)
);

NAND4xp25_ASAP7_75t_L g1687 ( 
.A(n_1651),
.B(n_1579),
.C(n_1611),
.D(n_1603),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1666),
.B(n_1640),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1663),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1651),
.A2(n_1591),
.B1(n_1602),
.B2(n_1641),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1673),
.B(n_1621),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1645),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1671),
.A2(n_1586),
.B1(n_1592),
.B2(n_1601),
.C(n_1632),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1645),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1645),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1675),
.B(n_1621),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1658),
.B(n_1593),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1677),
.B(n_1593),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1648),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1646),
.A2(n_1586),
.B1(n_1592),
.B2(n_1641),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1648),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1666),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1662),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1649),
.B(n_1665),
.Y(n_1705)
);

OAI33xp33_ASAP7_75t_L g1706 ( 
.A1(n_1668),
.A2(n_1521),
.A3(n_1507),
.B1(n_1597),
.B2(n_1506),
.B3(n_1514),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1646),
.A2(n_1625),
.B1(n_1599),
.B2(n_1594),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1660),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1654),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_R g1710 ( 
.A(n_1666),
.B(n_1633),
.Y(n_1710)
);

OAI31xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1646),
.A2(n_1599),
.A3(n_1590),
.B(n_1644),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1662),
.Y(n_1712)
);

INVx4_ASAP7_75t_L g1713 ( 
.A(n_1666),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1659),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1660),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1660),
.Y(n_1716)
);

NAND4xp25_ASAP7_75t_L g1717 ( 
.A(n_1671),
.B(n_1600),
.C(n_1583),
.D(n_1640),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1714),
.B(n_1667),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1697),
.B(n_1658),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1697),
.B(n_1658),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1692),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1705),
.B(n_1646),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1705),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1683),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1685),
.B(n_1667),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1683),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1694),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1689),
.Y(n_1728)
);

AND2x2_ASAP7_75t_SL g1729 ( 
.A(n_1686),
.B(n_1647),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1692),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1694),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1695),
.Y(n_1732)
);

NAND4xp25_ASAP7_75t_L g1733 ( 
.A(n_1679),
.B(n_1647),
.C(n_1658),
.D(n_1671),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1704),
.B(n_1661),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1705),
.B(n_1647),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1709),
.B(n_1647),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1704),
.B(n_1661),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1695),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1709),
.B(n_1655),
.Y(n_1739)
);

AND2x2_ASAP7_75t_SL g1740 ( 
.A(n_1711),
.B(n_1655),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1699),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1708),
.B(n_1669),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1708),
.B(n_1661),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1715),
.B(n_1672),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1699),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1715),
.B(n_1669),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1680),
.B(n_1655),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1680),
.B(n_1655),
.Y(n_1749)
);

NAND2xp33_ASAP7_75t_R g1750 ( 
.A(n_1682),
.B(n_1631),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1701),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1701),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1696),
.B(n_1656),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1702),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1716),
.B(n_1672),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1716),
.B(n_1703),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1731),
.A2(n_1674),
.B(n_1657),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1728),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1740),
.B(n_1723),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1748),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1728),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1742),
.B(n_1698),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1724),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1724),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1729),
.B(n_1702),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1748),
.B(n_1713),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1733),
.A2(n_1690),
.B1(n_1687),
.B2(n_1700),
.C(n_1693),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1731),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1726),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1729),
.A2(n_1707),
.B1(n_1713),
.B2(n_1612),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1754),
.B(n_1713),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1726),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1727),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1754),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1740),
.B(n_1691),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1729),
.B(n_1702),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1727),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1740),
.B(n_1691),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1742),
.B(n_1703),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1723),
.B(n_1696),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1738),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1754),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1723),
.B(n_1681),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1723),
.B(n_1681),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1722),
.B(n_1678),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1738),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1746),
.B(n_1712),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1741),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1731),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1733),
.B(n_1684),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1741),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1746),
.B(n_1712),
.Y(n_1793)
);

AOI32xp33_ASAP7_75t_L g1794 ( 
.A1(n_1736),
.A2(n_1656),
.A3(n_1688),
.B1(n_1652),
.B2(n_1653),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1725),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1722),
.B(n_1678),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1718),
.B(n_1664),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1732),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1718),
.B(n_1664),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1760),
.B(n_1725),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1766),
.B(n_1595),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1782),
.B(n_1736),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1774),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1763),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1765),
.B(n_1736),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1763),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1791),
.B(n_1753),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1774),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1795),
.B(n_1753),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1767),
.B(n_1702),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1775),
.B(n_1735),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1776),
.B(n_1750),
.C(n_1702),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1795),
.B(n_1753),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1795),
.B(n_1744),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1775),
.B(n_1778),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1758),
.B(n_1719),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1764),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1771),
.B(n_1616),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1774),
.B(n_1735),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1778),
.B(n_1735),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1795),
.B(n_1744),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1757),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1759),
.B(n_1739),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1771),
.B(n_1628),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1758),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1771),
.B(n_1770),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1795),
.B(n_1755),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1764),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1757),
.Y(n_1829)
);

NAND2xp33_ASAP7_75t_L g1830 ( 
.A(n_1759),
.B(n_1509),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1788),
.B(n_1755),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1761),
.B(n_1719),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1788),
.B(n_1761),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1797),
.B(n_1739),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1769),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1780),
.B(n_1739),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1825),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1804),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1812),
.A2(n_1794),
.B1(n_1717),
.B2(n_1799),
.C(n_1796),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1810),
.A2(n_1678),
.B1(n_1796),
.B2(n_1656),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1804),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1815),
.B(n_1780),
.Y(n_1842)
);

AOI322xp5_ASAP7_75t_L g1843 ( 
.A1(n_1826),
.A2(n_1783),
.A3(n_1784),
.B1(n_1749),
.B2(n_1747),
.C1(n_1785),
.C2(n_1656),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1815),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1806),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_SL g1846 ( 
.A(n_1812),
.B(n_1784),
.C(n_1783),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1800),
.B(n_1762),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1808),
.Y(n_1848)
);

OAI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1833),
.A2(n_1785),
.B(n_1762),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1811),
.B(n_1785),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1818),
.B(n_1773),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1805),
.A2(n_1820),
.B1(n_1811),
.B2(n_1824),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1806),
.Y(n_1853)
);

OAI32xp33_ASAP7_75t_L g1854 ( 
.A1(n_1809),
.A2(n_1720),
.A3(n_1769),
.B1(n_1792),
.B2(n_1772),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1820),
.B(n_1781),
.Y(n_1855)
);

OAI322xp33_ASAP7_75t_L g1856 ( 
.A1(n_1807),
.A2(n_1772),
.A3(n_1777),
.B1(n_1792),
.B2(n_1786),
.C1(n_1789),
.C2(n_1787),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1823),
.B(n_1779),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1802),
.A2(n_1649),
.B1(n_1720),
.B2(n_1581),
.Y(n_1858)
);

XNOR2x1_ASAP7_75t_L g1859 ( 
.A(n_1823),
.B(n_1669),
.Y(n_1859)
);

NAND4xp25_ASAP7_75t_L g1860 ( 
.A(n_1801),
.B(n_1786),
.C(n_1777),
.D(n_1789),
.Y(n_1860)
);

OAI222xp33_ASAP7_75t_L g1861 ( 
.A1(n_1813),
.A2(n_1793),
.B1(n_1787),
.B2(n_1779),
.C1(n_1659),
.C2(n_1756),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1817),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1838),
.Y(n_1863)
);

AOI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1846),
.A2(n_1830),
.B1(n_1819),
.B2(n_1808),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1851),
.A2(n_1819),
.B1(n_1814),
.B2(n_1827),
.Y(n_1865)
);

NAND4xp25_ASAP7_75t_L g1866 ( 
.A(n_1852),
.B(n_1821),
.C(n_1803),
.D(n_1819),
.Y(n_1866)
);

OAI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1839),
.A2(n_1831),
.B1(n_1803),
.B2(n_1834),
.Y(n_1867)
);

O2A1O1Ixp33_ASAP7_75t_SL g1868 ( 
.A1(n_1851),
.A2(n_1803),
.B(n_1835),
.C(n_1817),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1842),
.B(n_1836),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_L g1870 ( 
.A(n_1860),
.B(n_1830),
.C(n_1835),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1841),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1844),
.A2(n_1836),
.B1(n_1828),
.B2(n_1832),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1837),
.B(n_1828),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1842),
.B(n_1816),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1853),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1862),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1848),
.Y(n_1878)
);

OAI322xp33_ASAP7_75t_L g1879 ( 
.A1(n_1855),
.A2(n_1832),
.A3(n_1816),
.B1(n_1829),
.B2(n_1822),
.C1(n_1798),
.C2(n_1790),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1857),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1847),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1852),
.B(n_1793),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1874),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1878),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1868),
.A2(n_1856),
.B(n_1854),
.Y(n_1885)
);

AOI322xp5_ASAP7_75t_L g1886 ( 
.A1(n_1867),
.A2(n_1870),
.A3(n_1881),
.B1(n_1840),
.B2(n_1882),
.C1(n_1880),
.C2(n_1872),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1865),
.A2(n_1840),
.B1(n_1849),
.B2(n_1850),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1869),
.B(n_1850),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1865),
.B(n_1859),
.Y(n_1889)
);

AOI211xp5_ASAP7_75t_L g1890 ( 
.A1(n_1879),
.A2(n_1861),
.B(n_1858),
.C(n_1822),
.Y(n_1890)
);

OA22x2_ASAP7_75t_L g1891 ( 
.A1(n_1864),
.A2(n_1829),
.B1(n_1798),
.B2(n_1790),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1866),
.B(n_1859),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1863),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1873),
.A2(n_1877),
.B(n_1876),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1888),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1886),
.B(n_1884),
.Y(n_1896)
);

NOR3x1_ASAP7_75t_L g1897 ( 
.A(n_1892),
.B(n_1875),
.C(n_1871),
.Y(n_1897)
);

NOR2x1_ASAP7_75t_L g1898 ( 
.A(n_1885),
.B(n_1768),
.Y(n_1898)
);

AOI211xp5_ASAP7_75t_L g1899 ( 
.A1(n_1889),
.A2(n_1843),
.B(n_1650),
.C(n_1768),
.Y(n_1899)
);

NAND4xp25_ASAP7_75t_L g1900 ( 
.A(n_1883),
.B(n_1649),
.C(n_1536),
.D(n_1533),
.Y(n_1900)
);

NAND3xp33_ASAP7_75t_L g1901 ( 
.A(n_1890),
.B(n_1576),
.C(n_1674),
.Y(n_1901)
);

NAND5xp2_ASAP7_75t_L g1902 ( 
.A(n_1887),
.B(n_1674),
.C(n_1747),
.D(n_1749),
.E(n_1652),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_SL g1903 ( 
.A(n_1894),
.B(n_1893),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1887),
.B(n_1747),
.Y(n_1904)
);

OAI21xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1898),
.A2(n_1891),
.B(n_1749),
.Y(n_1905)
);

XOR2x2_ASAP7_75t_L g1906 ( 
.A(n_1896),
.B(n_1649),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1895),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1901),
.A2(n_1650),
.B1(n_1706),
.B2(n_1676),
.C(n_1743),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1897),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1903),
.B(n_1756),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1909),
.B(n_1907),
.Y(n_1911)
);

AOI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1905),
.A2(n_1904),
.B1(n_1910),
.B2(n_1900),
.C(n_1899),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1906),
.B(n_1734),
.Y(n_1913)
);

A2O1A1Ixp33_ASAP7_75t_L g1914 ( 
.A1(n_1908),
.A2(n_1902),
.B(n_1581),
.C(n_1721),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1909),
.A2(n_1737),
.B1(n_1734),
.B2(n_1743),
.C(n_1745),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1910),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1916),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1911),
.Y(n_1918)
);

NAND2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1913),
.B(n_1533),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1915),
.Y(n_1920)
);

NOR2xp67_ASAP7_75t_L g1921 ( 
.A(n_1912),
.B(n_1721),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1917),
.Y(n_1922)
);

NAND3xp33_ASAP7_75t_L g1923 ( 
.A(n_1918),
.B(n_1920),
.C(n_1921),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1918),
.B(n_1914),
.Y(n_1924)
);

AO22x2_ASAP7_75t_L g1925 ( 
.A1(n_1923),
.A2(n_1919),
.B1(n_1721),
.B2(n_1730),
.Y(n_1925)
);

OAI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1925),
.A2(n_1922),
.B1(n_1924),
.B2(n_1756),
.Y(n_1926)
);

NOR3xp33_ASAP7_75t_L g1927 ( 
.A(n_1926),
.B(n_1513),
.C(n_1568),
.Y(n_1927)
);

AO22x2_ASAP7_75t_L g1928 ( 
.A1(n_1926),
.A2(n_1730),
.B1(n_1752),
.B2(n_1732),
.Y(n_1928)
);

OAI22x1_ASAP7_75t_SL g1929 ( 
.A1(n_1927),
.A2(n_1492),
.B1(n_1547),
.B2(n_1559),
.Y(n_1929)
);

AOI222xp33_ASAP7_75t_L g1930 ( 
.A1(n_1928),
.A2(n_1751),
.B1(n_1745),
.B2(n_1730),
.C1(n_1732),
.C2(n_1752),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1930),
.B(n_1737),
.Y(n_1931)
);

AOI221xp5_ASAP7_75t_SL g1932 ( 
.A1(n_1929),
.A2(n_1751),
.B1(n_1752),
.B2(n_1509),
.C(n_1654),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1931),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1933),
.B(n_1932),
.Y(n_1934)
);

OAI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1934),
.A2(n_1509),
.B1(n_1492),
.B2(n_1559),
.Y(n_1935)
);

OAI221xp5_ASAP7_75t_R g1936 ( 
.A1(n_1935),
.A2(n_1654),
.B1(n_1575),
.B2(n_1547),
.C(n_1536),
.Y(n_1936)
);

AOI211xp5_ASAP7_75t_L g1937 ( 
.A1(n_1936),
.A2(n_1536),
.B(n_1533),
.C(n_1570),
.Y(n_1937)
);


endmodule