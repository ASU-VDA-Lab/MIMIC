module fake_jpeg_31470_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_61),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_0),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_74),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_48),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_46),
.B1(n_53),
.B2(n_45),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_87),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_52),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_0),
.C(n_1),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_89),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_53),
.B1(n_70),
.B2(n_44),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_69),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_49),
.B(n_42),
.Y(n_90)
);

OAI211xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_22),
.B(n_36),
.C(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_39),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_17),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_9),
.C(n_10),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_107),
.C(n_8),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_88),
.Y(n_101)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_87),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_108),
.C(n_16),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_1),
.B(n_2),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_7),
.B(n_8),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_21),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_112),
.B1(n_115),
.B2(n_100),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_118),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_120),
.B(n_100),
.C(n_95),
.D(n_103),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_124),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_94),
.C(n_120),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_116),
.C(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_127),
.C(n_128),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_12),
.B(n_14),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_20),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_24),
.C(n_25),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_110),
.B(n_28),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_26),
.Y(n_135)
);


endmodule