module fake_netlist_5_2472_n_1833 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1833);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1833;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1584;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1715;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_87),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_17),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_55),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_30),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_47),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_48),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_55),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_43),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_61),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_102),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_3),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_70),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_54),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_122),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_15),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_110),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_48),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_86),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_90),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_76),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_42),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_113),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_92),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_47),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_14),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_20),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_82),
.Y(n_211)
);

BUFx8_ASAP7_75t_SL g212 ( 
.A(n_46),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_10),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_35),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_41),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_22),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_85),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_1),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_150),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_104),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_144),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_40),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_133),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_31),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_152),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_101),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_35),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_142),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_37),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_167),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_79),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_57),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_8),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_114),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_103),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_154),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_19),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_8),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_43),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_119),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_89),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_28),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_137),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_161),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

INVxp33_ASAP7_75t_SL g257 ( 
.A(n_9),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_42),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_52),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_166),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_30),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_162),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_120),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_72),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_6),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_28),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_68),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_77),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_49),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_15),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_124),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_117),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_168),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_127),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_74),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_75),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_27),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_54),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_1),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_123),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_97),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_7),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_121),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_44),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_2),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_58),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_95),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_52),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_147),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_155),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_80),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_81),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_83),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_160),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_23),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_99),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_46),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_138),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_64),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_29),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_107),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_53),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_146),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_9),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_4),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_32),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_67),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_58),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_153),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_134),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_111),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_65),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_112),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_51),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_164),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_56),
.Y(n_317)
);

BUFx8_ASAP7_75t_SL g318 ( 
.A(n_93),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_94),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_125),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_3),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_36),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_39),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_140),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_36),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_24),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_21),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_96),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_22),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_13),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_130),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_33),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_91),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_19),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_45),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_78),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_71),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_63),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_57),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_34),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_222),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_222),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_224),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_210),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_302),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_318),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_212),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_171),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_222),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_222),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_222),
.Y(n_351)
);

BUFx6f_ASAP7_75t_SL g352 ( 
.A(n_190),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_222),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_226),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_296),
.B(n_339),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_174),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_222),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_222),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_222),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_247),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_175),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_263),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_210),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_184),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_273),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_185),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_173),
.B(n_181),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_247),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_210),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_316),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_186),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_176),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_177),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_325),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_173),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_210),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_302),
.B(n_0),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_182),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_210),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_210),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_198),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_337),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_325),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_198),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_203),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_203),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_215),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_281),
.B(n_4),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_303),
.B(n_5),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_215),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_182),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_214),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_206),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_218),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_214),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_176),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_237),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_189),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_193),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_237),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_280),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_280),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_292),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_305),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_194),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_181),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_196),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_303),
.B(n_5),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_305),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_197),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_305),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_200),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_202),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_187),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_187),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_204),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_178),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_201),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_394),
.B(n_238),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_281),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_372),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_379),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_378),
.A2(n_172),
.B1(n_285),
.B2(n_334),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_388),
.A2(n_249),
.B1(n_209),
.B2(n_257),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_206),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_377),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_380),
.A2(n_220),
.B(n_201),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_369),
.B(n_308),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_308),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_342),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_390),
.B(n_292),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_350),
.B(n_308),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_350),
.B(n_218),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_351),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_372),
.B(n_331),
.Y(n_457)
);

BUFx8_ASAP7_75t_L g458 ( 
.A(n_352),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_391),
.A2(n_404),
.B1(n_368),
.B2(n_375),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_413),
.B(n_190),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_419),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_353),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_353),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_360),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_357),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_321),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_357),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_321),
.Y(n_470)
);

OA21x2_ASAP7_75t_L g471 ( 
.A1(n_358),
.A2(n_235),
.B(n_220),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_420),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_358),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_359),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_359),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_372),
.B(n_331),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_392),
.B(n_183),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_408),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_395),
.B(n_205),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_387),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_387),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_384),
.B(n_195),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_373),
.A2(n_241),
.B(n_235),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_393),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_389),
.B(n_207),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_408),
.B(n_183),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_422),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_367),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_367),
.B(n_315),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_374),
.B(n_190),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_497),
.B(n_348),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_447),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_471),
.Y(n_502)
);

OR2x6_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_435),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_483),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_356),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_471),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_361),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_364),
.Y(n_509)
);

NOR3xp33_ASAP7_75t_L g510 ( 
.A(n_436),
.B(n_499),
.C(n_453),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_435),
.Y(n_511)
);

AND3x1_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_322),
.C(n_315),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_425),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_453),
.B(n_366),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_471),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_434),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_424),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_428),
.B(n_371),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_437),
.B(n_399),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_447),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_345),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_465),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_477),
.B(n_396),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_439),
.B(n_436),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_477),
.B(n_396),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_471),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_471),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_437),
.B(n_400),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_465),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_398),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_499),
.B(n_409),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_428),
.B(n_411),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_425),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_495),
.A2(n_322),
.B1(n_343),
.B2(n_298),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_485),
.B(n_415),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_445),
.B(n_297),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_433),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_498),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_440),
.B(n_398),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_489),
.B(n_417),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_495),
.A2(n_317),
.B1(n_267),
.B2(n_340),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_454),
.B(n_297),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_496),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_495),
.B(n_191),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_485),
.B(n_418),
.Y(n_549)
);

AND3x2_ASAP7_75t_L g550 ( 
.A(n_496),
.B(n_312),
.C(n_216),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_433),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_458),
.B(n_421),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_433),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_454),
.A2(n_241),
.B1(n_267),
.B2(n_298),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_440),
.B(n_401),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_498),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_456),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_440),
.B(n_401),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_498),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_447),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_449),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_447),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_493),
.B(n_236),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_459),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_463),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_424),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_447),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_459),
.B(n_191),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_463),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_493),
.B(n_252),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_455),
.B(n_211),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_424),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_463),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_455),
.B(n_213),
.Y(n_579)
);

CKINVDCx6p67_ASAP7_75t_R g580 ( 
.A(n_461),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_438),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_434),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_455),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_447),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_447),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_467),
.Y(n_586)
);

BUFx8_ASAP7_75t_SL g587 ( 
.A(n_468),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_438),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_438),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_454),
.A2(n_317),
.B1(n_335),
.B2(n_340),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_455),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_454),
.A2(n_335),
.B1(n_312),
.B2(n_352),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_458),
.B(n_346),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_468),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_441),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_424),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_441),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_458),
.B(n_347),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_467),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_455),
.A2(n_265),
.B(n_221),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_441),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_458),
.B(n_190),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_467),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_461),
.B(n_352),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_458),
.B(n_199),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_447),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_441),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_455),
.B(n_217),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

INVx4_ASAP7_75t_SL g610 ( 
.A(n_474),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_474),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_467),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_449),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_474),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_467),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_474),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_494),
.B(n_354),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_460),
.Y(n_618)
);

AND3x2_ASAP7_75t_L g619 ( 
.A(n_449),
.B(n_221),
.C(n_216),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_460),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_460),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_454),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

OR2x6_ASAP7_75t_L g625 ( 
.A(n_431),
.B(n_223),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_494),
.B(n_362),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_468),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_454),
.B(n_225),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_470),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_470),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_464),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_458),
.B(n_199),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_469),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_474),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_469),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_469),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_431),
.A2(n_248),
.B1(n_262),
.B2(n_261),
.Y(n_638)
);

CKINVDCx6p67_ASAP7_75t_R g639 ( 
.A(n_494),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_439),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_457),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_469),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_448),
.B(n_227),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_448),
.B(n_199),
.Y(n_644)
);

OAI21xp33_ASAP7_75t_L g645 ( 
.A1(n_462),
.A2(n_410),
.B(n_376),
.Y(n_645)
);

BUFx8_ASAP7_75t_SL g646 ( 
.A(n_448),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_448),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_490),
.A2(n_272),
.B1(n_223),
.B2(n_242),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_473),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_473),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_547),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_533),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_519),
.B(n_365),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_641),
.B(n_474),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_622),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_622),
.B(n_474),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_511),
.B(n_474),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_583),
.B(n_473),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_583),
.B(n_591),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_591),
.B(n_473),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_502),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_533),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_535),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_566),
.B(n_475),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_547),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_535),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_557),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_504),
.B(n_323),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_566),
.B(n_475),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_543),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_511),
.B(n_445),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_531),
.B(n_370),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_543),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_516),
.B(n_445),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_557),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_502),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_600),
.B(n_291),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_559),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_613),
.B(n_475),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_613),
.B(n_475),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_530),
.B(n_568),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_556),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_559),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_575),
.B(n_445),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_547),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_506),
.B(n_242),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_540),
.B(n_291),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_582),
.B(n_445),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_540),
.B(n_291),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_561),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_547),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_540),
.B(n_291),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_506),
.A2(n_476),
.B(n_457),
.C(n_462),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_563),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_556),
.Y(n_696)
);

OAI21xp33_ASAP7_75t_L g697 ( 
.A1(n_542),
.A2(n_423),
.B(n_466),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_582),
.B(n_445),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_563),
.Y(n_699)
);

INVx8_ASAP7_75t_L g700 ( 
.A(n_503),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_531),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_505),
.B(n_490),
.Y(n_702)
);

NOR2xp67_ASAP7_75t_SL g703 ( 
.A(n_507),
.B(n_243),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_539),
.B(n_490),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_549),
.B(n_490),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_518),
.B(n_383),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_570),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_628),
.B(n_490),
.Y(n_708)
);

INVx8_ASAP7_75t_L g709 ( 
.A(n_503),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_504),
.B(n_490),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_594),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_562),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_510),
.B(n_291),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_544),
.B(n_180),
.C(n_179),
.Y(n_714)
);

BUFx6f_ASAP7_75t_SL g715 ( 
.A(n_573),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_628),
.B(n_476),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_648),
.A2(n_448),
.B1(n_243),
.B2(n_250),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_503),
.A2(n_284),
.B1(n_250),
.B2(n_251),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_594),
.Y(n_719)
);

OAI221xp5_ASAP7_75t_L g720 ( 
.A1(n_545),
.A2(n_472),
.B1(n_482),
.B2(n_260),
.C(n_251),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_570),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_517),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_522),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_562),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_500),
.B(n_291),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_523),
.B(n_472),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_508),
.B(n_291),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_536),
.B(n_188),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_507),
.B(n_443),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_515),
.B(n_443),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_509),
.B(n_515),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_528),
.B(n_291),
.Y(n_732)
);

AND2x6_ASAP7_75t_L g733 ( 
.A(n_528),
.B(n_260),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_529),
.B(n_427),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_574),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_542),
.A2(n_482),
.B(n_426),
.C(n_429),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_574),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_517),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_647),
.B(n_291),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_578),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_521),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_503),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_558),
.B(n_192),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_630),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_578),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_631),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_521),
.B(n_423),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_503),
.B(n_432),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_513),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_548),
.B(n_264),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_517),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_513),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_523),
.B(n_432),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_527),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_527),
.B(n_532),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_532),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_586),
.B(n_442),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_524),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_517),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_558),
.A2(n_426),
.B(n_429),
.C(n_430),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_647),
.B(n_230),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_587),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_524),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_564),
.B(n_208),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_564),
.B(n_232),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_548),
.A2(n_277),
.B1(n_268),
.B2(n_264),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_580),
.B(n_514),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_629),
.B(n_233),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_586),
.B(n_442),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_576),
.B(n_234),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_580),
.B(n_219),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_525),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_579),
.A2(n_429),
.B(n_426),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_534),
.B(n_228),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_599),
.B(n_430),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_617),
.A2(n_300),
.B1(n_239),
.B2(n_245),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_599),
.B(n_430),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_525),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_517),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_608),
.B(n_254),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_619),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_626),
.B(n_229),
.Y(n_783)
);

INVxp33_ASAP7_75t_SL g784 ( 
.A(n_526),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_538),
.B(n_487),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_SL g786 ( 
.A(n_640),
.B(n_271),
.C(n_270),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_603),
.B(n_255),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_552),
.B(n_268),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_548),
.B(n_487),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_603),
.B(n_444),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_548),
.B(n_231),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_537),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_612),
.B(n_444),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_612),
.B(n_269),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_537),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_615),
.B(n_444),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_550),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_615),
.B(n_274),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_541),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_541),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_548),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_638),
.B(n_240),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_512),
.B(n_487),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_512),
.B(n_488),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_618),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_604),
.B(n_644),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_526),
.B(n_266),
.C(n_258),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_SL g808 ( 
.A(n_640),
.B(n_199),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_643),
.B(n_446),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_551),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_639),
.B(n_446),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_645),
.B(n_488),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_639),
.B(n_645),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_625),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_646),
.B(n_244),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_R g816 ( 
.A(n_569),
.B(n_275),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_551),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_553),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_501),
.B(n_450),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_654),
.A2(n_611),
.B(n_572),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_688),
.A2(n_693),
.B(n_690),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_674),
.A2(n_611),
.B(n_572),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_774),
.A2(n_520),
.B(n_501),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_657),
.A2(n_611),
.B(n_572),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_681),
.A2(n_806),
.B1(n_661),
.B2(n_813),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_711),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_716),
.B(n_625),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_711),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_652),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_807),
.B(n_598),
.C(n_593),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_756),
.B(n_592),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_702),
.A2(n_625),
.B1(n_605),
.B2(n_602),
.Y(n_832)
);

O2A1O1Ixp5_ASAP7_75t_L g833 ( 
.A1(n_703),
.A2(n_633),
.B(n_584),
.C(n_567),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_671),
.A2(n_572),
.B(n_606),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_668),
.B(n_573),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_704),
.A2(n_616),
.B(n_606),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_741),
.B(n_625),
.Y(n_837)
);

AND2x6_ASAP7_75t_L g838 ( 
.A(n_676),
.B(n_520),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_705),
.A2(n_616),
.B(n_606),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_656),
.A2(n_616),
.B(n_606),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_652),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_656),
.A2(n_616),
.B(n_606),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_728),
.B(n_625),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_700),
.B(n_546),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_662),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_726),
.B(n_555),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_755),
.A2(n_757),
.B(n_677),
.C(n_783),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_726),
.B(n_590),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_738),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_662),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_719),
.B(n_573),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_SL g852 ( 
.A(n_808),
.B(n_816),
.C(n_653),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_726),
.B(n_546),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_663),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_663),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_658),
.A2(n_577),
.B(n_571),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_658),
.A2(n_577),
.B(n_571),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_747),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_660),
.A2(n_577),
.B(n_571),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_676),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_666),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_670),
.B(n_573),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_660),
.A2(n_577),
.B(n_571),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_719),
.B(n_573),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_710),
.B(n_520),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_809),
.A2(n_596),
.B(n_571),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_744),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_713),
.A2(n_677),
.B(n_731),
.C(n_708),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_754),
.B(n_546),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_812),
.B(n_546),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_746),
.B(n_402),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_689),
.A2(n_596),
.B(n_584),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_698),
.A2(n_596),
.B(n_584),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_701),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_706),
.B(n_567),
.Y(n_875)
);

NOR2x1_ASAP7_75t_L g876 ( 
.A(n_768),
.B(n_567),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_743),
.B(n_765),
.C(n_775),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_676),
.B(n_546),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_713),
.A2(n_546),
.B1(n_272),
.B2(n_277),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_738),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_731),
.A2(n_621),
.B(n_649),
.C(n_642),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_667),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_738),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_803),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_690),
.A2(n_623),
.B(n_649),
.C(n_642),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_673),
.B(n_596),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_801),
.A2(n_284),
.B1(n_336),
.B2(n_304),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_772),
.B(n_290),
.C(n_295),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_797),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_734),
.A2(n_614),
.B(n_585),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_682),
.B(n_585),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_675),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_696),
.B(n_614),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_729),
.A2(n_730),
.B(n_659),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_659),
.A2(n_614),
.B(n_635),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_752),
.B(n_635),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_712),
.B(n_635),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_675),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_722),
.A2(n_565),
.B(n_588),
.Y(n_899)
);

INVx5_ASAP7_75t_L g900 ( 
.A(n_700),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_724),
.A2(n_336),
.B(n_295),
.C(n_299),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_804),
.B(n_623),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_693),
.A2(n_637),
.B(n_636),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_678),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_789),
.B(n_624),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_683),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_683),
.B(n_624),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_685),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_685),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_651),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_691),
.Y(n_911)
);

AOI21x1_ASAP7_75t_L g912 ( 
.A1(n_664),
.A2(n_627),
.B(n_637),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_738),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_722),
.A2(n_565),
.B(n_560),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_684),
.A2(n_636),
.B(n_634),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_718),
.A2(n_290),
.B(n_299),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_687),
.A2(n_733),
.B1(n_695),
.B2(n_699),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_691),
.B(n_627),
.Y(n_918)
);

AND2x6_ASAP7_75t_SL g919 ( 
.A(n_815),
.B(n_304),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_695),
.B(n_632),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_782),
.B(n_488),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_699),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_785),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_802),
.B(n_632),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_707),
.B(n_634),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_707),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_655),
.A2(n_650),
.B1(n_620),
.B2(n_609),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_732),
.A2(n_650),
.B(n_620),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_721),
.B(n_610),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_721),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_735),
.B(n_560),
.Y(n_931)
);

NOR2x1p5_ASAP7_75t_L g932 ( 
.A(n_701),
.B(n_246),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_791),
.B(n_723),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_735),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_737),
.B(n_581),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_737),
.B(n_581),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_740),
.B(n_745),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_722),
.A2(n_565),
.B(n_609),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_740),
.B(n_588),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_748),
.A2(n_565),
.B(n_607),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_732),
.A2(n_595),
.B(n_607),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_664),
.A2(n_565),
.B(n_601),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_745),
.B(n_589),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_665),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_811),
.B(n_610),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_694),
.A2(n_601),
.B(n_597),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_814),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_739),
.A2(n_597),
.B(n_595),
.C(n_589),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_749),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_787),
.A2(n_333),
.B1(n_282),
.B2(n_288),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_686),
.B(n_402),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_805),
.Y(n_952)
);

CKINVDCx10_ASAP7_75t_R g953 ( 
.A(n_715),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_669),
.A2(n_554),
.B(n_553),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_669),
.A2(n_565),
.B(n_554),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_679),
.A2(n_610),
.B(n_450),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_760),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_679),
.A2(n_610),
.B(n_450),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_680),
.A2(n_451),
.B(n_491),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_749),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_680),
.A2(n_451),
.B(n_491),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_753),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_725),
.A2(n_451),
.B(n_491),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_753),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_725),
.A2(n_492),
.B(n_491),
.Y(n_965)
);

NAND2x1p5_ASAP7_75t_L g966 ( 
.A(n_760),
.B(n_478),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_692),
.B(n_403),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_717),
.B(n_276),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_727),
.A2(n_492),
.B(n_486),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_727),
.A2(n_492),
.B(n_486),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_723),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_700),
.A2(n_319),
.B1(n_293),
.B2(n_294),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_766),
.B(n_253),
.Y(n_973)
);

INVx8_ASAP7_75t_L g974 ( 
.A(n_700),
.Y(n_974)
);

CKINVDCx6p67_ASAP7_75t_R g975 ( 
.A(n_715),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_759),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_697),
.B(n_310),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_687),
.B(n_311),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_763),
.B(n_777),
.Y(n_979)
);

O2A1O1Ixp5_ASAP7_75t_L g980 ( 
.A1(n_739),
.A2(n_492),
.B(n_486),
.C(n_480),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_720),
.A2(n_256),
.B(n_259),
.C(n_278),
.Y(n_981)
);

AO21x2_ASAP7_75t_L g982 ( 
.A1(n_787),
.A2(n_794),
.B(n_798),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_709),
.A2(n_328),
.B1(n_313),
.B2(n_314),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_766),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_672),
.B(n_403),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_736),
.A2(n_329),
.B(n_283),
.C(n_286),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_687),
.B(n_320),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_714),
.B(n_405),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_759),
.Y(n_989)
);

AOI211xp5_ASAP7_75t_L g990 ( 
.A1(n_767),
.A2(n_279),
.B(n_287),
.C(n_289),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_687),
.B(n_324),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_751),
.A2(n_486),
.B(n_480),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_687),
.A2(n_733),
.B(n_819),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_794),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_760),
.B(n_709),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_687),
.A2(n_480),
.B(n_338),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_761),
.A2(n_301),
.B(n_306),
.C(n_307),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_751),
.A2(n_480),
.B(n_481),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_709),
.A2(n_309),
.B1(n_327),
.B2(n_332),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_750),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_760),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_733),
.B(n_484),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_750),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_764),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_825),
.B(n_788),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_877),
.A2(n_742),
.B1(n_709),
.B2(n_750),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_923),
.B(n_788),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_849),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_923),
.B(n_733),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_894),
.A2(n_742),
.B(n_780),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_868),
.A2(n_742),
.B(n_780),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_971),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_874),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_SL g1014 ( 
.A(n_971),
.B(n_784),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_855),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_984),
.A2(n_742),
.B(n_798),
.C(n_762),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_870),
.A2(n_769),
.B(n_781),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_984),
.B(n_784),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_821),
.A2(n_733),
.B(n_770),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_844),
.A2(n_769),
.B(n_781),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_924),
.A2(n_750),
.B1(n_762),
.B2(n_771),
.Y(n_1021)
);

O2A1O1Ixp5_ASAP7_75t_L g1022 ( 
.A1(n_843),
.A2(n_771),
.B(n_776),
.C(n_778),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_858),
.B(n_758),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_855),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_SL g1025 ( 
.A1(n_917),
.A2(n_793),
.B(n_790),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_884),
.B(n_786),
.Y(n_1026)
);

OAI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_884),
.A2(n_796),
.B1(n_715),
.B2(n_810),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_924),
.B(n_733),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_994),
.B(n_764),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_888),
.A2(n_818),
.B(n_817),
.C(n_810),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_875),
.B(n_773),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_862),
.B(n_773),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_985),
.B(n_405),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_869),
.A2(n_818),
.B(n_817),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_822),
.A2(n_800),
.B(n_799),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_841),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_847),
.A2(n_800),
.B(n_799),
.C(n_795),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_862),
.B(n_837),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_852),
.B(n_116),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_888),
.A2(n_795),
.B(n_792),
.C(n_779),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_SL g1041 ( 
.A1(n_851),
.A2(n_412),
.B1(n_407),
.B2(n_406),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_SL g1042 ( 
.A1(n_847),
.A2(n_792),
.B(n_779),
.C(n_412),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_SL g1043 ( 
.A(n_851),
.B(n_407),
.C(n_406),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_830),
.B(n_484),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_953),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_875),
.A2(n_484),
.B(n_481),
.C(n_479),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_835),
.B(n_6),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_827),
.A2(n_484),
.B(n_481),
.C(n_479),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_902),
.B(n_952),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_849),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_830),
.B(n_484),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_867),
.B(n_10),
.Y(n_1052)
);

CKINVDCx14_ASAP7_75t_R g1053 ( 
.A(n_933),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_860),
.B(n_484),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_974),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_826),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_979),
.A2(n_831),
.B1(n_832),
.B2(n_864),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_909),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_860),
.B(n_905),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_849),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_826),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_828),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_981),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_932),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_846),
.B(n_484),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_981),
.A2(n_11),
.B(n_12),
.C(n_16),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_909),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_831),
.A2(n_481),
.B(n_479),
.C(n_478),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_848),
.B(n_481),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_867),
.B(n_16),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_865),
.A2(n_481),
.B(n_479),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_820),
.A2(n_481),
.B(n_479),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_828),
.B(n_479),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_974),
.B(n_158),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_951),
.B(n_479),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_967),
.B(n_479),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_898),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_878),
.A2(n_478),
.B(n_148),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_871),
.B(n_478),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_986),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_834),
.A2(n_478),
.B(n_141),
.Y(n_1081)
);

AND2x6_ASAP7_75t_L g1082 ( 
.A(n_853),
.B(n_898),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_865),
.B(n_478),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_973),
.B(n_478),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_849),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_896),
.B(n_478),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_947),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_993),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1088)
);

AO21x1_ASAP7_75t_L g1089 ( 
.A1(n_945),
.A2(n_25),
.B(n_26),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_921),
.B(n_29),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_945),
.A2(n_139),
.B(n_132),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_921),
.B(n_31),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_986),
.A2(n_997),
.B(n_917),
.C(n_833),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_975),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_836),
.A2(n_126),
.B(n_118),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_839),
.A2(n_866),
.B(n_824),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_896),
.B(n_32),
.Y(n_1097)
);

AND2x2_ASAP7_75t_SL g1098 ( 
.A(n_879),
.B(n_105),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_889),
.B(n_1000),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_919),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_879),
.A2(n_100),
.B1(n_98),
.B2(n_88),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_906),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_906),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_910),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_872),
.A2(n_84),
.B(n_73),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_988),
.A2(n_33),
.B(n_34),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_873),
.A2(n_69),
.B(n_66),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_900),
.A2(n_62),
.B1(n_38),
.B2(n_39),
.Y(n_1108)
);

BUFx12f_ASAP7_75t_L g1109 ( 
.A(n_1003),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_990),
.B(n_950),
.C(n_916),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_910),
.B(n_37),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_886),
.B(n_911),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_937),
.A2(n_38),
.B(n_40),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_944),
.B(n_41),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_900),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_900),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_915),
.A2(n_59),
.B(n_60),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_944),
.B(n_59),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_911),
.A2(n_922),
.B1(n_892),
.B2(n_904),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_997),
.A2(n_887),
.B(n_901),
.C(n_977),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_982),
.A2(n_886),
.B1(n_968),
.B2(n_972),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_974),
.B(n_900),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_999),
.B(n_891),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_903),
.A2(n_859),
.B(n_857),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_922),
.B(n_845),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1004),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_856),
.A2(n_863),
.B(n_890),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_880),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_829),
.B(n_861),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_907),
.A2(n_925),
.B(n_918),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_901),
.A2(n_897),
.B(n_893),
.C(n_983),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_850),
.B(n_854),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_908),
.A2(n_934),
.B1(n_930),
.B2(n_926),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1004),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_882),
.B(n_949),
.Y(n_1135)
);

OAI22x1_ASAP7_75t_L g1136 ( 
.A1(n_995),
.A2(n_876),
.B1(n_929),
.B2(n_989),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_962),
.B(n_964),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_982),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_960),
.B(n_976),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_920),
.B(n_943),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_880),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_931),
.B(n_935),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_957),
.B(n_1001),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_913),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_913),
.B(n_883),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_957),
.B(n_1001),
.Y(n_1146)
);

NOR2xp67_ASAP7_75t_L g1147 ( 
.A(n_978),
.B(n_987),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_913),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_883),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_936),
.B(n_939),
.Y(n_1150)
);

CKINVDCx11_ASAP7_75t_R g1151 ( 
.A(n_1012),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1036),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1018),
.B(n_991),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1010),
.A2(n_823),
.B(n_912),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1057),
.A2(n_1120),
.B(n_1021),
.C(n_1098),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1048),
.A2(n_940),
.A3(n_1002),
.B(n_970),
.Y(n_1156)
);

BUFx4_ASAP7_75t_SL g1157 ( 
.A(n_1094),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1033),
.B(n_995),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1035),
.A2(n_946),
.B(n_895),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1093),
.A2(n_980),
.B(n_965),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1056),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1020),
.A2(n_996),
.B(n_938),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1130),
.A2(n_899),
.B(n_914),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_1098),
.B(n_838),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1072),
.A2(n_941),
.B(n_928),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1014),
.B(n_927),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1104),
.B(n_840),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1117),
.A2(n_969),
.B1(n_963),
.B2(n_842),
.C(n_998),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_SL g1169 ( 
.A(n_1122),
.B(n_838),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1038),
.B(n_1023),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_1047),
.A2(n_1097),
.B1(n_1026),
.B2(n_1118),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1106),
.B(n_885),
.C(n_959),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1016),
.A2(n_948),
.B(n_881),
.C(n_958),
.Y(n_1173)
);

O2A1O1Ixp5_ASAP7_75t_L g1174 ( 
.A1(n_1097),
.A2(n_929),
.B(n_954),
.C(n_956),
.Y(n_1174)
);

INVx6_ASAP7_75t_L g1175 ( 
.A(n_1109),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1096),
.A2(n_1034),
.B(n_1127),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1013),
.B(n_942),
.Y(n_1177)
);

OA21x2_ASAP7_75t_L g1178 ( 
.A1(n_1046),
.A2(n_992),
.B(n_961),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1068),
.A2(n_955),
.A3(n_838),
.B(n_966),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1138),
.A2(n_1136),
.A3(n_1124),
.B(n_1011),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1022),
.A2(n_838),
.B(n_966),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1055),
.Y(n_1182)
);

INVx8_ASAP7_75t_L g1183 ( 
.A(n_1008),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1019),
.A2(n_1017),
.B(n_1140),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1087),
.Y(n_1185)
);

AO21x1_ASAP7_75t_L g1186 ( 
.A1(n_1005),
.A2(n_1028),
.B(n_1051),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1008),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1142),
.A2(n_1150),
.B(n_1031),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1049),
.B(n_1059),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1129),
.B(n_1137),
.Y(n_1190)
);

CKINVDCx11_ASAP7_75t_R g1191 ( 
.A(n_1064),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1037),
.A2(n_1089),
.A3(n_1088),
.B(n_1083),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1081),
.A2(n_1065),
.B(n_1069),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1008),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1133),
.A2(n_1086),
.A3(n_1006),
.B(n_1078),
.Y(n_1195)
);

OAI22x1_ASAP7_75t_L g1196 ( 
.A1(n_1047),
.A2(n_1118),
.B1(n_1111),
.B2(n_1114),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1061),
.Y(n_1197)
);

BUFx4f_ASAP7_75t_L g1198 ( 
.A(n_1008),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1063),
.A2(n_1066),
.B(n_1080),
.C(n_1027),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1027),
.A2(n_1110),
.B(n_1007),
.C(n_1115),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1147),
.A2(n_1071),
.B(n_1022),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1009),
.A2(n_1054),
.A3(n_1137),
.B(n_1105),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1025),
.A2(n_1131),
.B(n_1121),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1044),
.A2(n_1084),
.B(n_1132),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1075),
.A2(n_1076),
.B(n_1042),
.Y(n_1205)
);

O2A1O1Ixp5_ASAP7_75t_L g1206 ( 
.A1(n_1107),
.A2(n_1095),
.B(n_1091),
.C(n_1145),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1110),
.A2(n_1123),
.B(n_1043),
.C(n_1030),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1079),
.A2(n_1112),
.B(n_1040),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1090),
.A2(n_1070),
.B(n_1052),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1099),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1043),
.A2(n_1090),
.B(n_1032),
.C(n_1101),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1100),
.A2(n_1061),
.B1(n_1062),
.B2(n_1052),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1119),
.A2(n_1125),
.B1(n_1077),
.B2(n_1102),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1062),
.B(n_1073),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1082),
.A2(n_1119),
.B(n_1135),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1050),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1139),
.A2(n_1029),
.B(n_1103),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1143),
.A2(n_1146),
.B(n_1149),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1143),
.A2(n_1146),
.B(n_1149),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1045),
.Y(n_1220)
);

NOR4xp25_ASAP7_75t_L g1221 ( 
.A(n_1116),
.B(n_1108),
.C(n_1070),
.D(n_1092),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1113),
.A2(n_1134),
.B(n_1126),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1015),
.B(n_1024),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1058),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1053),
.B(n_1067),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1128),
.Y(n_1226)
);

NOR2xp67_ASAP7_75t_L g1227 ( 
.A(n_1144),
.B(n_1141),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1041),
.A2(n_1050),
.B1(n_1060),
.B2(n_1085),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1050),
.Y(n_1229)
);

AOI21x1_ASAP7_75t_SL g1230 ( 
.A1(n_1039),
.A2(n_1082),
.B(n_1060),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1060),
.B(n_1085),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1060),
.A2(n_1085),
.B(n_1082),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1082),
.B(n_1038),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1082),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1057),
.A2(n_681),
.B(n_877),
.C(n_510),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1237)
);

OAI22x1_ASAP7_75t_L g1238 ( 
.A1(n_1057),
.A2(n_526),
.B1(n_877),
.B2(n_851),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1033),
.B(n_711),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1026),
.A2(n_681),
.B(n_499),
.C(n_510),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1241)
);

NAND2xp33_ASAP7_75t_SL g1242 ( 
.A(n_1074),
.B(n_1012),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1036),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1020),
.A2(n_1130),
.B(n_844),
.Y(n_1245)
);

BUFx2_ASAP7_75t_SL g1246 ( 
.A(n_1012),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1018),
.B(n_521),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1098),
.A2(n_510),
.B1(n_681),
.B2(n_877),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1048),
.A2(n_1046),
.A3(n_1068),
.B(n_1093),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1013),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1018),
.B(n_681),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1055),
.B(n_900),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1253)
);

O2A1O1Ixp5_ASAP7_75t_L g1254 ( 
.A1(n_1117),
.A2(n_877),
.B(n_681),
.C(n_783),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1016),
.A2(n_1088),
.B(n_1093),
.C(n_843),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1038),
.B(n_1055),
.Y(n_1256)
);

AO32x2_ASAP7_75t_L g1257 ( 
.A1(n_1021),
.A2(n_825),
.A3(n_832),
.B1(n_1006),
.B2(n_1133),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1020),
.A2(n_1130),
.B(n_844),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1013),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_L g1260 ( 
.A(n_1013),
.B(n_984),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1049),
.B(n_681),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1013),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1048),
.A2(n_1046),
.A3(n_1068),
.B(n_1093),
.Y(n_1263)
);

AO21x2_ASAP7_75t_L g1264 ( 
.A1(n_1016),
.A2(n_1096),
.B(n_1011),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1018),
.B(n_681),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1033),
.B(n_711),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1055),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1093),
.A2(n_847),
.B(n_1022),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1055),
.B(n_900),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1093),
.A2(n_847),
.B(n_1022),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1020),
.A2(n_1130),
.B(n_844),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1020),
.A2(n_1130),
.B(n_844),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1012),
.Y(n_1276)
);

AO21x1_ASAP7_75t_L g1277 ( 
.A1(n_1021),
.A2(n_1117),
.B(n_1005),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1093),
.A2(n_847),
.B(n_1022),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1012),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1104),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1020),
.A2(n_1130),
.B(n_844),
.Y(n_1281)
);

AOI221x1_ASAP7_75t_L g1282 ( 
.A1(n_1117),
.A2(n_888),
.B1(n_1088),
.B2(n_877),
.C(n_510),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1048),
.A2(n_1046),
.A3(n_1068),
.B(n_1093),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1038),
.B(n_1055),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1014),
.B(n_672),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1049),
.B(n_681),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1010),
.A2(n_1035),
.B(n_1072),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1048),
.A2(n_1046),
.A3(n_1068),
.B(n_1093),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1020),
.A2(n_1130),
.B(n_844),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1093),
.A2(n_847),
.B(n_1022),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1046),
.A2(n_1068),
.B(n_1048),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1020),
.A2(n_1130),
.B(n_844),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1038),
.B(n_1055),
.Y(n_1294)
);

CKINVDCx11_ASAP7_75t_R g1295 ( 
.A(n_1012),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1055),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1049),
.B(n_681),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_SL g1298 ( 
.A1(n_1016),
.A2(n_1088),
.B(n_1093),
.C(n_843),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1098),
.A2(n_681),
.B1(n_825),
.B2(n_877),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1093),
.A2(n_847),
.B(n_1022),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1018),
.B(n_521),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1152),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1185),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1164),
.A2(n_1299),
.B1(n_1265),
.B2(n_1251),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1250),
.Y(n_1305)
);

CKINVDCx8_ASAP7_75t_R g1306 ( 
.A(n_1246),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1248),
.A2(n_1209),
.B1(n_1299),
.B2(n_1238),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1161),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1151),
.Y(n_1309)
);

BUFx2_ASAP7_75t_SL g1310 ( 
.A(n_1280),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1210),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1209),
.A2(n_1277),
.B1(n_1171),
.B2(n_1297),
.Y(n_1312)
);

INVx8_ASAP7_75t_L g1313 ( 
.A(n_1183),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1261),
.A2(n_1287),
.B1(n_1297),
.B2(n_1203),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1261),
.A2(n_1287),
.B1(n_1203),
.B2(n_1164),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1243),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1295),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1191),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1276),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1155),
.A2(n_1189),
.B1(n_1301),
.B2(n_1247),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1286),
.A2(n_1153),
.B1(n_1196),
.B2(n_1242),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1212),
.A2(n_1170),
.B1(n_1189),
.B2(n_1166),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1269),
.A2(n_1300),
.B1(n_1291),
.B2(n_1278),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1194),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1220),
.Y(n_1325)
);

CKINVDCx6p67_ASAP7_75t_R g1326 ( 
.A(n_1279),
.Y(n_1326)
);

AND2x4_ASAP7_75t_SL g1327 ( 
.A(n_1239),
.B(n_1266),
.Y(n_1327)
);

BUFx12f_ASAP7_75t_L g1328 ( 
.A(n_1259),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1197),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1198),
.Y(n_1330)
);

BUFx4f_ASAP7_75t_SL g1331 ( 
.A(n_1187),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1269),
.A2(n_1300),
.B1(n_1278),
.B2(n_1291),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1272),
.A2(n_1172),
.B1(n_1190),
.B2(n_1158),
.Y(n_1333)
);

INVx6_ASAP7_75t_L g1334 ( 
.A(n_1194),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_1214),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1169),
.A2(n_1225),
.B1(n_1233),
.B2(n_1228),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1194),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1217),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1224),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1262),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1272),
.A2(n_1172),
.B1(n_1190),
.B2(n_1214),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1226),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1260),
.B(n_1235),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1186),
.A2(n_1188),
.B1(n_1233),
.B2(n_1184),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1175),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1177),
.A2(n_1167),
.B1(n_1294),
.B2(n_1285),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1223),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1256),
.A2(n_1294),
.B1(n_1285),
.B2(n_1175),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1240),
.A2(n_1211),
.B1(n_1207),
.B2(n_1256),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1208),
.A2(n_1215),
.B1(n_1213),
.B2(n_1264),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1200),
.A2(n_1215),
.B1(n_1234),
.B2(n_1199),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1228),
.A2(n_1221),
.B1(n_1264),
.B2(n_1282),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1201),
.A2(n_1221),
.B1(n_1292),
.B2(n_1160),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1218),
.A2(n_1219),
.B1(n_1204),
.B2(n_1292),
.Y(n_1354)
);

BUFx8_ASAP7_75t_SL g1355 ( 
.A(n_1157),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1222),
.Y(n_1356)
);

BUFx4f_ASAP7_75t_L g1357 ( 
.A(n_1183),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1231),
.B(n_1198),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1160),
.A2(n_1254),
.B1(n_1205),
.B2(n_1162),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1257),
.A2(n_1290),
.B1(n_1245),
.B2(n_1258),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1274),
.A2(n_1275),
.B1(n_1281),
.B2(n_1293),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1183),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1181),
.A2(n_1257),
.B1(n_1178),
.B2(n_1298),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1216),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1255),
.B(n_1296),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1216),
.Y(n_1366)
);

BUFx2_ASAP7_75t_R g1367 ( 
.A(n_1182),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1181),
.A2(n_1257),
.B1(n_1178),
.B2(n_1193),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1182),
.A2(n_1296),
.B1(n_1268),
.B2(n_1270),
.Y(n_1369)
);

INVx8_ASAP7_75t_L g1370 ( 
.A(n_1268),
.Y(n_1370)
);

CKINVDCx6p67_ASAP7_75t_R g1371 ( 
.A(n_1230),
.Y(n_1371)
);

CKINVDCx16_ASAP7_75t_R g1372 ( 
.A(n_1252),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1252),
.A2(n_1270),
.B1(n_1232),
.B2(n_1229),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1227),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1163),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1173),
.A2(n_1192),
.B1(n_1284),
.B2(n_1263),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1168),
.A2(n_1192),
.B1(n_1249),
.B2(n_1289),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1180),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1176),
.A2(n_1159),
.B1(n_1288),
.B2(n_1237),
.Y(n_1379)
);

BUFx12f_ASAP7_75t_L g1380 ( 
.A(n_1174),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1165),
.A2(n_1244),
.B1(n_1283),
.B2(n_1273),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1192),
.A2(n_1289),
.B1(n_1263),
.B2(n_1284),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1180),
.Y(n_1383)
);

BUFx10_ASAP7_75t_L g1384 ( 
.A(n_1206),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1202),
.B(n_1195),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_SL g1386 ( 
.A1(n_1236),
.A2(n_1271),
.B1(n_1267),
.B2(n_1253),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1263),
.A2(n_1289),
.B1(n_1284),
.B2(n_1202),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1179),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1195),
.A2(n_1179),
.B(n_1241),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1154),
.A2(n_1195),
.B1(n_1156),
.B2(n_1179),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1156),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1156),
.A2(n_1164),
.B1(n_808),
.B2(n_653),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1194),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1164),
.A2(n_808),
.B1(n_653),
.B2(n_1098),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1248),
.A2(n_510),
.B1(n_1209),
.B2(n_1299),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1248),
.A2(n_510),
.B1(n_1209),
.B2(n_1299),
.Y(n_1396)
);

INVx6_ASAP7_75t_L g1397 ( 
.A(n_1194),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1250),
.Y(n_1398)
);

BUFx10_ASAP7_75t_L g1399 ( 
.A(n_1250),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1151),
.Y(n_1400)
);

INVx4_ASAP7_75t_SL g1401 ( 
.A(n_1256),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1152),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1248),
.A2(n_510),
.B1(n_1209),
.B2(n_1299),
.Y(n_1403)
);

INVx4_ASAP7_75t_SL g1404 ( 
.A(n_1256),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1164),
.A2(n_808),
.B1(n_1299),
.B2(n_1287),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1194),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1248),
.A2(n_510),
.B1(n_1209),
.B2(n_1299),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1185),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1185),
.Y(n_1409)
);

NAND2x1p5_ASAP7_75t_L g1410 ( 
.A(n_1194),
.B(n_900),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1151),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1248),
.A2(n_653),
.B(n_852),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1185),
.Y(n_1413)
);

CKINVDCx6p67_ASAP7_75t_R g1414 ( 
.A(n_1151),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1248),
.A2(n_510),
.B1(n_1209),
.B2(n_1299),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1151),
.Y(n_1416)
);

INVx6_ASAP7_75t_L g1417 ( 
.A(n_1194),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1299),
.A2(n_808),
.B1(n_499),
.B2(n_1164),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1254),
.A2(n_877),
.B(n_681),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1151),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1164),
.A2(n_808),
.B1(n_653),
.B2(n_1098),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1185),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1248),
.A2(n_1299),
.B1(n_1261),
.B2(n_1297),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1394),
.B(n_1421),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1323),
.B(n_1332),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1323),
.B(n_1332),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1356),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1356),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1381),
.A2(n_1361),
.B(n_1338),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1381),
.A2(n_1361),
.B(n_1338),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1388),
.Y(n_1431)
);

AOI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1349),
.A2(n_1385),
.B(n_1351),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1307),
.B(n_1341),
.Y(n_1433)
);

AND2x6_ASAP7_75t_L g1434 ( 
.A(n_1365),
.B(n_1388),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1307),
.B(n_1341),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1342),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1378),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1391),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1383),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1355),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1329),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1380),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1371),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1376),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1359),
.A2(n_1389),
.B(n_1353),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1401),
.B(n_1404),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1384),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1418),
.A2(n_1423),
.B1(n_1343),
.B2(n_1320),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1384),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1352),
.B(n_1333),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1379),
.A2(n_1359),
.B(n_1390),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1302),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1387),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1390),
.A2(n_1344),
.B(n_1368),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1387),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1333),
.B(n_1312),
.Y(n_1456)
);

OAI21xp33_ASAP7_75t_L g1457 ( 
.A1(n_1395),
.A2(n_1407),
.B(n_1415),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1316),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1322),
.B(n_1321),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1375),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1402),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1382),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1308),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1339),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1314),
.B(n_1322),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1377),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1312),
.B(n_1353),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1344),
.A2(n_1368),
.B(n_1350),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1347),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1314),
.B(n_1315),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1377),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1354),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1354),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1315),
.B(n_1412),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1324),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1350),
.A2(n_1363),
.B(n_1419),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1324),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1363),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1395),
.B(n_1396),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_L g1480 ( 
.A(n_1396),
.B(n_1403),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1365),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1403),
.B(n_1407),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1304),
.B(n_1415),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1346),
.A2(n_1360),
.B(n_1386),
.Y(n_1484)
);

AO21x1_ASAP7_75t_SL g1485 ( 
.A1(n_1346),
.A2(n_1348),
.B(n_1366),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1405),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1405),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1373),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1327),
.B(n_1311),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1369),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1369),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1392),
.A2(n_1336),
.B1(n_1319),
.B2(n_1335),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1310),
.B(n_1370),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1303),
.B(n_1422),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1334),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_SL g1496 ( 
.A1(n_1358),
.A2(n_1367),
.B(n_1306),
.C(n_1326),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1303),
.B(n_1408),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1334),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1327),
.B(n_1340),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1408),
.B(n_1413),
.Y(n_1500)
);

INVxp67_ASAP7_75t_R g1501 ( 
.A(n_1414),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1409),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1413),
.B(n_1364),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1337),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1372),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1480),
.A2(n_1317),
.B(n_1374),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_SL g1507 ( 
.A1(n_1474),
.A2(n_1420),
.B(n_1309),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1441),
.B(n_1319),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1458),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1452),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1500),
.B(n_1399),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1497),
.Y(n_1512)
);

AOI21xp33_ASAP7_75t_L g1513 ( 
.A1(n_1459),
.A2(n_1370),
.B(n_1411),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1451),
.A2(n_1417),
.B(n_1406),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_SL g1515 ( 
.A1(n_1465),
.A2(n_1416),
.B(n_1370),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1500),
.B(n_1399),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_SL g1517 ( 
.A1(n_1483),
.A2(n_1432),
.B(n_1470),
.Y(n_1517)
);

OR2x2_ASAP7_75t_SL g1518 ( 
.A(n_1460),
.B(n_1318),
.Y(n_1518)
);

AO32x2_ASAP7_75t_L g1519 ( 
.A1(n_1436),
.A2(n_1331),
.A3(n_1393),
.B1(n_1406),
.B2(n_1397),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1503),
.B(n_1362),
.Y(n_1520)
);

O2A1O1Ixp33_ASAP7_75t_SL g1521 ( 
.A1(n_1424),
.A2(n_1400),
.B(n_1345),
.C(n_1397),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1439),
.B(n_1305),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1457),
.A2(n_1357),
.B(n_1330),
.C(n_1313),
.Y(n_1523)
);

OAI211xp5_ASAP7_75t_L g1524 ( 
.A1(n_1448),
.A2(n_1398),
.B(n_1313),
.C(n_1325),
.Y(n_1524)
);

O2A1O1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1479),
.A2(n_1410),
.B(n_1357),
.C(n_1393),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_SL g1526 ( 
.A1(n_1432),
.A2(n_1313),
.B(n_1328),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1484),
.Y(n_1527)
);

BUFx4f_ASAP7_75t_SL g1528 ( 
.A(n_1443),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1482),
.A2(n_1435),
.B(n_1433),
.Y(n_1529)
);

AO32x2_ASAP7_75t_L g1530 ( 
.A1(n_1475),
.A2(n_1477),
.A3(n_1471),
.B1(n_1466),
.B2(n_1462),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1433),
.B(n_1435),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1532)
);

OAI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1476),
.A2(n_1456),
.B(n_1450),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1492),
.A2(n_1443),
.B1(n_1460),
.B2(n_1497),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1451),
.A2(n_1476),
.B(n_1454),
.Y(n_1535)
);

NOR2x1_ASAP7_75t_SL g1536 ( 
.A(n_1460),
.B(n_1485),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1444),
.B(n_1462),
.Y(n_1537)
);

AO22x2_ASAP7_75t_L g1538 ( 
.A1(n_1466),
.A2(n_1471),
.B1(n_1455),
.B2(n_1453),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1437),
.Y(n_1539)
);

NAND2xp33_ASAP7_75t_R g1540 ( 
.A(n_1446),
.B(n_1445),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1502),
.B(n_1463),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1463),
.B(n_1486),
.Y(n_1542)
);

OAI211xp5_ASAP7_75t_L g1543 ( 
.A1(n_1487),
.A2(n_1456),
.B(n_1467),
.C(n_1426),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1437),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1487),
.B(n_1425),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1442),
.A2(n_1489),
.B1(n_1494),
.B2(n_1505),
.Y(n_1546)
);

A2O1A1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1468),
.A2(n_1426),
.B(n_1454),
.C(n_1473),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1447),
.B(n_1449),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1442),
.A2(n_1499),
.B1(n_1446),
.B2(n_1491),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1431),
.B(n_1446),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1427),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1442),
.B(n_1481),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1535),
.B(n_1445),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1527),
.B(n_1478),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1535),
.B(n_1445),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1545),
.B(n_1488),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1510),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1517),
.A2(n_1442),
.B1(n_1445),
.B2(n_1473),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1550),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1535),
.B(n_1472),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1547),
.B(n_1472),
.Y(n_1561)
);

NAND2x1_ASAP7_75t_L g1562 ( 
.A(n_1526),
.B(n_1434),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1531),
.B(n_1481),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1543),
.A2(n_1490),
.B1(n_1491),
.B2(n_1446),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1547),
.B(n_1468),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1533),
.B(n_1429),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1509),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1551),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1519),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1550),
.B(n_1438),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1514),
.B(n_1429),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1529),
.A2(n_1490),
.B1(n_1484),
.B2(n_1434),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1469),
.Y(n_1575)
);

AND2x2_ASAP7_75t_SL g1576 ( 
.A(n_1514),
.B(n_1484),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1538),
.B(n_1469),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1548),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1538),
.B(n_1428),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1519),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1575),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1575),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1554),
.B(n_1577),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1569),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1554),
.B(n_1537),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1577),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1553),
.A2(n_1430),
.B(n_1552),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1568),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1557),
.Y(n_1589)
);

INVx5_ASAP7_75t_SL g1590 ( 
.A(n_1576),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1568),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_L g1592 ( 
.A(n_1564),
.B(n_1440),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1568),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1569),
.B(n_1541),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1579),
.B(n_1512),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1569),
.Y(n_1596)
);

OAI31xp33_ASAP7_75t_L g1597 ( 
.A1(n_1564),
.A2(n_1524),
.A3(n_1534),
.B(n_1521),
.Y(n_1597)
);

NOR3xp33_ASAP7_75t_L g1598 ( 
.A(n_1565),
.B(n_1513),
.C(n_1506),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1578),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1559),
.B(n_1571),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_L g1601 ( 
.A(n_1558),
.B(n_1573),
.C(n_1565),
.Y(n_1601)
);

OR2x2_ASAP7_75t_SL g1602 ( 
.A(n_1556),
.B(n_1508),
.Y(n_1602)
);

INVx5_ASAP7_75t_L g1603 ( 
.A(n_1570),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1579),
.B(n_1532),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1573),
.A2(n_1521),
.B1(n_1542),
.B2(n_1549),
.C(n_1546),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1578),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1574),
.B(n_1537),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1570),
.B(n_1539),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1558),
.A2(n_1523),
.B(n_1525),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1580),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1576),
.B(n_1530),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1530),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1574),
.B(n_1544),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1566),
.B(n_1530),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1588),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1610),
.B(n_1566),
.Y(n_1617)
);

AND2x2_ASAP7_75t_SL g1618 ( 
.A(n_1592),
.B(n_1566),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1583),
.B(n_1563),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1610),
.B(n_1553),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1583),
.B(n_1563),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1606),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1600),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1610),
.B(n_1553),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1581),
.B(n_1582),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1599),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1591),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1581),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1600),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1591),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1593),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1603),
.B(n_1555),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1582),
.B(n_1561),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1586),
.B(n_1561),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1586),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1585),
.B(n_1556),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1585),
.B(n_1561),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1596),
.B(n_1559),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1590),
.B(n_1559),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1614),
.B(n_1560),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1560),
.Y(n_1643)
);

NOR3xp33_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1552),
.C(n_1523),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1555),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1589),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1603),
.B(n_1614),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1603),
.B(n_1555),
.Y(n_1648)
);

NAND4xp25_ASAP7_75t_L g1649 ( 
.A(n_1597),
.B(n_1522),
.C(n_1560),
.D(n_1496),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1603),
.B(n_1572),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1572),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1604),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1613),
.B(n_1567),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1593),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1617),
.B(n_1590),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1653),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1653),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1615),
.Y(n_1658)
);

AOI21xp33_ASAP7_75t_L g1659 ( 
.A1(n_1626),
.A2(n_1601),
.B(n_1597),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1617),
.B(n_1590),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1615),
.Y(n_1661)
);

INVxp33_ASAP7_75t_L g1662 ( 
.A(n_1649),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1647),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1625),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1616),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1647),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1617),
.B(n_1590),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1625),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1634),
.B(n_1602),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1619),
.B(n_1595),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1629),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1634),
.B(n_1602),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1628),
.Y(n_1673)
);

OR2x2_ASAP7_75t_SL g1674 ( 
.A(n_1636),
.B(n_1587),
.Y(n_1674)
);

OAI32xp33_ASAP7_75t_L g1675 ( 
.A1(n_1644),
.A2(n_1611),
.A3(n_1598),
.B1(n_1612),
.B2(n_1609),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1635),
.B(n_1604),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1647),
.B(n_1590),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1622),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1628),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1631),
.Y(n_1680)
);

O2A1O1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1649),
.A2(n_1609),
.B(n_1598),
.C(n_1605),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1619),
.B(n_1595),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1616),
.B(n_1603),
.Y(n_1683)
);

INVx3_ASAP7_75t_SL g1684 ( 
.A(n_1618),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1631),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1621),
.B(n_1611),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1640),
.B(n_1611),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1635),
.B(n_1638),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1632),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1632),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1654),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1638),
.B(n_1608),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1654),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1618),
.A2(n_1605),
.B1(n_1515),
.B2(n_1434),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1652),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1684),
.B(n_1627),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1663),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1689),
.B(n_1626),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1683),
.B(n_1623),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1681),
.B(n_1621),
.Y(n_1702)
);

AOI21xp33_ASAP7_75t_SL g1703 ( 
.A1(n_1662),
.A2(n_1659),
.B(n_1675),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1658),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1658),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1697),
.B(n_1644),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1661),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1683),
.B(n_1618),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1678),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1684),
.B(n_1627),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1671),
.B(n_1637),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1661),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1664),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1669),
.B(n_1637),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1684),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1683),
.Y(n_1716)
);

NOR3xp33_ASAP7_75t_L g1717 ( 
.A(n_1675),
.B(n_1622),
.C(n_1516),
.Y(n_1717)
);

NAND2x1_ASAP7_75t_SL g1718 ( 
.A(n_1677),
.B(n_1655),
.Y(n_1718)
);

OR2x6_ASAP7_75t_L g1719 ( 
.A(n_1665),
.B(n_1493),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1677),
.B(n_1623),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1688),
.B(n_1623),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1664),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1689),
.B(n_1642),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1668),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1669),
.B(n_1612),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1688),
.B(n_1623),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1663),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1672),
.B(n_1642),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1655),
.B(n_1630),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1668),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1660),
.B(n_1667),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1672),
.B(n_1612),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1723),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1705),
.Y(n_1735)
);

OAI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1703),
.A2(n_1696),
.B1(n_1676),
.B2(n_1666),
.C(n_1670),
.Y(n_1736)
);

AOI21xp33_ASAP7_75t_L g1737 ( 
.A1(n_1715),
.A2(n_1657),
.B(n_1656),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1723),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1717),
.A2(n_1702),
.B1(n_1732),
.B2(n_1706),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1732),
.B(n_1660),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1698),
.B(n_1667),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_R g1742 ( 
.A(n_1698),
.B(n_1501),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1709),
.B(n_1666),
.C(n_1695),
.Y(n_1744)
);

O2A1O1Ixp33_ASAP7_75t_SL g1745 ( 
.A1(n_1716),
.A2(n_1695),
.B(n_1682),
.C(n_1686),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1718),
.A2(n_1676),
.B1(n_1693),
.B2(n_1687),
.C(n_1691),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1710),
.B(n_1687),
.Y(n_1747)
);

INVx2_ASAP7_75t_SL g1748 ( 
.A(n_1718),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1710),
.B(n_1693),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1716),
.B(n_1679),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1726),
.A2(n_1633),
.B(n_1648),
.C(n_1645),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1708),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1713),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1721),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1708),
.A2(n_1643),
.B1(n_1630),
.B2(n_1540),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1708),
.B(n_1528),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1713),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1729),
.B(n_1690),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1729),
.B(n_1673),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1741),
.B(n_1720),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1739),
.B(n_1714),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1748),
.A2(n_1674),
.B1(n_1733),
.B2(n_1711),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1742),
.B(n_1700),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1748),
.A2(n_1507),
.B(n_1704),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1734),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1741),
.B(n_1720),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1749),
.B(n_1700),
.Y(n_1767)
);

AOI322xp5_ASAP7_75t_L g1768 ( 
.A1(n_1737),
.A2(n_1624),
.A3(n_1620),
.B1(n_1643),
.B2(n_1633),
.C1(n_1645),
.C2(n_1648),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1756),
.A2(n_1730),
.B1(n_1727),
.B2(n_1721),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1740),
.Y(n_1770)
);

OAI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1747),
.A2(n_1730),
.B(n_1727),
.Y(n_1771)
);

AOI322xp5_ASAP7_75t_L g1772 ( 
.A1(n_1744),
.A2(n_1620),
.A3(n_1624),
.B1(n_1645),
.B2(n_1633),
.C1(n_1648),
.C2(n_1650),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1735),
.Y(n_1773)
);

OAI21xp33_ASAP7_75t_SL g1774 ( 
.A1(n_1752),
.A2(n_1728),
.B(n_1724),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1736),
.B(n_1724),
.Y(n_1775)
);

OAI31xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1746),
.A2(n_1701),
.A3(n_1699),
.B(n_1725),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1740),
.B(n_1738),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1735),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1738),
.B(n_1699),
.Y(n_1779)
);

XOR2xp5_ASAP7_75t_L g1780 ( 
.A(n_1761),
.B(n_1769),
.Y(n_1780)
);

OAI321xp33_ASAP7_75t_L g1781 ( 
.A1(n_1775),
.A2(n_1755),
.A3(n_1757),
.B1(n_1743),
.B2(n_1753),
.C(n_1750),
.Y(n_1781)
);

NOR2x1_ASAP7_75t_L g1782 ( 
.A(n_1773),
.B(n_1743),
.Y(n_1782)
);

INVxp33_ASAP7_75t_L g1783 ( 
.A(n_1763),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1760),
.B(n_1754),
.Y(n_1784)
);

A2O1A1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1776),
.A2(n_1751),
.B(n_1754),
.C(n_1758),
.Y(n_1785)
);

AOI211xp5_ASAP7_75t_L g1786 ( 
.A1(n_1774),
.A2(n_1745),
.B(n_1757),
.C(n_1753),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1777),
.B(n_1758),
.C(n_1759),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1770),
.B(n_1766),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1762),
.A2(n_1759),
.B1(n_1728),
.B2(n_1731),
.C(n_1722),
.Y(n_1789)
);

INVxp67_ASAP7_75t_SL g1790 ( 
.A(n_1765),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1765),
.Y(n_1791)
);

NAND4xp25_ASAP7_75t_L g1792 ( 
.A(n_1787),
.B(n_1764),
.C(n_1771),
.D(n_1767),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1781),
.B(n_1764),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1783),
.B(n_1779),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1790),
.B(n_1778),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1791),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1784),
.B(n_1768),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1782),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1788),
.Y(n_1799)
);

OAI211xp5_ASAP7_75t_L g1800 ( 
.A1(n_1786),
.A2(n_1772),
.B(n_1712),
.C(n_1707),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1780),
.Y(n_1801)
);

OAI211xp5_ASAP7_75t_L g1802 ( 
.A1(n_1793),
.A2(n_1785),
.B(n_1789),
.C(n_1781),
.Y(n_1802)
);

NAND4xp25_ASAP7_75t_L g1803 ( 
.A(n_1801),
.B(n_1701),
.C(n_1511),
.D(n_1501),
.Y(n_1803)
);

NOR3xp33_ASAP7_75t_L g1804 ( 
.A(n_1794),
.B(n_1701),
.C(n_1520),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1797),
.A2(n_1719),
.B1(n_1528),
.B2(n_1680),
.Y(n_1805)
);

AOI221x1_ASAP7_75t_L g1806 ( 
.A1(n_1798),
.A2(n_1673),
.B1(n_1694),
.B2(n_1680),
.C(n_1685),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_SL g1807 ( 
.A1(n_1803),
.A2(n_1792),
.B1(n_1799),
.B2(n_1795),
.C(n_1796),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1802),
.B(n_1800),
.Y(n_1808)
);

NAND2xp33_ASAP7_75t_SL g1809 ( 
.A(n_1806),
.B(n_1800),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1804),
.A2(n_1694),
.B1(n_1685),
.B2(n_1650),
.C(n_1651),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1805),
.A2(n_1651),
.B(n_1650),
.C(n_1674),
.Y(n_1811)
);

OAI211xp5_ASAP7_75t_L g1812 ( 
.A1(n_1802),
.A2(n_1651),
.B(n_1692),
.C(n_1562),
.Y(n_1812)
);

INVx2_ASAP7_75t_SL g1813 ( 
.A(n_1808),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1809),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1807),
.B(n_1719),
.Y(n_1815)
);

AO22x2_ASAP7_75t_L g1816 ( 
.A1(n_1812),
.A2(n_1692),
.B1(n_1630),
.B2(n_1646),
.Y(n_1816)
);

XOR2x2_ASAP7_75t_L g1817 ( 
.A(n_1811),
.B(n_1536),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1814),
.Y(n_1818)
);

AO22x2_ASAP7_75t_L g1819 ( 
.A1(n_1813),
.A2(n_1810),
.B1(n_1630),
.B2(n_1641),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_SL g1820 ( 
.A1(n_1815),
.A2(n_1719),
.B1(n_1518),
.B2(n_1493),
.Y(n_1820)
);

XOR2x2_ASAP7_75t_L g1821 ( 
.A(n_1818),
.B(n_1817),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1821),
.B(n_1719),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1822),
.A2(n_1820),
.B1(n_1816),
.B2(n_1819),
.Y(n_1823)
);

OAI22x1_ASAP7_75t_L g1824 ( 
.A1(n_1822),
.A2(n_1641),
.B1(n_1639),
.B2(n_1596),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1823),
.B(n_1641),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1824),
.A2(n_1641),
.B1(n_1624),
.B2(n_1620),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1825),
.A2(n_1641),
.B1(n_1599),
.B2(n_1639),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1826),
.B(n_1639),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1493),
.B(n_1562),
.Y(n_1829)
);

A2O1A1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1829),
.A2(n_1827),
.B(n_1639),
.C(n_1613),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1830),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1831),
.A2(n_1639),
.B1(n_1584),
.B2(n_1607),
.C(n_1594),
.Y(n_1832)
);

AOI211xp5_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1498),
.B(n_1495),
.C(n_1504),
.Y(n_1833)
);


endmodule