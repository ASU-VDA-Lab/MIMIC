module fake_jpeg_29309_n_465 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_465);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_465;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_52),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_27),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_58),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_61),
.B(n_98),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_13),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_66),
.B(n_74),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_67),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_69),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_10),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_82),
.Y(n_155)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_42),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_6),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_19),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_92),
.B(n_46),
.Y(n_137)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_14),
.B(n_6),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_44),
.Y(n_150)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_39),
.B1(n_36),
.B2(n_41),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_102),
.A2(n_110),
.B1(n_131),
.B2(n_134),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_48),
.B(n_33),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_107),
.B(n_138),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_36),
.B1(n_41),
.B2(n_46),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_133),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_124),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_84),
.A2(n_18),
.B1(n_41),
.B2(n_37),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_90),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_64),
.A2(n_18),
.B1(n_41),
.B2(n_37),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

INVx2_ASAP7_75t_R g138 ( 
.A(n_55),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_37),
.B1(n_34),
.B2(n_46),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_72),
.B1(n_97),
.B2(n_96),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_32),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_49),
.B(n_44),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_43),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

CKINVDCx12_ASAP7_75t_R g175 ( 
.A(n_158),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_50),
.A2(n_32),
.B1(n_23),
.B2(n_46),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_88),
.B1(n_71),
.B2(n_68),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_77),
.A2(n_7),
.B(n_48),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_23),
.Y(n_173)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_38),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_168),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_167),
.A2(n_122),
.B1(n_104),
.B2(n_147),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_47),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

CKINVDCx12_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_47),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_190),
.Y(n_237)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

BUFx4f_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_181),
.Y(n_223)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_105),
.B(n_91),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_188),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_194),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_78),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_187),
.B(n_123),
.C(n_106),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_118),
.B(n_99),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_38),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_191),
.B(n_197),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_155),
.B(n_33),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_134),
.A2(n_93),
.B1(n_83),
.B2(n_52),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_193),
.A2(n_196),
.B1(n_199),
.B2(n_204),
.Y(n_227)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_129),
.B(n_75),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_124),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_43),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_198),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_145),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_201),
.Y(n_238)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_143),
.A2(n_54),
.B1(n_85),
.B2(n_79),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_202),
.A2(n_207),
.B1(n_102),
.B2(n_62),
.Y(n_214)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_208),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_131),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_205),
.B(n_122),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_72),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_123),
.B(n_87),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_139),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_209),
.B(n_210),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_214),
.A2(n_170),
.B1(n_196),
.B2(n_169),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_176),
.A2(n_143),
.B1(n_154),
.B2(n_109),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_217),
.B1(n_220),
.B2(n_225),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_183),
.B1(n_166),
.B2(n_178),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_147),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_195),
.C(n_194),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_144),
.B1(n_154),
.B2(n_130),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_109),
.B1(n_136),
.B2(n_130),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_240),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_136),
.B1(n_110),
.B2(n_161),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_231),
.B1(n_235),
.B2(n_164),
.Y(n_250)
);

AO22x1_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_181),
.B1(n_175),
.B2(n_140),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_165),
.A2(n_127),
.B1(n_125),
.B2(n_120),
.Y(n_235)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_190),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_252),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_251),
.B1(n_260),
.B2(n_267),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_217),
.A2(n_191),
.B1(n_163),
.B2(n_174),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_187),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_195),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_257),
.Y(n_284)
);

INVx5_ASAP7_75t_SL g254 ( 
.A(n_241),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_255),
.A2(n_244),
.B1(n_223),
.B2(n_234),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_233),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_209),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_259),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_203),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_214),
.A2(n_198),
.B1(n_172),
.B2(n_180),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

OA21x2_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_181),
.B(n_124),
.Y(n_299)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_31),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_227),
.A2(n_127),
.B1(n_125),
.B2(n_171),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_231),
.A2(n_104),
.B1(n_140),
.B2(n_182),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_211),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_31),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_273),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_228),
.A2(n_127),
.B1(n_152),
.B2(n_201),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_218),
.B1(n_223),
.B2(n_241),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_205),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_229),
.C(n_242),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_220),
.B(n_216),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_276),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_218),
.B1(n_240),
.B2(n_216),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_278),
.A2(n_283),
.B1(n_261),
.B2(n_253),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_282),
.A2(n_296),
.B1(n_268),
.B2(n_280),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_218),
.B1(n_226),
.B2(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_238),
.B(n_222),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_299),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_255),
.A2(n_234),
.B1(n_219),
.B2(n_244),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_260),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_291),
.B(n_271),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_250),
.A2(n_244),
.B1(n_221),
.B2(n_242),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_302),
.B(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_257),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_310),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_316),
.C(n_324),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_292),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_275),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_259),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_311),
.B(n_312),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_287),
.B(n_249),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_319),
.B1(n_276),
.B2(n_289),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_266),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_295),
.B(n_273),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_317),
.B(n_318),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_251),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_292),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_325),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_258),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_321),
.B(n_323),
.Y(n_344)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_281),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_322),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_262),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_252),
.C(n_270),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_263),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_293),
.B1(n_283),
.B2(n_278),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_329),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_277),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_308),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_280),
.B1(n_282),
.B2(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_303),
.A2(n_305),
.B1(n_313),
.B2(n_319),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_336),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_313),
.A2(n_299),
.B(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_338),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_303),
.A2(n_290),
.B1(n_286),
.B2(n_280),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_313),
.A2(n_299),
.B(n_291),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_299),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_339),
.Y(n_355)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_323),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_340),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_305),
.A2(n_311),
.B1(n_290),
.B2(n_316),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_341),
.A2(n_345),
.B1(n_349),
.B2(n_326),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_317),
.A2(n_267),
.B1(n_306),
.B2(n_274),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_309),
.A2(n_282),
.B1(n_292),
.B2(n_294),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_358),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_328),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_359),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_339),
.A2(n_343),
.B(n_351),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_357),
.A2(n_349),
.B(n_346),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_324),
.C(n_325),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_324),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_310),
.C(n_318),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_370),
.C(n_375),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_307),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_361),
.Y(n_377)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_331),
.Y(n_362)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_362),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_363),
.A2(n_336),
.B1(n_347),
.B2(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_365),
.Y(n_391)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_372),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_339),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_342),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_321),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_348),
.B(n_344),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_371),
.B(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_347),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_322),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_315),
.C(n_302),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_376),
.B(n_370),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_366),
.A2(n_338),
.B(n_335),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_380),
.Y(n_398)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_382),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_374),
.B(n_236),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_390),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_387),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_346),
.C(n_342),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_392),
.C(n_394),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_355),
.B1(n_368),
.B2(n_354),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_359),
.B(n_304),
.C(n_294),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_356),
.A2(n_320),
.B1(n_297),
.B2(n_301),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_393),
.A2(n_363),
.B1(n_368),
.B2(n_369),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_297),
.C(n_301),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_375),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_402),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_388),
.B(n_377),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_400),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_406),
.Y(n_413)
);

BUFx12f_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

FAx1_ASAP7_75t_SL g411 ( 
.A(n_401),
.B(n_379),
.CI(n_386),
.CON(n_411),
.SN(n_411)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_360),
.Y(n_402)
);

INVx5_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_404),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_352),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_378),
.C(n_385),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_393),
.A2(n_354),
.B1(n_355),
.B2(n_371),
.Y(n_409)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_382),
.A2(n_357),
.B1(n_299),
.B2(n_292),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_410),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_415),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_394),
.C(n_381),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_416),
.C(n_424),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_387),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_386),
.C(n_389),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_245),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_400),
.A2(n_391),
.B(n_385),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_272),
.B(n_229),
.Y(n_435)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_391),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_422),
.B(n_407),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_398),
.C(n_401),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_427),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_404),
.B1(n_400),
.B2(n_405),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_426),
.B(n_430),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_420),
.A2(n_300),
.B1(n_248),
.B2(n_247),
.Y(n_427)
);

OA22x2_ASAP7_75t_L g428 ( 
.A1(n_415),
.A2(n_421),
.B1(n_413),
.B2(n_422),
.Y(n_428)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_428),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_423),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_269),
.Y(n_431)
);

NOR4xp25_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_436),
.C(n_411),
.D(n_413),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_300),
.B(n_265),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_433),
.A2(n_435),
.B(n_164),
.Y(n_442)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_412),
.Y(n_434)
);

AOI21xp33_ASAP7_75t_L g444 ( 
.A1(n_434),
.A2(n_254),
.B(n_221),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_439),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_414),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_429),
.A2(n_416),
.B(n_245),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_442),
.Y(n_451)
);

AOI322xp5_ASAP7_75t_L g448 ( 
.A1(n_444),
.A2(n_446),
.A3(n_185),
.B1(n_186),
.B2(n_116),
.C1(n_152),
.C2(n_434),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_429),
.A2(n_221),
.B(n_230),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_445),
.B(n_432),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_428),
.A2(n_254),
.B1(n_185),
.B2(n_186),
.Y(n_446)
);

AO21x1_ASAP7_75t_L g455 ( 
.A1(n_447),
.A2(n_448),
.B(n_450),
.Y(n_455)
);

AOI322xp5_ASAP7_75t_L g450 ( 
.A1(n_437),
.A2(n_441),
.A3(n_428),
.B1(n_446),
.B2(n_425),
.C1(n_443),
.C2(n_185),
.Y(n_450)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_70),
.B1(n_65),
.B2(n_56),
.Y(n_453)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_453),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_449),
.A2(n_451),
.B(n_53),
.Y(n_454)
);

AOI21x1_ASAP7_75t_SL g458 ( 
.A1(n_454),
.A2(n_456),
.B(n_0),
.Y(n_458)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_0),
.C(n_1),
.Y(n_456)
);

AOI21xp33_ASAP7_75t_L g461 ( 
.A1(n_458),
.A2(n_459),
.B(n_1),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_455),
.B(n_1),
.Y(n_459)
);

BUFx24_ASAP7_75t_SL g460 ( 
.A(n_457),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_460),
.B(n_461),
.C(n_1),
.Y(n_462)
);

OAI221xp5_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_3),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_464),
.A2(n_3),
.B1(n_4),
.B2(n_342),
.Y(n_465)
);


endmodule