module fake_jpeg_928_n_119 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_3),
.B(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_29),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_39),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_34),
.B1(n_38),
.B2(n_36),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_35),
.B(n_38),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_68),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_33),
.B(n_34),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_67),
.B1(n_4),
.B2(n_5),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_46),
.B1(n_44),
.B2(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_59),
.B1(n_53),
.B2(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_82),
.B1(n_7),
.B2(n_8),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_2),
.C(n_3),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_59),
.C(n_58),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_21),
.C(n_28),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_81),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_2),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_6),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_4),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_58),
.B1(n_35),
.B2(n_6),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_13),
.B(n_14),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_91),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_12),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_16),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_77),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_17),
.C(n_27),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_78),
.C(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_23),
.C(n_26),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_95),
.C(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_86),
.B1(n_85),
.B2(n_92),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_108),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_99),
.C(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_110),
.B(n_111),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_97),
.C(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_112),
.A2(n_109),
.B1(n_101),
.B2(n_108),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_103),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_113),
.B(n_24),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_30),
.C(n_15),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_13),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_15),
.Y(n_119)
);


endmodule