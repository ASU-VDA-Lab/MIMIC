module fake_aes_7974_n_719 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_719);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_719;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_71), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_38), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_49), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_67), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_29), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_65), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_24), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_6), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_43), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_3), .Y(n_90) );
BUFx8_ASAP7_75t_SL g91 ( .A(n_18), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_42), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
BUFx2_ASAP7_75t_L g96 ( .A(n_54), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_33), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_68), .Y(n_98) );
INVxp33_ASAP7_75t_L g99 ( .A(n_77), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_45), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_37), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_28), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_76), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_62), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_2), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_34), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_17), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_60), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_36), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_53), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_1), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_11), .Y(n_113) );
BUFx5_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
BUFx5_ASAP7_75t_L g115 ( .A(n_27), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_41), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_32), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_46), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_57), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_19), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_21), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_22), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_64), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_59), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_31), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_56), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_2), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_3), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_114), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_91), .Y(n_130) );
AO22x1_ASAP7_75t_L g131 ( .A1(n_99), .A2(n_0), .B1(n_1), .B2(n_4), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_99), .B(n_103), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_96), .B(n_0), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_112), .B(n_4), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_103), .B(n_5), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_114), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_90), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_87), .B(n_5), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_90), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_128), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_128), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_88), .Y(n_146) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_95), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_114), .B(n_6), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_91), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_82), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_80), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
INVx1_ASAP7_75t_SL g155 ( .A(n_82), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_115), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_115), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_86), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_102), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_92), .B(n_7), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_93), .B(n_48), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_98), .B(n_8), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_101), .Y(n_167) );
XOR2xp5_ASAP7_75t_L g168 ( .A(n_102), .B(n_8), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_84), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_81), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_105), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_125), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_135), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_164), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_132), .B(n_120), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_140), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_132), .B(n_124), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_164), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_134), .B(n_110), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_171), .B(n_107), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_163), .B(n_153), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_137), .B(n_113), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_152), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_136), .B(n_117), .Y(n_184) );
OR2x2_ASAP7_75t_L g185 ( .A(n_147), .B(n_122), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_135), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_163), .B(n_115), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_153), .B(n_123), .Y(n_190) );
NOR2xp33_ASAP7_75t_SL g191 ( .A(n_130), .B(n_85), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_136), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_170), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_154), .B(n_121), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_154), .B(n_89), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_137), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_160), .B(n_97), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_160), .B(n_115), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_129), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_129), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_165), .B(n_119), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_155), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_130), .B(n_116), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_156), .B(n_118), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_150), .B(n_165), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_162), .B(n_115), .Y(n_209) );
OR2x2_ASAP7_75t_L g210 ( .A(n_150), .B(n_104), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
NOR2x1p5_ASAP7_75t_L g212 ( .A(n_169), .B(n_100), .Y(n_212) );
BUFx3_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_151), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_142), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g216 ( .A(n_133), .B(n_109), .C(n_108), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_151), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_165), .B(n_111), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_131), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_170), .B(n_106), .Y(n_220) );
AO22x2_ASAP7_75t_L g221 ( .A1(n_168), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_141), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_166), .B(n_115), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_143), .B(n_12), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_169), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_151), .B(n_13), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_162), .B(n_52), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_161), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_138), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_144), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_162), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_162), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_162), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_145), .B(n_14), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_224), .Y(n_236) );
NAND3xp33_ASAP7_75t_SL g237 ( .A(n_229), .B(n_159), .C(n_157), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_208), .B(n_164), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
INVx5_ASAP7_75t_L g240 ( .A(n_184), .Y(n_240) );
AND2x6_ASAP7_75t_SL g241 ( .A(n_176), .B(n_168), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_204), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_175), .B(n_203), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_234), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_192), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_203), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_175), .B(n_164), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_197), .A2(n_164), .B1(n_144), .B2(n_172), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_177), .B(n_131), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_235), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_232), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_195), .A2(n_157), .B1(n_159), .B2(n_167), .Y(n_255) );
AND2x6_ASAP7_75t_L g256 ( .A(n_178), .B(n_167), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_181), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_182), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_218), .B(n_172), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_184), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_218), .B(n_172), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_174), .B(n_167), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_190), .B(n_172), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_196), .B(n_172), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_181), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_198), .B(n_167), .Y(n_266) );
NOR2xp33_ASAP7_75t_R g267 ( .A(n_225), .B(n_15), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_193), .B(n_167), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_180), .B(n_16), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_206), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_178), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_184), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_188), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_213), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_185), .B(n_158), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_226), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_212), .B(n_16), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_194), .A2(n_158), .B(n_149), .C(n_146), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_179), .B(n_149), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_194), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_184), .A2(n_158), .B1(n_149), .B2(n_146), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_223), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_200), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_184), .A2(n_158), .B1(n_149), .B2(n_146), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_213), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_179), .B(n_149), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
BUFx4f_ASAP7_75t_L g291 ( .A(n_205), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_216), .B(n_158), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_210), .B(n_20), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_215), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_174), .B(n_23), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_200), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_220), .B(n_138), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_220), .B(n_138), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_186), .B(n_146), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_186), .B(n_146), .Y(n_300) );
NOR3xp33_ASAP7_75t_SL g301 ( .A(n_222), .B(n_26), .C(n_30), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_209), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_201), .B(n_138), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_283), .A2(n_202), .B(n_173), .C(n_187), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_242), .A2(n_191), .B1(n_221), .B2(n_217), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_290), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_299), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_260), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_260), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_240), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
OAI21x1_ASAP7_75t_SL g313 ( .A1(n_274), .A2(n_173), .B(n_187), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_258), .B(n_183), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_238), .A2(n_214), .B(n_209), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_249), .A2(n_211), .B(n_199), .Y(n_318) );
CKINVDCx14_ASAP7_75t_R g319 ( .A(n_294), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_240), .Y(n_320) );
INVx4_ASAP7_75t_SL g321 ( .A(n_256), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_241), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_252), .A2(n_211), .B(n_199), .C(n_231), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_272), .B(n_228), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_246), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_248), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
BUFx6f_ASAP7_75t_SL g328 ( .A(n_280), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_240), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_237), .A2(n_228), .B(n_221), .C(n_47), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_258), .B(n_39), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_248), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_270), .B(n_221), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_246), .B(n_230), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_243), .B(n_40), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_244), .B(n_50), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_247), .B(n_51), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_236), .A2(n_230), .B1(n_227), .B2(n_61), .Y(n_338) );
INVx4_ASAP7_75t_L g339 ( .A(n_285), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_291), .B(n_55), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_271), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_250), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_250), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_278), .B(n_58), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_268), .Y(n_345) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_237), .B(n_230), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_239), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_259), .A2(n_230), .B(n_227), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_253), .A2(n_265), .B(n_257), .C(n_266), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_236), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_271), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_273), .B(n_63), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_282), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_289), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_256), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_267), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_346), .A2(n_261), .B(n_298), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_316), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_312), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_333), .A2(n_280), .B1(n_269), .B2(n_293), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_309), .B(n_295), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_353), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_325), .B(n_293), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_354), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_304), .Y(n_366) );
INVx6_ASAP7_75t_L g367 ( .A(n_339), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_325), .B(n_275), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_349), .A2(n_264), .B(n_263), .C(n_255), .Y(n_369) );
AOI21x1_ASAP7_75t_L g370 ( .A1(n_348), .A2(n_297), .B(n_303), .Y(n_370) );
O2A1O1Ixp33_ASAP7_75t_SL g371 ( .A1(n_335), .A2(n_281), .B(n_292), .C(n_262), .Y(n_371) );
INVx2_ASAP7_75t_SL g372 ( .A(n_309), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_307), .A2(n_291), .B1(n_268), .B2(n_267), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_342), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_301), .B(n_251), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_343), .B(n_295), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_347), .B(n_286), .Y(n_378) );
OAI21x1_ASAP7_75t_SL g379 ( .A1(n_313), .A2(n_251), .B(n_296), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_305), .B(n_301), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_287), .B(n_284), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_330), .A2(n_266), .B(n_300), .Y(n_382) );
AOI22xp33_ASAP7_75t_SL g383 ( .A1(n_328), .A2(n_256), .B1(n_288), .B2(n_271), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_315), .A2(n_318), .B(n_335), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_350), .B(n_332), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_352), .A2(n_287), .B(n_284), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_356), .B(n_302), .Y(n_387) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_337), .A2(n_344), .B(n_318), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_317), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_337), .A2(n_279), .B(n_254), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_364), .A2(n_322), .B1(n_339), .B2(n_314), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_364), .B(n_345), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_359), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_359), .A2(n_355), .B1(n_340), .B2(n_331), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_380), .A2(n_328), .B1(n_361), .B2(n_377), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_370), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_363), .Y(n_397) );
INVx3_ASAP7_75t_L g398 ( .A(n_389), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_384), .A2(n_315), .B(n_344), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_373), .A2(n_319), .B(n_330), .C(n_326), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_336), .B1(n_324), .B2(n_323), .C(n_338), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_360), .A2(n_334), .B1(n_306), .B2(n_308), .C(n_324), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_370), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_380), .A2(n_310), .B1(n_317), .B2(n_355), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_371), .A2(n_351), .B(n_341), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_365), .A2(n_329), .B(n_327), .C(n_320), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_365), .A2(n_245), .B(n_320), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_387), .A2(n_310), .B1(n_329), .B2(n_327), .C(n_311), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_368), .A2(n_317), .B1(n_311), .B2(n_351), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_377), .A2(n_256), .B1(n_341), .B2(n_351), .Y(n_414) );
INVxp33_ASAP7_75t_SL g415 ( .A(n_383), .Y(n_415) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_387), .A2(n_341), .B1(n_288), .B2(n_276), .C(n_271), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g417 ( .A1(n_358), .A2(n_256), .B(n_321), .Y(n_417) );
AO31x2_ASAP7_75t_L g418 ( .A1(n_366), .A2(n_321), .A3(n_227), .B(n_70), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_377), .B(n_389), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_393), .Y(n_420) );
BUFx6f_ASAP7_75t_SL g421 ( .A(n_419), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_413), .B(n_366), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_415), .A2(n_377), .B1(n_376), .B2(n_382), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_397), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_413), .B(n_389), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_398), .B(n_357), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_397), .B(n_376), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_401), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_396), .Y(n_430) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_405), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_401), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_410), .B(n_376), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_419), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_419), .B(n_376), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_392), .B(n_382), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_418), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_398), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_398), .B(n_382), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_418), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_395), .B(n_388), .Y(n_442) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_399), .A2(n_390), .B(n_379), .Y(n_443) );
INVx4_ASAP7_75t_L g444 ( .A(n_392), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_404), .B(n_368), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_418), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_418), .B(n_388), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_418), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_408), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_417), .B(n_388), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_394), .B(n_378), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_416), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_403), .B(n_378), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_444), .B(n_391), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_425), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_429), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_436), .B(n_388), .Y(n_460) );
NAND4xp25_ASAP7_75t_SL g461 ( .A(n_420), .B(n_415), .C(n_406), .D(n_414), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_444), .B(n_385), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_430), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_430), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_429), .B(n_385), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_445), .B(n_367), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_444), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_436), .B(n_357), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_436), .B(n_357), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_426), .Y(n_470) );
NOR3xp33_ASAP7_75t_SL g471 ( .A(n_452), .B(n_400), .C(n_402), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_428), .B(n_357), .Y(n_472) );
INVx3_ASAP7_75t_L g473 ( .A(n_426), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_424), .B(n_369), .C(n_407), .D(n_367), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_432), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_444), .B(n_412), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_428), .B(n_390), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_435), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_428), .B(n_372), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_442), .B(n_372), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_422), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_449), .B(n_362), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_442), .B(n_362), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g488 ( .A1(n_444), .A2(n_367), .B1(n_362), .B2(n_379), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_435), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_433), .B(n_367), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_442), .B(n_66), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_420), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_422), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_433), .B(n_69), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_452), .A2(n_386), .B1(n_381), .B2(n_321), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_433), .B(n_72), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_422), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_431), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_437), .B(n_386), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_431), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_440), .B(n_73), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_437), .B(n_381), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_440), .B(n_75), .Y(n_503) );
OAI211xp5_ASAP7_75t_SL g504 ( .A1(n_445), .A2(n_78), .B(n_79), .C(n_227), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_440), .B(n_276), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_457), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_457), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_458), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_467), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_463), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_462), .B(n_445), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_460), .B(n_451), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_462), .B(n_434), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_467), .B(n_449), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_460), .B(n_451), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_458), .B(n_434), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_467), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_459), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_459), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_472), .B(n_451), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_475), .B(n_434), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_467), .B(n_423), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_475), .B(n_434), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_463), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_485), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_485), .B(n_434), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_500), .B(n_447), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_479), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_472), .B(n_447), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_482), .B(n_447), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_492), .B(n_455), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_492), .B(n_455), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_479), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_482), .B(n_423), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_500), .B(n_423), .Y(n_537) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_476), .B(n_439), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_489), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_466), .B(n_454), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_464), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_489), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_466), .B(n_454), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_489), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_490), .B(n_423), .Y(n_545) );
OR2x6_ASAP7_75t_L g546 ( .A(n_483), .B(n_448), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_465), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_465), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_468), .B(n_423), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_498), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_498), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_468), .B(n_446), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_469), .B(n_446), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_461), .A2(n_454), .B1(n_421), .B2(n_453), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_469), .B(n_441), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_488), .A2(n_453), .B(n_441), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_461), .A2(n_421), .B1(n_453), .B2(n_424), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_486), .B(n_438), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_486), .B(n_438), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_481), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_478), .B(n_481), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_456), .B(n_439), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_478), .B(n_448), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_471), .A2(n_448), .B1(n_438), .B2(n_450), .C(n_427), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_557), .A2(n_456), .B1(n_476), .B2(n_471), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_506), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_561), .B(n_487), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_528), .B(n_490), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_561), .B(n_473), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_528), .B(n_483), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_529), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_512), .B(n_483), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_512), .B(n_497), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_547), .B(n_497), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_548), .B(n_499), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_530), .B(n_470), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_470), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_509), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_550), .B(n_499), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_521), .B(n_470), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_521), .B(n_470), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_506), .Y(n_582) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_518), .B(n_488), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_509), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_516), .B(n_487), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_518), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_507), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_523), .B(n_480), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_507), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_526), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_516), .B(n_487), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_550), .B(n_502), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g595 ( .A1(n_515), .A2(n_484), .B(n_504), .C(n_494), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_551), .B(n_532), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_560), .B(n_480), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_551), .B(n_502), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_511), .B(n_493), .Y(n_599) );
OR2x6_ASAP7_75t_L g600 ( .A(n_538), .B(n_480), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_533), .B(n_493), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_519), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_531), .B(n_545), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_537), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_520), .B(n_493), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_549), .B(n_473), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_529), .B(n_477), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_517), .Y(n_608) );
NAND3xp33_ASAP7_75t_SL g609 ( .A(n_554), .B(n_496), .C(n_494), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_534), .B(n_477), .Y(n_610) );
AOI221x1_ASAP7_75t_L g611 ( .A1(n_556), .A2(n_504), .B1(n_474), .B2(n_491), .C(n_501), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_535), .B(n_477), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_549), .B(n_473), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_537), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_531), .B(n_464), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_540), .B(n_421), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_539), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_600), .A2(n_538), .B1(n_523), .B2(n_543), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_596), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_596), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_573), .B(n_563), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_609), .A2(n_538), .B1(n_546), .B2(n_514), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_608), .B(n_552), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_593), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_603), .B(n_562), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_583), .A2(n_523), .B(n_546), .Y(n_627) );
NOR4xp25_ASAP7_75t_L g628 ( .A(n_595), .B(n_564), .C(n_474), .D(n_524), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_618), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_595), .A2(n_527), .B(n_495), .C(n_545), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_584), .Y(n_631) );
OAI322xp33_ASAP7_75t_SL g632 ( .A1(n_575), .A2(n_542), .A3(n_544), .B1(n_525), .B2(n_541), .C1(n_510), .C2(n_513), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_578), .Y(n_633) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_565), .A2(n_546), .B1(n_495), .B2(n_553), .C(n_552), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_616), .B(n_563), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_604), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_611), .A2(n_496), .B(n_491), .Y(n_637) );
AOI221x1_ASAP7_75t_L g638 ( .A1(n_565), .A2(n_503), .B1(n_501), .B2(n_427), .C(n_450), .Y(n_638) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_586), .A2(n_546), .B1(n_555), .B2(n_553), .C(n_487), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_572), .B(n_555), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_602), .Y(n_641) );
AOI21xp33_ASAP7_75t_SL g642 ( .A1(n_600), .A2(n_503), .B(n_536), .Y(n_642) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_567), .A2(n_559), .B(n_558), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_588), .B(n_513), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_566), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_615), .B(n_536), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g647 ( .A1(n_574), .A2(n_473), .B1(n_541), .B2(n_525), .C(n_510), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_613), .B(n_559), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_582), .Y(n_649) );
AOI221xp5_ASAP7_75t_SL g650 ( .A1(n_575), .A2(n_558), .B1(n_505), .B2(n_464), .C(n_421), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_617), .A2(n_421), .B1(n_427), .B2(n_505), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_587), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_574), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_597), .B(n_427), .C(n_426), .D(n_443), .Y(n_654) );
OAI32xp33_ASAP7_75t_L g655 ( .A1(n_570), .A2(n_427), .A3(n_426), .B1(n_443), .B2(n_276), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_579), .B(n_443), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_588), .A2(n_443), .B1(n_276), .B2(n_288), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_629), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_620), .B(n_594), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_636), .B(n_569), .Y(n_660) );
NAND2x1_ASAP7_75t_L g661 ( .A(n_627), .B(n_600), .Y(n_661) );
AOI22xp5_ASAP7_75t_SL g662 ( .A1(n_636), .A2(n_619), .B1(n_629), .B2(n_653), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_621), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_634), .A2(n_614), .B1(n_606), .B2(n_576), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_630), .A2(n_623), .B(n_628), .C(n_642), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_625), .Y(n_666) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_644), .B(n_633), .Y(n_667) );
NAND2xp33_ASAP7_75t_R g668 ( .A(n_637), .B(n_585), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_631), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_635), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_641), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_645), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_L g673 ( .A1(n_654), .A2(n_577), .B(n_591), .C(n_580), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_622), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_630), .B(n_594), .C(n_598), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_649), .Y(n_676) );
OAI31xp33_ASAP7_75t_SL g677 ( .A1(n_623), .A2(n_581), .A3(n_589), .B(n_590), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_653), .B(n_598), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_626), .A2(n_568), .B1(n_579), .B2(n_592), .Y(n_679) );
AO22x1_ASAP7_75t_L g680 ( .A1(n_632), .A2(n_571), .B1(n_605), .B2(n_607), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_652), .Y(n_681) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_669), .Y(n_682) );
XNOR2xp5_ASAP7_75t_L g683 ( .A(n_664), .B(n_624), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_668), .A2(n_639), .B1(n_643), .B2(n_650), .Y(n_684) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_661), .B(n_647), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_675), .B(n_648), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_662), .A2(n_640), .B1(n_646), .B2(n_651), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_658), .Y(n_688) );
AOI211xp5_ASAP7_75t_SL g689 ( .A1(n_673), .A2(n_669), .B(n_665), .C(n_678), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_665), .A2(n_656), .B(n_655), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_667), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_680), .A2(n_638), .B(n_605), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_677), .A2(n_601), .B(n_599), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_672), .Y(n_694) );
AOI21xp5_ASAP7_75t_SL g695 ( .A1(n_667), .A2(n_657), .B(n_607), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_685), .B(n_660), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_689), .A2(n_679), .B1(n_659), .B2(n_663), .C(n_671), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_686), .B(n_659), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_694), .Y(n_699) );
OAI221xp5_ASAP7_75t_SL g700 ( .A1(n_684), .A2(n_674), .B1(n_670), .B2(n_666), .C(n_681), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_682), .Y(n_701) );
AOI211xp5_ASAP7_75t_SL g702 ( .A1(n_687), .A2(n_676), .B(n_610), .C(n_612), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_692), .A2(n_610), .B(n_612), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_700), .A2(n_683), .B1(n_691), .B2(n_695), .Y(n_704) );
NOR2xp67_ASAP7_75t_SL g705 ( .A(n_701), .B(n_691), .Y(n_705) );
NAND5xp2_ASAP7_75t_L g706 ( .A(n_702), .B(n_690), .C(n_693), .D(n_688), .E(n_691), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_699), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_703), .B(n_443), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_707), .Y(n_709) );
NOR4xp25_ASAP7_75t_L g710 ( .A(n_704), .B(n_700), .C(n_697), .D(n_696), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_705), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_709), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_711), .Y(n_713) );
XNOR2xp5_ASAP7_75t_L g714 ( .A(n_713), .B(n_710), .Y(n_714) );
INVx4_ASAP7_75t_L g715 ( .A(n_712), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_715), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_714), .B(n_698), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_717), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_706), .B1(n_708), .B2(n_288), .Y(n_719) );
endmodule