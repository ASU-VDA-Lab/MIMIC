module real_jpeg_29674_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_0),
.B(n_70),
.Y(n_88)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_2),
.A2(n_21),
.B1(n_43),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_3),
.A2(n_7),
.B(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_3),
.A2(n_16),
.B1(n_28),
.B2(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_3),
.A2(n_16),
.B1(n_23),
.B2(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_3),
.A2(n_16),
.B1(n_21),
.B2(n_43),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_4),
.B(n_29),
.Y(n_80)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_5),
.A2(n_21),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_5),
.A2(n_23),
.B1(n_42),
.B2(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_72),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_71),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_61),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_13),
.B(n_61),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_35),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B(n_20),
.C(n_23),
.Y(n_15)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_16),
.A2(n_21),
.B(n_39),
.C(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_16),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_17),
.B(n_23),
.Y(n_58)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_18),
.A2(n_19),
.B1(n_21),
.B2(n_43),
.Y(n_54)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_21),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_23),
.A2(n_54),
.B(n_57),
.C(n_58),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B(n_33),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_27),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_27),
.B(n_33),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_28),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_31),
.B(n_33),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_31),
.B(n_91),
.Y(n_100)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_49),
.B1(n_50),
.B2(n_60),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_37),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.C(n_67),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_84),
.B(n_109),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_81),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_74),
.B(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_95),
.B(n_108),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_101),
.B(n_107),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);


endmodule