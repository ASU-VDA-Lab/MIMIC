module fake_jpeg_24932_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

HB1xp67_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_20),
.A2(n_23),
.B1(n_11),
.B2(n_15),
.Y(n_29)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_24),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_16),
.B1(n_15),
.B2(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_21),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_41),
.B1(n_42),
.B2(n_27),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_22),
.C(n_26),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_39),
.C(n_40),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_9),
.B(n_13),
.C(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_33),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_25),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_28),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_30),
.B(n_31),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_21),
.B1(n_14),
.B2(n_19),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_13),
.B(n_17),
.Y(n_43)
);

XNOR2x1_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_19),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_35),
.C(n_42),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_39),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.C(n_57),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_48),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_44),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_62),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_47),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_27),
.B1(n_33),
.B2(n_14),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_44),
.B1(n_19),
.B2(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_60),
.A3(n_63),
.B1(n_8),
.B2(n_3),
.C(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_66),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_63),
.B1(n_8),
.B2(n_4),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_69),
.C(n_68),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_71),
.Y(n_74)
);


endmodule