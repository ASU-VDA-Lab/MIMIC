module real_aes_18102_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1845;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1853;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_1779;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1802;
wire n_727;
wire n_397;
wire n_1056;
wire n_1855;
wire n_1083;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_1838;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_1851;
wire n_780;
wire n_931;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1868;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_394;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI211xp5_ASAP7_75t_L g1461 ( .A1(n_0), .A2(n_703), .B(n_1294), .C(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1473 ( .A(n_0), .Y(n_1473) );
INVx1_ASAP7_75t_L g563 ( .A(n_1), .Y(n_563) );
OAI211xp5_ASAP7_75t_L g626 ( .A1(n_1), .A2(n_627), .B(n_629), .C(n_638), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g1590 ( .A1(n_2), .A2(n_96), .B1(n_1557), .B2(n_1562), .Y(n_1590) );
INVx1_ASAP7_75t_L g358 ( .A(n_3), .Y(n_358) );
AND2x2_ASAP7_75t_L g405 ( .A(n_3), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g495 ( .A(n_3), .B(n_244), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_3), .B(n_368), .Y(n_715) );
INVx1_ASAP7_75t_L g1142 ( .A(n_4), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_5), .A2(n_143), .B1(n_681), .B2(n_1284), .Y(n_1283) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_5), .A2(n_143), .B1(n_699), .B2(n_709), .Y(n_1297) );
OAI22xp33_ASAP7_75t_L g1397 ( .A1(n_6), .A2(n_279), .B1(n_1072), .B2(n_1398), .Y(n_1397) );
OAI22xp33_ASAP7_75t_L g1404 ( .A1(n_6), .A2(n_279), .B1(n_1062), .B2(n_1063), .Y(n_1404) );
OAI22xp33_ASAP7_75t_L g1286 ( .A1(n_7), .A2(n_271), .B1(n_360), .B2(n_895), .Y(n_1286) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_7), .A2(n_271), .B1(n_698), .B2(n_1230), .Y(n_1292) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_8), .A2(n_72), .B1(n_605), .B2(n_606), .Y(n_1140) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_8), .A2(n_18), .B1(n_844), .B2(n_1169), .C(n_1171), .Y(n_1168) );
INVx1_ASAP7_75t_L g1336 ( .A(n_9), .Y(n_1336) );
INVx1_ASAP7_75t_L g379 ( .A(n_10), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_11), .A2(n_171), .B1(n_615), .B2(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g630 ( .A(n_11), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1853 ( .A1(n_12), .A2(n_24), .B1(n_534), .B2(n_1127), .Y(n_1853) );
INVx1_ASAP7_75t_L g1881 ( .A(n_12), .Y(n_1881) );
OAI211xp5_ASAP7_75t_L g800 ( .A1(n_13), .A2(n_703), .B(n_801), .C(n_805), .Y(n_800) );
INVx1_ASAP7_75t_L g814 ( .A(n_13), .Y(n_814) );
INVx1_ASAP7_75t_L g1200 ( .A(n_14), .Y(n_1200) );
INVx1_ASAP7_75t_L g1250 ( .A(n_15), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1778 ( .A1(n_16), .A2(n_338), .B1(n_1518), .B2(n_1520), .C(n_1779), .Y(n_1778) );
OAI21xp33_ASAP7_75t_SL g1816 ( .A1(n_16), .A2(n_1488), .B(n_1504), .Y(n_1816) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_17), .Y(n_1025) );
AOI22xp33_ASAP7_75t_SL g1157 ( .A1(n_18), .A2(n_227), .B1(n_1127), .B2(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g780 ( .A(n_19), .Y(n_780) );
INVx2_ASAP7_75t_L g391 ( .A(n_20), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_21), .A2(n_343), .B1(n_507), .B2(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g529 ( .A(n_21), .Y(n_529) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_22), .A2(n_283), .B1(n_360), .B2(n_691), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_22), .A2(n_283), .B1(n_1229), .B2(n_1230), .Y(n_1228) );
OAI22xp33_ASAP7_75t_L g1794 ( .A1(n_23), .A2(n_281), .B1(n_1795), .B2(n_1798), .Y(n_1794) );
INVx1_ASAP7_75t_L g1814 ( .A(n_23), .Y(n_1814) );
AOI221xp5_ASAP7_75t_L g1865 ( .A1(n_24), .A2(n_40), .B1(n_508), .B2(n_1866), .C(n_1868), .Y(n_1865) );
INVx1_ASAP7_75t_L g1421 ( .A(n_25), .Y(n_1421) );
INVx1_ASAP7_75t_L g1150 ( .A(n_26), .Y(n_1150) );
INVx1_ASAP7_75t_L g1349 ( .A(n_27), .Y(n_1349) );
OA222x2_ASAP7_75t_L g1480 ( .A1(n_28), .A2(n_81), .B1(n_238), .B2(n_1481), .C1(n_1484), .C2(n_1488), .Y(n_1480) );
INVx1_ASAP7_75t_L g1530 ( .A(n_28), .Y(n_1530) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_29), .Y(n_353) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_29), .B(n_351), .Y(n_1558) );
INVx1_ASAP7_75t_L g986 ( .A(n_30), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_31), .A2(n_318), .B1(n_636), .B2(n_637), .Y(n_1094) );
INVxp67_ASAP7_75t_SL g1111 ( .A(n_31), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_32), .A2(n_199), .B1(n_475), .B2(n_477), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_32), .A2(n_260), .B1(n_548), .B2(n_550), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g1854 ( .A1(n_33), .A2(n_207), .B1(n_867), .B2(n_1457), .Y(n_1854) );
INVx1_ASAP7_75t_L g1870 ( .A(n_33), .Y(n_1870) );
INVx1_ASAP7_75t_L g419 ( .A(n_34), .Y(n_419) );
INVx1_ASAP7_75t_L g1207 ( .A(n_35), .Y(n_1207) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_36), .Y(n_1033) );
XNOR2xp5_ASAP7_75t_L g767 ( .A(n_37), .B(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_37), .A2(n_75), .B1(n_1565), .B2(n_1574), .Y(n_1589) );
OAI22xp33_ASAP7_75t_L g1391 ( .A1(n_38), .A2(n_181), .B1(n_809), .B2(n_938), .Y(n_1391) );
OAI22xp33_ASAP7_75t_L g1405 ( .A1(n_38), .A2(n_181), .B1(n_360), .B2(n_691), .Y(n_1405) );
INVx1_ASAP7_75t_L g903 ( .A(n_39), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g1856 ( .A1(n_40), .A2(n_311), .B1(n_1127), .B2(n_1857), .Y(n_1856) );
INVxp67_ASAP7_75t_SL g1149 ( .A(n_41), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_41), .A2(n_170), .B1(n_964), .B2(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1342 ( .A(n_42), .Y(n_1342) );
INVx1_ASAP7_75t_L g912 ( .A(n_43), .Y(n_912) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_44), .A2(n_665), .B(n_668), .C(n_671), .Y(n_664) );
INVx1_ASAP7_75t_L g706 ( .A(n_44), .Y(n_706) );
INVx1_ASAP7_75t_L g1246 ( .A(n_45), .Y(n_1246) );
OAI211xp5_ASAP7_75t_L g1222 ( .A1(n_46), .A2(n_812), .B(n_889), .C(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1233 ( .A(n_46), .Y(n_1233) );
CKINVDCx5p33_ASAP7_75t_R g1501 ( .A(n_47), .Y(n_1501) );
INVx1_ASAP7_75t_L g1163 ( .A(n_48), .Y(n_1163) );
INVx1_ASAP7_75t_L g599 ( .A(n_49), .Y(n_599) );
AOI21xp33_ASAP7_75t_L g639 ( .A1(n_49), .A2(n_640), .B(n_641), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g1099 ( .A1(n_50), .A2(n_255), .B1(n_636), .B2(n_1100), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_50), .A2(n_232), .B1(n_1113), .B2(n_1114), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g1146 ( .A(n_51), .Y(n_1146) );
INVx1_ASAP7_75t_L g1189 ( .A(n_52), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_53), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g1855 ( .A1(n_54), .A2(n_69), .B1(n_1139), .B2(n_1153), .Y(n_1855) );
INVx1_ASAP7_75t_L g1869 ( .A(n_54), .Y(n_1869) );
INVx1_ASAP7_75t_L g727 ( .A(n_55), .Y(n_727) );
OAI22xp33_ASAP7_75t_SL g1088 ( .A1(n_56), .A2(n_241), .B1(n_737), .B2(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1128 ( .A(n_56), .Y(n_1128) );
INVx1_ASAP7_75t_L g583 ( .A(n_57), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_57), .A2(n_304), .B1(n_623), .B2(n_625), .Y(n_622) );
XNOR2xp5_ASAP7_75t_L g1331 ( .A(n_58), .B(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g990 ( .A(n_59), .Y(n_990) );
INVx1_ASAP7_75t_L g1302 ( .A(n_60), .Y(n_1302) );
AOI21xp33_ASAP7_75t_L g852 ( .A1(n_61), .A2(n_472), .B(n_853), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_61), .A2(n_262), .B1(n_867), .B2(n_875), .C(n_877), .Y(n_874) );
CKINVDCx5p33_ASAP7_75t_R g1849 ( .A(n_62), .Y(n_1849) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_63), .A2(n_113), .B1(n_1565), .B2(n_1574), .Y(n_1573) );
AOI22xp5_ASAP7_75t_L g1581 ( .A1(n_64), .A2(n_249), .B1(n_1565), .B2(n_1574), .Y(n_1581) );
INVx1_ASAP7_75t_L g1203 ( .A(n_65), .Y(n_1203) );
OAI222xp33_ASAP7_75t_L g829 ( .A1(n_66), .A2(n_79), .B1(n_86), .B2(n_381), .C1(n_830), .C2(n_831), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g1051 ( .A1(n_67), .A2(n_122), .B1(n_360), .B2(n_821), .Y(n_1051) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_67), .A2(n_122), .B1(n_698), .B2(n_809), .Y(n_1065) );
AOI21xp33_ASAP7_75t_L g502 ( .A1(n_68), .A2(n_503), .B(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_68), .A2(n_199), .B1(n_531), .B2(n_534), .Y(n_530) );
INVx1_ASAP7_75t_L g1885 ( .A(n_69), .Y(n_1885) );
INVx1_ASAP7_75t_L g1370 ( .A(n_70), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g1379 ( .A1(n_70), .A2(n_889), .B(n_1380), .C(n_1383), .Y(n_1379) );
INVx1_ASAP7_75t_L g1269 ( .A(n_71), .Y(n_1269) );
OAI211xp5_ASAP7_75t_L g1273 ( .A1(n_71), .A2(n_589), .B(n_872), .C(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1188 ( .A(n_72), .Y(n_1188) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_73), .A2(n_80), .B1(n_897), .B2(n_898), .Y(n_896) );
OAI22xp33_ASAP7_75t_L g945 ( .A1(n_73), .A2(n_80), .B1(n_709), .B2(n_946), .Y(n_945) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_74), .Y(n_836) );
AOI21xp33_ASAP7_75t_L g1800 ( .A1(n_76), .A2(n_1801), .B(n_1802), .Y(n_1800) );
AOI221xp5_ASAP7_75t_L g1829 ( .A1(n_76), .A2(n_110), .B1(n_1493), .B2(n_1830), .C(n_1831), .Y(n_1829) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_77), .Y(n_458) );
INVx1_ASAP7_75t_L g1245 ( .A(n_78), .Y(n_1245) );
OAI221xp5_ASAP7_75t_L g1517 ( .A1(n_81), .A2(n_191), .B1(n_1518), .B2(n_1520), .C(n_1522), .Y(n_1517) );
OAI22xp5_ASAP7_75t_L g1874 ( .A1(n_82), .A2(n_298), .B1(n_688), .B2(n_964), .Y(n_1874) );
INVx1_ASAP7_75t_L g1887 ( .A(n_82), .Y(n_1887) );
INVx1_ASAP7_75t_L g1495 ( .A(n_83), .Y(n_1495) );
AOI22xp33_ASAP7_75t_L g1544 ( .A1(n_83), .A2(n_131), .B1(n_546), .B2(n_548), .Y(n_1544) );
INVx1_ASAP7_75t_L g921 ( .A(n_84), .Y(n_921) );
XOR2x2_ASAP7_75t_L g952 ( .A(n_85), .B(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g1596 ( .A1(n_85), .A2(n_235), .B1(n_1565), .B2(n_1574), .Y(n_1596) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_86), .A2(n_340), .B1(n_625), .B2(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g1422 ( .A(n_87), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g1226 ( .A1(n_88), .A2(n_169), .B1(n_817), .B2(n_961), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g1234 ( .A1(n_88), .A2(n_169), .B1(n_1072), .B2(n_1235), .Y(n_1234) );
AOI22xp5_ASAP7_75t_L g1556 ( .A1(n_89), .A2(n_243), .B1(n_1557), .B2(n_1562), .Y(n_1556) );
XOR2x2_ASAP7_75t_L g1772 ( .A(n_89), .B(n_1773), .Y(n_1772) );
AOI22xp33_ASAP7_75t_L g1837 ( .A1(n_89), .A2(n_1838), .B1(n_1841), .B2(n_1888), .Y(n_1837) );
AOI22xp5_ASAP7_75t_L g1564 ( .A1(n_90), .A2(n_103), .B1(n_1565), .B2(n_1567), .Y(n_1564) );
AO22x1_ASAP7_75t_L g1587 ( .A1(n_91), .A2(n_251), .B1(n_1557), .B2(n_1562), .Y(n_1587) );
INVx1_ASAP7_75t_L g958 ( .A(n_92), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_93), .A2(n_159), .B1(n_477), .B2(n_507), .Y(n_854) );
INVx1_ASAP7_75t_L g869 ( .A(n_93), .Y(n_869) );
INVx1_ASAP7_75t_L g1340 ( .A(n_94), .Y(n_1340) );
XNOR2xp5_ASAP7_75t_L g1236 ( .A(n_95), .B(n_1237), .Y(n_1236) );
CKINVDCx5p33_ASAP7_75t_R g1162 ( .A(n_97), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_98), .A2(n_315), .B1(n_1153), .B2(n_1155), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_98), .A2(n_205), .B1(n_508), .B2(n_636), .C(n_1186), .Y(n_1185) );
OAI211xp5_ASAP7_75t_L g1287 ( .A1(n_99), .A2(n_665), .B(n_668), .C(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1296 ( .A(n_99), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1780 ( .A1(n_100), .A2(n_209), .B1(n_1781), .B2(n_1783), .Y(n_1780) );
INVxp67_ASAP7_75t_SL g1825 ( .A(n_100), .Y(n_1825) );
OAI22xp33_ASAP7_75t_L g1460 ( .A1(n_101), .A2(n_154), .B1(n_585), .B2(n_809), .Y(n_1460) );
OAI22xp33_ASAP7_75t_L g1467 ( .A1(n_101), .A2(n_154), .B1(n_360), .B2(n_691), .Y(n_1467) );
AOI222xp33_ASAP7_75t_L g1803 ( .A1(n_102), .A2(n_153), .B1(n_331), .B2(n_412), .C1(n_546), .C2(n_758), .Y(n_1803) );
INVx1_ASAP7_75t_L g1832 ( .A(n_102), .Y(n_1832) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_104), .A2(n_142), .B1(n_894), .B2(n_895), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_104), .A2(n_142), .B1(n_938), .B2(n_940), .Y(n_937) );
INVx1_ASAP7_75t_L g1224 ( .A(n_105), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_106), .A2(n_178), .B1(n_709), .B2(n_809), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_106), .A2(n_210), .B1(n_817), .B2(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g1440 ( .A(n_107), .Y(n_1440) );
INVx1_ASAP7_75t_L g613 ( .A(n_108), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_108), .A2(n_248), .B1(n_636), .B2(n_637), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_109), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g1786 ( .A1(n_110), .A2(n_220), .B1(n_1787), .B2(n_1788), .C(n_1789), .Y(n_1786) );
INVx1_ASAP7_75t_L g351 ( .A(n_111), .Y(n_351) );
INVx1_ASAP7_75t_L g1339 ( .A(n_112), .Y(n_1339) );
XOR2x2_ASAP7_75t_L g1388 ( .A(n_113), .B(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g776 ( .A(n_114), .Y(n_776) );
AO221x2_ASAP7_75t_L g1674 ( .A1(n_115), .A2(n_330), .B1(n_1557), .B2(n_1562), .C(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1777 ( .A(n_116), .Y(n_1777) );
OAI21xp33_ASAP7_75t_L g1810 ( .A1(n_116), .A2(n_1484), .B(n_1811), .Y(n_1810) );
OAI211xp5_ASAP7_75t_L g955 ( .A1(n_117), .A2(n_668), .B(n_956), .C(n_957), .Y(n_955) );
INVx1_ASAP7_75t_L g972 ( .A(n_117), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_118), .A2(n_341), .B1(n_681), .B2(n_685), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_118), .A2(n_126), .B1(n_698), .B2(n_699), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_119), .A2(n_152), .B1(n_817), .B2(n_961), .Y(n_1270) );
OAI22xp33_ASAP7_75t_L g1276 ( .A1(n_119), .A2(n_152), .B1(n_1235), .B2(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1290 ( .A(n_120), .Y(n_1290) );
OAI211xp5_ASAP7_75t_L g1293 ( .A1(n_120), .A2(n_589), .B(n_1294), .C(n_1295), .Y(n_1293) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_121), .A2(n_147), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1132 ( .A(n_121), .B(n_699), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g1862 ( .A(n_123), .Y(n_1862) );
INVx1_ASAP7_75t_L g1449 ( .A(n_124), .Y(n_1449) );
INVx1_ASAP7_75t_L g1204 ( .A(n_125), .Y(n_1204) );
OAI22xp33_ASAP7_75t_L g690 ( .A1(n_126), .A2(n_314), .B1(n_360), .B2(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g998 ( .A(n_127), .Y(n_998) );
INVx1_ASAP7_75t_L g1418 ( .A(n_128), .Y(n_1418) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_129), .A2(n_275), .B1(n_604), .B2(n_606), .Y(n_603) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_129), .A2(n_504), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g1268 ( .A(n_130), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_131), .A2(n_175), .B1(n_511), .B2(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1241 ( .A(n_132), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_133), .A2(n_325), .B1(n_817), .B2(n_961), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_133), .A2(n_325), .B1(n_699), .B2(n_967), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g1508 ( .A1(n_134), .A2(n_191), .B1(n_1509), .B2(n_1512), .Y(n_1508) );
INVx1_ASAP7_75t_L g1531 ( .A(n_134), .Y(n_1531) );
INVx1_ASAP7_75t_L g1442 ( .A(n_135), .Y(n_1442) );
INVx1_ASAP7_75t_L g1444 ( .A(n_136), .Y(n_1444) );
OAI211xp5_ASAP7_75t_L g1052 ( .A1(n_137), .A2(n_668), .B(n_1053), .C(n_1055), .Y(n_1052) );
INVx1_ASAP7_75t_L g1070 ( .A(n_137), .Y(n_1070) );
OAI22xp33_ASAP7_75t_L g962 ( .A1(n_138), .A2(n_183), .B1(n_821), .B2(n_963), .Y(n_962) );
OAI22xp33_ASAP7_75t_L g973 ( .A1(n_138), .A2(n_183), .B1(n_585), .B2(n_974), .Y(n_973) );
AO22x1_ASAP7_75t_L g1578 ( .A1(n_139), .A2(n_333), .B1(n_1557), .B2(n_1562), .Y(n_1578) );
INVx1_ASAP7_75t_L g915 ( .A(n_140), .Y(n_915) );
INVx1_ASAP7_75t_L g784 ( .A(n_141), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g1103 ( .A1(n_144), .A2(n_321), .B1(n_956), .B2(n_1104), .C(n_1105), .Y(n_1103) );
INVx1_ASAP7_75t_L g1123 ( .A(n_144), .Y(n_1123) );
INVx1_ASAP7_75t_L g1092 ( .A(n_145), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_145), .A2(n_255), .B1(n_1113), .B2(n_1119), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g1096 ( .A(n_146), .Y(n_1096) );
INVx1_ASAP7_75t_L g1126 ( .A(n_147), .Y(n_1126) );
INVx1_ASAP7_75t_L g1396 ( .A(n_148), .Y(n_1396) );
OAI211xp5_ASAP7_75t_L g1400 ( .A1(n_148), .A2(n_1382), .B(n_1401), .C(n_1402), .Y(n_1400) );
INVx1_ASAP7_75t_L g807 ( .A(n_149), .Y(n_807) );
OAI211xp5_ASAP7_75t_SL g811 ( .A1(n_149), .A2(n_668), .B(n_812), .C(n_813), .Y(n_811) );
OAI22xp33_ASAP7_75t_L g1371 ( .A1(n_150), .A2(n_252), .B1(n_698), .B2(n_974), .Y(n_1371) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_150), .A2(n_252), .B1(n_895), .B2(n_1375), .Y(n_1374) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_151), .A2(n_210), .B1(n_698), .B2(n_799), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g820 ( .A1(n_151), .A2(n_178), .B1(n_360), .B2(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g1822 ( .A(n_153), .Y(n_1822) );
INVx1_ASAP7_75t_L g1289 ( .A(n_155), .Y(n_1289) );
INVx1_ASAP7_75t_L g1416 ( .A(n_156), .Y(n_1416) );
INVx1_ASAP7_75t_L g1337 ( .A(n_157), .Y(n_1337) );
INVx1_ASAP7_75t_L g1346 ( .A(n_158), .Y(n_1346) );
INVxp67_ASAP7_75t_SL g878 ( .A(n_159), .Y(n_878) );
INVx1_ASAP7_75t_L g1463 ( .A(n_160), .Y(n_1463) );
OAI22xp33_ASAP7_75t_L g1364 ( .A1(n_161), .A2(n_188), .B1(n_709), .B2(n_1235), .Y(n_1364) );
OAI22xp33_ASAP7_75t_L g1376 ( .A1(n_161), .A2(n_188), .B1(n_681), .B2(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1210 ( .A(n_162), .Y(n_1210) );
INVx1_ASAP7_75t_L g1253 ( .A(n_163), .Y(n_1253) );
AO22x1_ASAP7_75t_L g1585 ( .A1(n_164), .A2(n_334), .B1(n_1565), .B2(n_1586), .Y(n_1585) );
CKINVDCx16_ASAP7_75t_R g1676 ( .A(n_165), .Y(n_1676) );
INVx1_ASAP7_75t_L g1419 ( .A(n_166), .Y(n_1419) );
INVx1_ASAP7_75t_L g1446 ( .A(n_167), .Y(n_1446) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_168), .A2(n_327), .B1(n_467), .B2(n_469), .C(n_472), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_168), .A2(n_343), .B1(n_544), .B2(n_545), .Y(n_543) );
INVxp67_ASAP7_75t_SL g1165 ( .A(n_170), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_171), .A2(n_275), .B1(n_636), .B2(n_637), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g1500 ( .A(n_172), .Y(n_1500) );
INVx1_ASAP7_75t_L g1078 ( .A(n_173), .Y(n_1078) );
INVx1_ASAP7_75t_L g721 ( .A(n_174), .Y(n_721) );
INVx1_ASAP7_75t_L g1540 ( .A(n_175), .Y(n_1540) );
XNOR2xp5_ASAP7_75t_L g1193 ( .A(n_176), .B(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g672 ( .A(n_177), .Y(n_672) );
INVx1_ASAP7_75t_L g989 ( .A(n_179), .Y(n_989) );
INVx1_ASAP7_75t_L g1252 ( .A(n_180), .Y(n_1252) );
INVx1_ASAP7_75t_L g959 ( .A(n_182), .Y(n_959) );
OAI211xp5_ASAP7_75t_L g968 ( .A1(n_182), .A2(n_703), .B(n_969), .C(n_971), .Y(n_968) );
INVx1_ASAP7_75t_L g1413 ( .A(n_184), .Y(n_1413) );
INVx1_ASAP7_75t_L g851 ( .A(n_185), .Y(n_851) );
AOI221x1_ASAP7_75t_SL g866 ( .A1(n_185), .A2(n_258), .B1(n_792), .B2(n_867), .C(n_868), .Y(n_866) );
AOI221x1_ASAP7_75t_SL g1490 ( .A1(n_186), .A2(n_253), .B1(n_1491), .B2(n_1493), .C(n_1494), .Y(n_1490) );
AOI21xp33_ASAP7_75t_L g1542 ( .A1(n_186), .A2(n_758), .B(n_1543), .Y(n_1542) );
AOI21xp33_ASAP7_75t_L g858 ( .A1(n_187), .A2(n_503), .B(n_504), .Y(n_858) );
INVx1_ASAP7_75t_L g879 ( .A(n_187), .Y(n_879) );
INVx2_ASAP7_75t_L g1560 ( .A(n_189), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_189), .B(n_1561), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_189), .B(n_295), .Y(n_1568) );
INVx1_ASAP7_75t_L g732 ( .A(n_190), .Y(n_732) );
INVx1_ASAP7_75t_L g738 ( .A(n_192), .Y(n_738) );
INVx1_ASAP7_75t_L g891 ( .A(n_193), .Y(n_891) );
INVx1_ASAP7_75t_L g1395 ( .A(n_194), .Y(n_1395) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_195), .A2(n_377), .B1(n_556), .B2(n_557), .Y(n_376) );
INVxp67_ASAP7_75t_L g557 ( .A(n_195), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g1496 ( .A(n_196), .Y(n_1496) );
INVx1_ASAP7_75t_L g747 ( .A(n_197), .Y(n_747) );
OAI211xp5_ASAP7_75t_L g888 ( .A1(n_198), .A2(n_778), .B(n_889), .C(n_890), .Y(n_888) );
INVx1_ASAP7_75t_L g944 ( .A(n_198), .Y(n_944) );
XOR2x2_ASAP7_75t_L g1279 ( .A(n_200), .B(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1464 ( .A(n_201), .Y(n_1464) );
OAI211xp5_ASAP7_75t_L g1468 ( .A1(n_201), .A2(n_846), .B(n_1469), .C(n_1472), .Y(n_1468) );
XOR2x2_ASAP7_75t_L g1009 ( .A(n_202), .B(n_1010), .Y(n_1009) );
INVx1_ASAP7_75t_L g1198 ( .A(n_203), .Y(n_1198) );
OAI221xp5_ASAP7_75t_SL g434 ( .A1(n_204), .A2(n_291), .B1(n_435), .B2(n_443), .C(n_451), .Y(n_434) );
INVx1_ASAP7_75t_L g489 ( .A(n_204), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_205), .A2(n_301), .B1(n_792), .B2(n_1139), .Y(n_1138) );
XNOR2xp5_ASAP7_75t_L g661 ( .A(n_206), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g1883 ( .A(n_207), .Y(n_1883) );
INVx2_ASAP7_75t_L g393 ( .A(n_208), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_208), .B(n_391), .Y(n_418) );
INVx1_ASAP7_75t_L g555 ( .A(n_208), .Y(n_555) );
INVxp67_ASAP7_75t_SL g1806 ( .A(n_209), .Y(n_1806) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_211), .A2(n_217), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
OAI22xp33_ASAP7_75t_L g1071 ( .A1(n_211), .A2(n_217), .B1(n_799), .B2(n_1072), .Y(n_1071) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_212), .Y(n_1023) );
INVx1_ASAP7_75t_L g806 ( .A(n_213), .Y(n_806) );
INVx1_ASAP7_75t_L g827 ( .A(n_214), .Y(n_827) );
INVx1_ASAP7_75t_L g750 ( .A(n_215), .Y(n_750) );
INVx1_ASAP7_75t_L g783 ( .A(n_216), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g1265 ( .A1(n_218), .A2(n_250), .B1(n_360), .B2(n_691), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_218), .A2(n_250), .B1(n_974), .B2(n_1229), .Y(n_1272) );
BUFx3_ASAP7_75t_L g385 ( .A(n_219), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g1818 ( .A(n_220), .B(n_1819), .Y(n_1818) );
INVx1_ASAP7_75t_L g1790 ( .A(n_221), .Y(n_1790) );
AOI22xp33_ASAP7_75t_L g1597 ( .A1(n_222), .A2(n_225), .B1(n_1557), .B2(n_1562), .Y(n_1597) );
INVx1_ASAP7_75t_L g399 ( .A(n_223), .Y(n_399) );
INVx1_ASAP7_75t_L g1206 ( .A(n_224), .Y(n_1206) );
OAI22xp5_ASAP7_75t_SL g839 ( .A1(n_226), .A2(n_276), .B1(n_454), .B2(n_460), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_226), .Y(n_849) );
INVx1_ASAP7_75t_L g1187 ( .A(n_227), .Y(n_1187) );
INVx1_ASAP7_75t_L g981 ( .A(n_228), .Y(n_981) );
INVx1_ASAP7_75t_L g1225 ( .A(n_229), .Y(n_1225) );
OAI211xp5_ASAP7_75t_SL g1231 ( .A1(n_229), .A2(n_703), .B(n_872), .C(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1411 ( .A(n_230), .Y(n_1411) );
CKINVDCx5p33_ASAP7_75t_R g1019 ( .A(n_231), .Y(n_1019) );
AOI21xp33_ASAP7_75t_L g1093 ( .A1(n_232), .A2(n_503), .B(n_504), .Y(n_1093) );
INVx1_ASAP7_75t_L g1305 ( .A(n_233), .Y(n_1305) );
INVx1_ASAP7_75t_L g911 ( .A(n_234), .Y(n_911) );
INVx1_ASAP7_75t_L g1415 ( .A(n_236), .Y(n_1415) );
INVx1_ASAP7_75t_L g781 ( .A(n_237), .Y(n_781) );
INVx1_ASAP7_75t_L g1523 ( .A(n_238), .Y(n_1523) );
INVx1_ASAP7_75t_L g576 ( .A(n_239), .Y(n_576) );
INVx1_ASAP7_75t_L g1348 ( .A(n_240), .Y(n_1348) );
INVx1_ASAP7_75t_L g1131 ( .A(n_241), .Y(n_1131) );
INVx1_ASAP7_75t_L g717 ( .A(n_242), .Y(n_717) );
BUFx3_ASAP7_75t_L g368 ( .A(n_244), .Y(n_368) );
INVx1_ASAP7_75t_L g406 ( .A(n_244), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g1678 ( .A(n_245), .Y(n_1678) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_246), .A2(n_265), .B1(n_1557), .B2(n_1562), .Y(n_1580) );
OAI22xp33_ASAP7_75t_L g1465 ( .A1(n_247), .A2(n_299), .B1(n_1277), .B2(n_1398), .Y(n_1465) );
OAI22xp5_ASAP7_75t_L g1474 ( .A1(n_247), .A2(n_299), .B1(n_817), .B2(n_961), .Y(n_1474) );
INVx1_ASAP7_75t_L g602 ( .A(n_248), .Y(n_602) );
INVx1_ASAP7_75t_L g1539 ( .A(n_253), .Y(n_1539) );
INVx1_ASAP7_75t_L g773 ( .A(n_254), .Y(n_773) );
INVx1_ASAP7_75t_L g1478 ( .A(n_256), .Y(n_1478) );
INVx1_ASAP7_75t_L g774 ( .A(n_257), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_258), .A2(n_262), .B1(n_477), .B2(n_507), .Y(n_859) );
INVx1_ASAP7_75t_L g1311 ( .A(n_259), .Y(n_1311) );
INVx1_ASAP7_75t_L g497 ( .A(n_260), .Y(n_497) );
INVx1_ASAP7_75t_L g892 ( .A(n_261), .Y(n_892) );
OAI211xp5_ASAP7_75t_L g941 ( .A1(n_261), .A2(n_589), .B(n_753), .C(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g1248 ( .A(n_263), .Y(n_1248) );
INVx1_ASAP7_75t_L g984 ( .A(n_264), .Y(n_984) );
INVx1_ASAP7_75t_L g1792 ( .A(n_266), .Y(n_1792) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_267), .Y(n_1027) );
INVx1_ASAP7_75t_L g916 ( .A(n_268), .Y(n_916) );
INVx1_ASAP7_75t_L g1310 ( .A(n_269), .Y(n_1310) );
INVx1_ASAP7_75t_L g1447 ( .A(n_270), .Y(n_1447) );
CKINVDCx5p33_ASAP7_75t_R g1863 ( .A(n_272), .Y(n_1863) );
AOI22xp5_ASAP7_75t_L g1572 ( .A1(n_273), .A2(n_337), .B1(n_1557), .B2(n_1562), .Y(n_1572) );
AO22x1_ASAP7_75t_L g1577 ( .A1(n_274), .A2(n_280), .B1(n_1565), .B2(n_1574), .Y(n_1577) );
INVx1_ASAP7_75t_L g843 ( .A(n_276), .Y(n_843) );
INVx1_ASAP7_75t_L g1307 ( .A(n_277), .Y(n_1307) );
INVx1_ASAP7_75t_L g388 ( .A(n_278), .Y(n_388) );
INVx1_ASAP7_75t_L g450 ( .A(n_278), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_280), .A2(n_559), .B1(n_560), .B2(n_659), .Y(n_558) );
INVxp67_ASAP7_75t_L g659 ( .A(n_280), .Y(n_659) );
INVxp67_ASAP7_75t_SL g1809 ( .A(n_281), .Y(n_1809) );
INVx1_ASAP7_75t_L g1314 ( .A(n_282), .Y(n_1314) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_284), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_285), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_285), .A2(n_328), .B1(n_645), .B2(n_646), .C(n_649), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g1266 ( .A1(n_286), .A2(n_812), .B(n_889), .C(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1275 ( .A(n_286), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_287), .Y(n_1021) );
INVx1_ASAP7_75t_L g856 ( .A(n_288), .Y(n_856) );
INVx1_ASAP7_75t_L g1450 ( .A(n_289), .Y(n_1450) );
INVx1_ASAP7_75t_L g1369 ( .A(n_290), .Y(n_1369) );
INVx1_ASAP7_75t_L g513 ( .A(n_291), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_292), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_293), .A2(n_885), .B1(n_886), .B2(n_947), .Y(n_884) );
INVxp67_ASAP7_75t_SL g947 ( .A(n_293), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g1859 ( .A(n_294), .Y(n_1859) );
INVx1_ASAP7_75t_L g1561 ( .A(n_295), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_295), .B(n_1560), .Y(n_1566) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_296), .Y(n_1032) );
OAI211xp5_ASAP7_75t_SL g1365 ( .A1(n_297), .A2(n_589), .B(n_1366), .C(n_1368), .Y(n_1365) );
INVx1_ASAP7_75t_L g1384 ( .A(n_297), .Y(n_1384) );
INVx1_ASAP7_75t_L g1850 ( .A(n_298), .Y(n_1850) );
INVx1_ASAP7_75t_L g979 ( .A(n_300), .Y(n_979) );
INVx1_ASAP7_75t_L g1173 ( .A(n_301), .Y(n_1173) );
INVx1_ASAP7_75t_L g740 ( .A(n_302), .Y(n_740) );
INVx1_ASAP7_75t_L g676 ( .A(n_303), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_303), .A2(n_701), .B(n_703), .C(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g586 ( .A(n_304), .Y(n_586) );
INVx1_ASAP7_75t_L g1102 ( .A(n_305), .Y(n_1102) );
INVx1_ASAP7_75t_L g1060 ( .A(n_306), .Y(n_1060) );
OAI211xp5_ASAP7_75t_L g1066 ( .A1(n_306), .A2(n_703), .B(n_1067), .C(n_1069), .Y(n_1066) );
INVx1_ASAP7_75t_L g1242 ( .A(n_307), .Y(n_1242) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_308), .Y(n_611) );
INVx1_ASAP7_75t_L g1313 ( .A(n_309), .Y(n_1313) );
INVx1_ASAP7_75t_L g777 ( .A(n_310), .Y(n_777) );
AOI211xp5_ASAP7_75t_SL g1878 ( .A1(n_311), .A2(n_1879), .B(n_1880), .C(n_1882), .Y(n_1878) );
AOI21xp5_ASAP7_75t_SL g1097 ( .A1(n_312), .A2(n_503), .B(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1110 ( .A(n_312), .Y(n_1110) );
INVx1_ASAP7_75t_L g1211 ( .A(n_313), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_314), .A2(n_341), .B1(n_708), .B2(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g1172 ( .A(n_315), .Y(n_1172) );
INVx1_ASAP7_75t_L g1437 ( .A(n_316), .Y(n_1437) );
XOR2x2_ASAP7_75t_L g1432 ( .A(n_317), .B(n_1433), .Y(n_1432) );
INVxp67_ASAP7_75t_L g1117 ( .A(n_318), .Y(n_1117) );
OAI211xp5_ASAP7_75t_L g1392 ( .A1(n_319), .A2(n_703), .B(n_1393), .C(n_1394), .Y(n_1392) );
INVx1_ASAP7_75t_L g1403 ( .A(n_319), .Y(n_1403) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_320), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1130 ( .A(n_321), .Y(n_1130) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_322), .Y(n_364) );
INVx1_ASAP7_75t_L g906 ( .A(n_323), .Y(n_906) );
INVx1_ASAP7_75t_L g922 ( .A(n_324), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_326), .Y(n_1514) );
INVx1_ASAP7_75t_L g524 ( .A(n_327), .Y(n_524) );
INVx1_ASAP7_75t_L g570 ( .A(n_328), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g1842 ( .A1(n_329), .A2(n_1843), .B1(n_1844), .B2(n_1845), .Y(n_1842) );
CKINVDCx5p33_ASAP7_75t_R g1843 ( .A(n_329), .Y(n_1843) );
AOI21xp33_ASAP7_75t_L g1823 ( .A1(n_331), .A2(n_982), .B(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g995 ( .A(n_332), .Y(n_995) );
INVx1_ASAP7_75t_L g1308 ( .A(n_335), .Y(n_1308) );
INVx1_ASAP7_75t_L g397 ( .A(n_336), .Y(n_397) );
INVx1_ASAP7_75t_L g439 ( .A(n_336), .Y(n_439) );
INVx2_ASAP7_75t_L g519 ( .A(n_336), .Y(n_519) );
INVx1_ASAP7_75t_L g1812 ( .A(n_338), .Y(n_1812) );
CKINVDCx5p33_ASAP7_75t_R g1515 ( .A(n_339), .Y(n_1515) );
INVx1_ASAP7_75t_L g838 ( .A(n_340), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g1851 ( .A(n_342), .Y(n_1851) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_369), .B(n_1548), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_354), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g1836 ( .A(n_348), .B(n_357), .Y(n_1836) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g1840 ( .A(n_350), .B(n_353), .Y(n_1840) );
INVx1_ASAP7_75t_L g1892 ( .A(n_350), .Y(n_1892) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g1894 ( .A(n_353), .B(n_1892), .Y(n_1894) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g694 ( .A(n_357), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g473 ( .A(n_358), .B(n_367), .Y(n_473) );
AND2x4_ASAP7_75t_L g505 ( .A(n_358), .B(n_368), .Y(n_505) );
INVx1_ASAP7_75t_L g894 ( .A(n_359), .Y(n_894) );
INVxp67_ASAP7_75t_SL g1375 ( .A(n_359), .Y(n_1375) );
AND2x4_ASAP7_75t_SL g1835 ( .A(n_359), .B(n_1836), .Y(n_1835) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_361), .B(n_366), .Y(n_360) );
OR2x6_ASAP7_75t_L g683 ( .A(n_361), .B(n_684), .Y(n_683) );
BUFx4f_ASAP7_75t_L g994 ( .A(n_361), .Y(n_994) );
INVx1_ASAP7_75t_L g1362 ( .A(n_361), .Y(n_1362) );
INVxp67_ASAP7_75t_L g1439 ( .A(n_361), .Y(n_1439) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx4f_ASAP7_75t_L g720 ( .A(n_362), .Y(n_720) );
INVx3_ASAP7_75t_L g964 ( .A(n_362), .Y(n_964) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx2_ASAP7_75t_L g408 ( .A(n_364), .Y(n_408) );
AND2x2_ASAP7_75t_L g431 ( .A(n_364), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g471 ( .A(n_364), .B(n_365), .Y(n_471) );
INVx2_ASAP7_75t_L g479 ( .A(n_364), .Y(n_479) );
NAND2x1_ASAP7_75t_L g501 ( .A(n_364), .B(n_365), .Y(n_501) );
INVx1_ASAP7_75t_L g653 ( .A(n_364), .Y(n_653) );
INVx1_ASAP7_75t_L g409 ( .A(n_365), .Y(n_409) );
INVx2_ASAP7_75t_L g432 ( .A(n_365), .Y(n_432) );
AND2x2_ASAP7_75t_L g478 ( .A(n_365), .B(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g488 ( .A(n_365), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_365), .B(n_479), .Y(n_689) );
OR2x2_ASAP7_75t_L g731 ( .A(n_365), .B(n_408), .Y(n_731) );
OR2x6_ASAP7_75t_L g963 ( .A(n_366), .B(n_964), .Y(n_963) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g670 ( .A(n_367), .Y(n_670) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx2_ASAP7_75t_L g675 ( .A(n_368), .Y(n_675) );
AND2x4_ASAP7_75t_L g679 ( .A(n_368), .B(n_652), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_1329), .B2(n_1547), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
XNOR2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_949), .Y(n_371) );
XOR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_825), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_660), .B2(n_824), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
XOR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_558), .Y(n_375) );
INVx1_ASAP7_75t_L g556 ( .A(n_377), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_398), .C(n_433), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_379), .A2(n_510), .B1(n_513), .B2(n_514), .Y(n_509) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx5_ASAP7_75t_L g1166 ( .A(n_381), .Y(n_1166) );
OR2x6_ASAP7_75t_L g381 ( .A(n_382), .B(n_394), .Y(n_381) );
INVx2_ASAP7_75t_L g1776 ( .A(n_382), .Y(n_1776) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_383), .B(n_389), .Y(n_382) );
BUFx3_ASAP7_75t_L g533 ( .A(n_383), .Y(n_533) );
INVx8_ASAP7_75t_L g549 ( .A(n_383), .Y(n_549) );
BUFx3_ASAP7_75t_L g605 ( .A(n_383), .Y(n_605) );
HB1xp67_ASAP7_75t_L g1528 ( .A(n_383), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_383), .B(n_1797), .Y(n_1796) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AND2x4_ASAP7_75t_L g425 ( .A(n_384), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g413 ( .A(n_385), .B(n_387), .Y(n_413) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_385), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_385), .B(n_450), .Y(n_457) );
AND2x4_ASAP7_75t_L g535 ( .A(n_385), .B(n_449), .Y(n_535) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g426 ( .A(n_388), .Y(n_426) );
AND2x4_ASAP7_75t_L g437 ( .A(n_389), .B(n_438), .Y(n_437) );
AND2x6_ASAP7_75t_L g1519 ( .A(n_389), .B(n_440), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_389), .B(n_447), .Y(n_1521) );
INVx1_ASAP7_75t_L g1525 ( .A(n_389), .Y(n_1525) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
NAND3x1_ASAP7_75t_L g553 ( .A(n_390), .B(n_554), .C(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g565 ( .A(n_390), .Y(n_565) );
OR2x6_ASAP7_75t_L g568 ( .A(n_390), .B(n_528), .Y(n_568) );
OR2x4_ASAP7_75t_L g585 ( .A(n_390), .B(n_413), .Y(n_585) );
AND2x4_ASAP7_75t_L g590 ( .A(n_390), .B(n_535), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g1007 ( .A(n_390), .B(n_555), .Y(n_1007) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp33_ASAP7_75t_SL g538 ( .A(n_391), .B(n_393), .Y(n_538) );
BUFx3_ASAP7_75t_L g574 ( .A(n_391), .Y(n_574) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_393), .Y(n_593) );
AND3x4_ASAP7_75t_L g882 ( .A(n_393), .B(n_574), .C(n_658), .Y(n_882) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_393), .B(n_574), .Y(n_1793) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g403 ( .A(n_395), .Y(n_403) );
INVx1_ASAP7_75t_L g695 ( .A(n_395), .Y(n_695) );
OR2x2_ASAP7_75t_L g1512 ( .A(n_395), .B(n_651), .Y(n_1512) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_419), .B2(n_420), .Y(n_398) );
INVxp67_ASAP7_75t_L g830 ( .A(n_400), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_410), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g1513 ( .A1(n_402), .A2(n_428), .B1(n_1514), .B2(n_1515), .Y(n_1513) );
AOI211xp5_ASAP7_75t_L g1808 ( .A1(n_402), .A2(n_1809), .B(n_1810), .C(n_1816), .Y(n_1808) );
AND2x4_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
AND2x4_ASAP7_75t_L g428 ( .A(n_403), .B(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_404), .Y(n_624) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
AND2x2_ASAP7_75t_L g429 ( .A(n_405), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g510 ( .A(n_405), .B(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_SL g515 ( .A(n_405), .B(n_470), .Y(n_515) );
AND2x4_ASAP7_75t_L g628 ( .A(n_405), .B(n_430), .Y(n_628) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_405), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_405), .B(n_439), .Y(n_1487) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_406), .Y(n_684) );
INVx3_ASAP7_75t_L g476 ( .A(n_407), .Y(n_476) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_407), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_407), .B(n_495), .Y(n_645) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_408), .Y(n_485) );
OR2x6_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_411), .A2(n_717), .B1(n_738), .B2(n_753), .Y(n_752) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_411), .A2(n_765), .B1(n_773), .B2(n_780), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_411), .A2(n_701), .B1(n_774), .B2(n_781), .Y(n_796) );
INVx2_ASAP7_75t_SL g905 ( .A(n_411), .Y(n_905) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g871 ( .A(n_412), .Y(n_871) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x4_ASAP7_75t_L g588 ( .A(n_413), .B(n_565), .Y(n_588) );
BUFx4f_ASAP7_75t_L g764 ( .A(n_413), .Y(n_764) );
BUFx3_ASAP7_75t_L g1018 ( .A(n_413), .Y(n_1018) );
BUFx3_ASAP7_75t_L g1199 ( .A(n_413), .Y(n_1199) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g422 ( .A(n_415), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g454 ( .A(n_416), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g460 ( .A(n_416), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g1144 ( .A(n_416), .Y(n_1144) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g537 ( .A(n_417), .B(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_417), .Y(n_595) );
INVx1_ASAP7_75t_L g745 ( .A(n_417), .Y(n_745) );
AND2x2_ASAP7_75t_SL g992 ( .A(n_417), .B(n_505), .Y(n_992) );
INVx1_ASAP7_75t_L g1534 ( .A(n_418), .Y(n_1534) );
INVx1_ASAP7_75t_L g1797 ( .A(n_418), .Y(n_1797) );
INVx1_ASAP7_75t_L g831 ( .A(n_420), .Y(n_831) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_421), .B(n_427), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g1116 ( .A(n_423), .Y(n_1116) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g544 ( .A(n_424), .Y(n_544) );
BUFx2_ASAP7_75t_L g610 ( .A(n_424), .Y(n_610) );
OR2x6_ASAP7_75t_SL g1781 ( .A(n_424), .B(n_1782), .Y(n_1781) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_425), .Y(n_523) );
BUFx8_ASAP7_75t_L g758 ( .A(n_425), .Y(n_758) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_425), .Y(n_789) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g1805 ( .A(n_428), .B(n_1806), .Y(n_1805) );
INVx1_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_430), .Y(n_503) );
INVx2_ASAP7_75t_L g1178 ( .A(n_430), .Y(n_1178) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g634 ( .A(n_431), .Y(n_634) );
AND2x4_ASAP7_75t_L g692 ( .A(n_431), .B(n_684), .Y(n_692) );
BUFx3_ASAP7_75t_L g853 ( .A(n_431), .Y(n_853) );
NOR3xp33_ASAP7_75t_SL g433 ( .A(n_434), .B(n_464), .C(n_520), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g1161 ( .A1(n_436), .A2(n_444), .B1(n_540), .B2(n_1162), .C(n_1163), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1861 ( .A1(n_436), .A2(n_444), .B1(n_540), .B2(n_1862), .C(n_1863), .Y(n_1861) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_437), .B(n_440), .Y(n_436) );
AND2x4_ASAP7_75t_SL g444 ( .A(n_437), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g540 ( .A(n_437), .B(n_541), .Y(n_540) );
NAND2x1_ASAP7_75t_L g835 ( .A(n_437), .B(n_440), .Y(n_835) );
AND2x4_ASAP7_75t_L g837 ( .A(n_437), .B(n_445), .Y(n_837) );
OR2x2_ASAP7_75t_L g1483 ( .A(n_438), .B(n_645), .Y(n_1483) );
INVx1_ASAP7_75t_L g1827 ( .A(n_438), .Y(n_1827) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g554 ( .A(n_439), .Y(n_554) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_442), .B(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g546 ( .A(n_442), .B(n_448), .Y(n_546) );
BUFx2_ASAP7_75t_L g575 ( .A(n_442), .Y(n_575) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g463 ( .A(n_450), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_458), .B2(n_459), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_452), .B(n_482), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g1145 ( .A1(n_453), .A2(n_459), .B1(n_1146), .B2(n_1147), .C1(n_1149), .C2(n_1150), .Y(n_1145) );
AOI222xp33_ASAP7_75t_L g1848 ( .A1(n_453), .A2(n_459), .B1(n_1147), .B2(n_1849), .C1(n_1850), .C2(n_1851), .Y(n_1848) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_456), .Y(n_601) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g528 ( .A(n_457), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_458), .A2(n_484), .B1(n_486), .B2(n_489), .C(n_490), .Y(n_483) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g702 ( .A(n_461), .Y(n_702) );
INVx4_ASAP7_75t_L g873 ( .A(n_461), .Y(n_873) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_461), .Y(n_909) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g755 ( .A(n_462), .Y(n_755) );
BUFx2_ASAP7_75t_L g804 ( .A(n_462), .Y(n_804) );
BUFx2_ASAP7_75t_L g579 ( .A(n_463), .Y(n_579) );
AOI31xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_496), .A3(n_509), .B(n_516), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_474), .B(n_480), .Y(n_465) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g1176 ( .A1(n_469), .A2(n_1142), .B1(n_1163), .B2(n_1177), .C(n_1179), .Y(n_1176) );
BUFx2_ASAP7_75t_L g1493 ( .A(n_469), .Y(n_1493) );
AOI221xp5_ASAP7_75t_L g1873 ( .A1(n_469), .A2(n_1177), .B1(n_1859), .B2(n_1863), .C(n_1874), .Y(n_1873) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x6_ASAP7_75t_L g654 ( .A(n_470), .B(n_495), .Y(n_654) );
AND2x2_ASAP7_75t_L g669 ( .A(n_470), .B(n_670), .Y(n_669) );
BUFx3_ASAP7_75t_L g1824 ( .A(n_470), .Y(n_1824) );
BUFx3_ASAP7_75t_L g1879 ( .A(n_470), .Y(n_1879) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g492 ( .A(n_471), .Y(n_492) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g641 ( .A(n_473), .Y(n_641) );
INVx1_ASAP7_75t_L g1098 ( .A(n_473), .Y(n_1098) );
OAI221xp5_ASAP7_75t_L g1171 ( .A1(n_473), .A2(n_857), .B1(n_932), .B2(n_1172), .C(n_1173), .Y(n_1171) );
OAI221xp5_ASAP7_75t_L g1868 ( .A1(n_473), .A2(n_857), .B1(n_1869), .B2(n_1870), .C(n_1871), .Y(n_1868) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g482 ( .A(n_476), .Y(n_482) );
INVx1_ASAP7_75t_L g507 ( .A(n_476), .Y(n_507) );
INVx2_ASAP7_75t_L g1503 ( .A(n_476), .Y(n_1503) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g508 ( .A(n_478), .Y(n_508) );
INVx2_ASAP7_75t_L g512 ( .A(n_478), .Y(n_512) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_478), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B(n_493), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_484), .A2(n_836), .B1(n_848), .B2(n_849), .Y(n_847) );
INVx1_ASAP7_75t_L g1105 ( .A(n_484), .Y(n_1105) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_484), .A2(n_848), .B1(n_1146), .B2(n_1162), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1877 ( .A1(n_484), .A2(n_488), .B1(n_1849), .B2(n_1862), .Y(n_1877) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g1104 ( .A(n_486), .Y(n_1104) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_487), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g674 ( .A(n_488), .B(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g848 ( .A(n_488), .Y(n_848) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_488), .B(n_675), .Y(n_1056) );
INVx1_ASAP7_75t_L g1511 ( .A(n_488), .Y(n_1511) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g1471 ( .A(n_492), .Y(n_1471) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g842 ( .A1(n_494), .A2(n_843), .B(n_844), .C(n_845), .Y(n_842) );
A2O1A1Ixp33_ASAP7_75t_SL g1101 ( .A1(n_494), .A2(n_844), .B(n_1102), .C(n_1103), .Y(n_1101) );
A2O1A1Ixp33_ASAP7_75t_L g1875 ( .A1(n_494), .A2(n_636), .B(n_1851), .C(n_1876), .Y(n_1875) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g648 ( .A(n_495), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_495), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g1507 ( .A(n_495), .B(n_519), .Y(n_1507) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_502), .C(n_506), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_498), .A2(n_735), .B1(n_780), .B2(n_781), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_498), .A2(n_1044), .B1(n_1203), .B2(n_1206), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_498), .A2(n_1044), .B1(n_1245), .B2(n_1248), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_498), .A2(n_932), .B1(n_1310), .B2(n_1311), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_498), .A2(n_1339), .B1(n_1342), .B2(n_1354), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g1356 ( .A1(n_498), .A2(n_1337), .B1(n_1349), .B2(n_1357), .Y(n_1356) );
OAI22xp5_ASAP7_75t_L g1445 ( .A1(n_498), .A2(n_1041), .B1(n_1446), .B2(n_1447), .Y(n_1445) );
INVx5_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
BUFx3_ASAP7_75t_L g631 ( .A(n_500), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_500), .B(n_1183), .Y(n_1182) );
BUFx2_ASAP7_75t_SL g1217 ( .A(n_500), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1488 ( .A(n_500), .B(n_1487), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1876 ( .A(n_500), .B(n_1877), .Y(n_1876) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_501), .Y(n_667) );
BUFx3_ASAP7_75t_L g1819 ( .A(n_503), .Y(n_1819) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_505), .B(n_744), .Y(n_743) );
AND2x4_ASAP7_75t_L g1047 ( .A(n_505), .B(n_744), .Y(n_1047) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_505), .A2(n_667), .B1(n_737), .B2(n_1187), .C(n_1188), .Y(n_1186) );
OAI21xp33_ASAP7_75t_L g1880 ( .A1(n_505), .A2(n_737), .B(n_1881), .Y(n_1880) );
INVx2_ASAP7_75t_L g625 ( .A(n_510), .Y(n_625) );
AND2x4_ASAP7_75t_L g1485 ( .A(n_511), .B(n_1486), .Y(n_1485) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g1100 ( .A(n_512), .Y(n_1100) );
AOI211xp5_ASAP7_75t_SL g643 ( .A1(n_514), .A2(n_576), .B(n_644), .C(n_654), .Y(n_643) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g863 ( .A(n_515), .Y(n_863) );
OAI31xp67_ASAP7_75t_L g1516 ( .A1(n_516), .A2(n_1517), .A3(n_1526), .B(n_1535), .Y(n_1516) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g714 ( .A(n_518), .B(n_715), .Y(n_714) );
OR2x6_ASAP7_75t_L g1006 ( .A(n_518), .B(n_1007), .Y(n_1006) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g658 ( .A(n_519), .Y(n_658) );
OAI211xp5_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_536), .B(n_539), .C(n_542), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_524), .B1(n_525), .B2(n_529), .C(n_530), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g564 ( .A(n_523), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g1022 ( .A(n_523), .Y(n_1022) );
BUFx6f_ASAP7_75t_L g1109 ( .A(n_523), .Y(n_1109) );
BUFx6f_ASAP7_75t_L g1457 ( .A(n_523), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_525), .A2(n_1021), .B1(n_1022), .B2(n_1023), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1426 ( .A1(n_525), .A2(n_1415), .B1(n_1421), .B2(n_1427), .Y(n_1426) );
OAI22xp5_ASAP7_75t_L g1428 ( .A1(n_525), .A2(n_793), .B1(n_1416), .B2(n_1422), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g1455 ( .A1(n_525), .A2(n_1444), .B1(n_1450), .B2(n_1456), .Y(n_1455) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g794 ( .A(n_527), .Y(n_794) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx3_ASAP7_75t_L g759 ( .A(n_528), .Y(n_759) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_534), .A2(n_867), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
BUFx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g541 ( .A(n_535), .Y(n_541) );
INVx2_ASAP7_75t_L g551 ( .A(n_535), .Y(n_551) );
BUFx2_ASAP7_75t_L g581 ( .A(n_535), .Y(n_581) );
BUFx2_ASAP7_75t_L g1119 ( .A(n_535), .Y(n_1119) );
BUFx3_ASAP7_75t_L g1124 ( .A(n_535), .Y(n_1124) );
BUFx2_ASAP7_75t_L g1158 ( .A(n_535), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1799 ( .A(n_535), .B(n_1797), .Y(n_1799) );
OAI33xp33_ASAP7_75t_L g751 ( .A1(n_536), .A2(n_619), .A3(n_752), .B1(n_756), .B2(n_760), .B3(n_762), .Y(n_751) );
OAI33xp33_ASAP7_75t_L g785 ( .A1(n_536), .A2(n_786), .A3(n_787), .B1(n_790), .B2(n_795), .B3(n_796), .Y(n_785) );
OAI33xp33_ASAP7_75t_L g1196 ( .A1(n_536), .A2(n_1028), .A3(n_1197), .B1(n_1202), .B2(n_1205), .B3(n_1209), .Y(n_1196) );
OAI33xp33_ASAP7_75t_L g1315 ( .A1(n_536), .A2(n_619), .A3(n_1316), .B1(n_1319), .B2(n_1320), .B3(n_1323), .Y(n_1315) );
OAI33xp33_ASAP7_75t_L g1334 ( .A1(n_536), .A2(n_619), .A3(n_1335), .B1(n_1338), .B2(n_1341), .B3(n_1347), .Y(n_1334) );
BUFx4f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx4f_ASAP7_75t_L g608 ( .A(n_537), .Y(n_608) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_537), .Y(n_1000) );
BUFx8_ASAP7_75t_L g1013 ( .A(n_537), .Y(n_1013) );
BUFx2_ASAP7_75t_L g1543 ( .A(n_538), .Y(n_1543) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_540), .A2(n_552), .B1(n_866), .B2(n_874), .C(n_881), .Y(n_865) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .C(n_552), .Y(n_542) );
INVx1_ASAP7_75t_L g598 ( .A(n_544), .Y(n_598) );
INVx1_ASAP7_75t_L g1249 ( .A(n_544), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_545), .A2(n_1102), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
BUFx12f_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx3_ASAP7_75t_L g867 ( .A(n_546), .Y(n_867) );
BUFx3_ASAP7_75t_L g1139 ( .A(n_546), .Y(n_1139) );
INVx5_ASAP7_75t_L g1156 ( .A(n_546), .Y(n_1156) );
AND2x4_ASAP7_75t_L g1784 ( .A(n_546), .B(n_1534), .Y(n_1784) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g1113 ( .A(n_549), .Y(n_1113) );
INVx8_ASAP7_75t_L g1127 ( .A(n_549), .Y(n_1127) );
INVx2_ASAP7_75t_L g1148 ( .A(n_549), .Y(n_1148) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g606 ( .A(n_551), .Y(n_606) );
INVx2_ASAP7_75t_L g1114 ( .A(n_551), .Y(n_1114) );
INVx1_ASAP7_75t_L g1857 ( .A(n_551), .Y(n_1857) );
INVx2_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
INVx2_ASAP7_75t_L g795 ( .A(n_552), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_552), .Y(n_1028) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx3_ASAP7_75t_L g919 ( .A(n_553), .Y(n_919) );
OAI33xp33_ASAP7_75t_L g1451 ( .A1(n_553), .A2(n_1013), .A3(n_1452), .B1(n_1454), .B2(n_1455), .B3(n_1458), .Y(n_1451) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI211xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_591), .B(n_596), .C(n_620), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g561 ( .A(n_562), .B(n_569), .C(n_582), .D(n_589), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B1(n_566), .B2(n_567), .Y(n_562) );
INVx1_ASAP7_75t_L g708 ( .A(n_564), .Y(n_708) );
INVx2_ASAP7_75t_L g809 ( .A(n_564), .Y(n_809) );
INVx2_ASAP7_75t_L g940 ( .A(n_564), .Y(n_940) );
INVx1_ASAP7_75t_L g974 ( .A(n_564), .Y(n_974) );
INVx1_ASAP7_75t_L g1230 ( .A(n_564), .Y(n_1230) );
INVx2_ASAP7_75t_L g967 ( .A(n_567), .Y(n_967) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx3_ASAP7_75t_L g709 ( .A(n_568), .Y(n_709) );
INVx1_ASAP7_75t_L g1073 ( .A(n_568), .Y(n_1073) );
INVx1_ASAP7_75t_L g1278 ( .A(n_568), .Y(n_1278) );
AOI222xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_576), .B2(n_577), .C1(n_580), .C2(n_581), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_571), .A2(n_577), .B1(n_1268), .B2(n_1275), .Y(n_1274) );
AOI22xp33_ASAP7_75t_SL g1394 ( .A1(n_571), .A2(n_578), .B1(n_1395), .B2(n_1396), .Y(n_1394) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g943 ( .A(n_572), .Y(n_943) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x4_ASAP7_75t_L g578 ( .A(n_573), .B(n_579), .Y(n_578) );
AND2x4_ASAP7_75t_L g705 ( .A(n_573), .B(n_575), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g1121 ( .A1(n_573), .A2(n_1122), .B(n_1125), .C(n_1129), .Y(n_1121) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_577), .A2(n_891), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1232 ( .A1(n_577), .A2(n_943), .B1(n_1224), .B2(n_1233), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_577), .A2(n_943), .B1(n_1289), .B2(n_1296), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_577), .A2(n_943), .B1(n_1369), .B2(n_1370), .Y(n_1368) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_578), .A2(n_672), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_578), .A2(n_705), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_578), .A2(n_705), .B1(n_958), .B2(n_972), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_578), .A2(n_705), .B1(n_1057), .B2(n_1070), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1129 ( .A1(n_578), .A2(n_705), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_578), .A2(n_705), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_580), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g618 ( .A(n_581), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B1(n_586), .B2(n_587), .Y(n_582) );
INVx2_ASAP7_75t_L g698 ( .A(n_584), .Y(n_698) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_SL g939 ( .A(n_585), .Y(n_939) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_585), .Y(n_1229) );
INVx2_ASAP7_75t_L g799 ( .A(n_587), .Y(n_799) );
INVx1_ASAP7_75t_L g946 ( .A(n_587), .Y(n_946) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g699 ( .A(n_588), .Y(n_699) );
BUFx2_ASAP7_75t_L g1235 ( .A(n_588), .Y(n_1235) );
BUFx3_ASAP7_75t_L g1398 ( .A(n_588), .Y(n_1398) );
CKINVDCx8_ASAP7_75t_R g589 ( .A(n_590), .Y(n_589) );
CKINVDCx8_ASAP7_75t_R g703 ( .A(n_590), .Y(n_703) );
OAI31xp33_ASAP7_75t_L g1120 ( .A1(n_590), .A2(n_1121), .A3(n_1132), .B(n_1133), .Y(n_1120) );
OAI31xp33_ASAP7_75t_L g797 ( .A1(n_591), .A2(n_798), .A3(n_800), .B(n_808), .Y(n_797) );
OAI31xp33_ASAP7_75t_L g1064 ( .A1(n_591), .A2(n_1065), .A3(n_1066), .B(n_1071), .Y(n_1064) );
CKINVDCx14_ASAP7_75t_R g1298 ( .A(n_591), .Y(n_1298) );
OAI31xp33_ASAP7_75t_L g1390 ( .A1(n_591), .A2(n_1391), .A3(n_1392), .B(n_1397), .Y(n_1390) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
AND2x2_ASAP7_75t_SL g710 ( .A(n_592), .B(n_594), .Y(n_710) );
AND2x2_ASAP7_75t_L g975 ( .A(n_592), .B(n_594), .Y(n_975) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_592), .B(n_594), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_592), .B(n_594), .Y(n_1372) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_607), .B1(n_609), .B2(n_619), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_600), .B2(n_602), .C(n_603), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_598), .A2(n_913), .B1(n_1307), .B2(n_1313), .Y(n_1319) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_600), .A2(n_1025), .B1(n_1026), .B2(n_1027), .Y(n_1024) );
OAI221xp5_ASAP7_75t_L g1107 ( .A1(n_600), .A2(n_1108), .B1(n_1110), .B2(n_1111), .C(n_1112), .Y(n_1107) );
OAI221xp5_ASAP7_75t_L g1115 ( .A1(n_600), .A2(n_1096), .B1(n_1116), .B2(n_1117), .C(n_1118), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_600), .A2(n_788), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1244 ( .A1(n_600), .A2(n_1026), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
OAI22xp5_ASAP7_75t_L g1454 ( .A1(n_600), .A2(n_1116), .B1(n_1442), .B2(n_1449), .Y(n_1454) );
OAI22xp5_ASAP7_75t_L g1538 ( .A1(n_600), .A2(n_1427), .B1(n_1539), .B2(n_1540), .Y(n_1538) );
CKINVDCx8_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
INVx3_ASAP7_75t_L g612 ( .A(n_601), .Y(n_612) );
INVx3_ASAP7_75t_L g913 ( .A(n_601), .Y(n_913) );
INVx1_ASAP7_75t_L g1003 ( .A(n_601), .Y(n_1003) );
INVx3_ASAP7_75t_L g1208 ( .A(n_601), .Y(n_1208) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g616 ( .A(n_605), .Y(n_616) );
INVx2_ASAP7_75t_SL g1791 ( .A(n_605), .Y(n_1791) );
OAI33xp33_ASAP7_75t_L g901 ( .A1(n_607), .A2(n_902), .A3(n_910), .B1(n_914), .B2(n_917), .B3(n_920), .Y(n_901) );
OAI22xp33_ASAP7_75t_L g1106 ( .A1(n_607), .A2(n_795), .B1(n_1107), .B2(n_1115), .Y(n_1106) );
BUFx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_612), .B2(n_613), .C(n_614), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_610), .A2(n_984), .B1(n_995), .B2(n_1003), .Y(n_1002) );
OAI211xp5_ASAP7_75t_SL g638 ( .A1(n_611), .A2(n_631), .B(n_639), .C(n_642), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_612), .A2(n_732), .B1(n_750), .B2(n_761), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_612), .A2(n_986), .B1(n_998), .B2(n_1005), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g1320 ( .A1(n_612), .A2(n_1308), .B1(n_1314), .B2(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_643), .B(n_655), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B(n_632), .C(n_635), .Y(n_629) );
BUFx2_ASAP7_75t_L g812 ( .A(n_631), .Y(n_812) );
INVx1_ASAP7_75t_L g1054 ( .A(n_631), .Y(n_1054) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g640 ( .A(n_634), .Y(n_640) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_636), .Y(n_844) );
A2O1A1Ixp33_ASAP7_75t_L g1181 ( .A1(n_636), .A2(n_1150), .B(n_1182), .C(n_1184), .Y(n_1181) );
INVx3_ASAP7_75t_L g1867 ( .A(n_636), .Y(n_1867) );
INVx1_ASAP7_75t_L g1170 ( .A(n_637), .Y(n_1170) );
INVx2_ASAP7_75t_L g1492 ( .A(n_640), .Y(n_1492) );
INVx1_ASAP7_75t_L g1828 ( .A(n_645), .Y(n_1828) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g1184 ( .A(n_648), .Y(n_1184) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_656), .Y(n_864) );
BUFx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g1081 ( .A(n_657), .Y(n_1081) );
OAI31xp33_ASAP7_75t_L g1167 ( .A1(n_657), .A2(n_1168), .A3(n_1174), .B(n_1185), .Y(n_1167) );
OAI31xp33_ASAP7_75t_L g1864 ( .A1(n_657), .A2(n_1865), .A3(n_1872), .B(n_1878), .Y(n_1864) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g1804 ( .A(n_658), .Y(n_1804) );
INVx1_ASAP7_75t_L g824 ( .A(n_660), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_766), .B1(n_767), .B2(n_823), .Y(n_660) );
INVx1_ASAP7_75t_L g823 ( .A(n_661), .Y(n_823) );
NAND3xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_696), .C(n_711), .Y(n_662) );
OAI31xp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_680), .A3(n_690), .B(n_693), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g850 ( .A1(n_665), .A2(n_851), .B(n_852), .C(n_854), .Y(n_850) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g739 ( .A(n_666), .Y(n_739) );
INVx1_ASAP7_75t_L g846 ( .A(n_666), .Y(n_846) );
INVx2_ASAP7_75t_L g857 ( .A(n_666), .Y(n_857) );
INVx4_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx4f_ASAP7_75t_L g733 ( .A(n_667), .Y(n_733) );
BUFx4f_ASAP7_75t_L g778 ( .A(n_667), .Y(n_778) );
BUFx6f_ASAP7_75t_L g956 ( .A(n_667), .Y(n_956) );
BUFx4f_ASAP7_75t_L g1089 ( .A(n_667), .Y(n_1089) );
BUFx4f_ASAP7_75t_L g1382 ( .A(n_667), .Y(n_1382) );
OR2x6_ASAP7_75t_L g1504 ( .A(n_667), .B(n_1505), .Y(n_1504) );
INVx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g889 ( .A(n_669), .Y(n_889) );
INVx1_ASAP7_75t_L g1401 ( .A(n_669), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_670), .B(n_1471), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_676), .B2(n_677), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_673), .A2(n_806), .B1(n_814), .B2(n_815), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_673), .A2(n_815), .B1(n_891), .B2(n_892), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_673), .A2(n_815), .B1(n_1289), .B2(n_1290), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_673), .A2(n_1058), .B1(n_1369), .B2(n_1384), .Y(n_1383) );
BUFx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_674), .A2(n_679), .B1(n_958), .B2(n_959), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_674), .A2(n_679), .B1(n_1268), .B2(n_1269), .Y(n_1267) );
OR2x2_ASAP7_75t_L g687 ( .A(n_675), .B(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_677), .A2(n_1056), .B1(n_1463), .B2(n_1473), .Y(n_1472) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx3_ASAP7_75t_L g815 ( .A(n_679), .Y(n_815) );
INVx2_ASAP7_75t_L g1059 ( .A(n_679), .Y(n_1059) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_683), .Y(n_817) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_683), .Y(n_897) );
BUFx2_ASAP7_75t_L g1062 ( .A(n_683), .Y(n_1062) );
INVx2_ASAP7_75t_L g1285 ( .A(n_685), .Y(n_1285) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g819 ( .A(n_687), .Y(n_819) );
INVx2_ASAP7_75t_L g899 ( .A(n_687), .Y(n_899) );
INVx8_ASAP7_75t_L g725 ( .A(n_688), .Y(n_725) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx4_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g821 ( .A(n_692), .Y(n_821) );
INVx3_ASAP7_75t_SL g895 ( .A(n_692), .Y(n_895) );
OAI31xp33_ASAP7_75t_L g1050 ( .A1(n_693), .A2(n_1051), .A3(n_1052), .B(n_1061), .Y(n_1050) );
OAI31xp33_ASAP7_75t_L g1220 ( .A1(n_693), .A2(n_1221), .A3(n_1222), .B(n_1226), .Y(n_1220) );
OAI31xp33_ASAP7_75t_L g1466 ( .A1(n_693), .A2(n_1467), .A3(n_1468), .B(n_1474), .Y(n_1466) );
BUFx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_SL g822 ( .A(n_694), .Y(n_822) );
OAI31xp33_ASAP7_75t_L g887 ( .A1(n_694), .A2(n_888), .A3(n_893), .B(n_896), .Y(n_887) );
INVx1_ASAP7_75t_L g1281 ( .A(n_694), .Y(n_1281) );
OAI31xp33_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_700), .A3(n_707), .B(n_710), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g1209 ( .A1(n_701), .A2(n_870), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g880 ( .A(n_702), .Y(n_880) );
OAI31xp33_ASAP7_75t_L g936 ( .A1(n_710), .A2(n_937), .A3(n_941), .B(n_945), .Y(n_936) );
OAI31xp33_ASAP7_75t_L g1227 ( .A1(n_710), .A2(n_1228), .A3(n_1231), .B(n_1234), .Y(n_1227) );
OAI31xp33_ASAP7_75t_L g1271 ( .A1(n_710), .A2(n_1272), .A3(n_1273), .B(n_1276), .Y(n_1271) );
NOR2xp33_ASAP7_75t_SL g711 ( .A(n_712), .B(n_751), .Y(n_711) );
OAI33xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_716), .A3(n_726), .B1(n_734), .B2(n_741), .B3(n_746), .Y(n_712) );
OAI33xp33_ASAP7_75t_L g923 ( .A1(n_713), .A2(n_741), .A3(n_924), .B1(n_931), .B2(n_934), .B3(n_935), .Y(n_923) );
INVx1_ASAP7_75t_L g1497 ( .A(n_713), .Y(n_1497) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx4_ASAP7_75t_L g771 ( .A(n_714), .Y(n_771) );
INVx2_ASAP7_75t_L g982 ( .A(n_714), .Y(n_982) );
INVx2_ASAP7_75t_L g1036 ( .A(n_714), .Y(n_1036) );
INVx1_ASAP7_75t_L g1351 ( .A(n_714), .Y(n_1351) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_721), .B2(n_722), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_718), .A2(n_747), .B1(n_748), .B2(n_750), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_718), .A2(n_722), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_718), .A2(n_748), .B1(n_783), .B2(n_784), .Y(n_782) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g1257 ( .A(n_719), .Y(n_1257) );
INVx2_ASAP7_75t_L g1263 ( .A(n_719), .Y(n_1263) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g927 ( .A(n_720), .Y(n_927) );
INVx4_ASAP7_75t_L g1884 ( .A(n_720), .Y(n_1884) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_721), .A2(n_740), .B1(n_763), .B2(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g1436 ( .A1(n_724), .A2(n_1437), .B1(n_1438), .B2(n_1440), .Y(n_1436) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g749 ( .A(n_725), .Y(n_749) );
INVx4_ASAP7_75t_L g930 ( .A(n_725), .Y(n_930) );
BUFx6f_ASAP7_75t_L g997 ( .A(n_725), .Y(n_997) );
INVx2_ASAP7_75t_L g1049 ( .A(n_725), .Y(n_1049) );
INVx2_ASAP7_75t_L g1087 ( .A(n_725), .Y(n_1087) );
INVx2_ASAP7_75t_L g1180 ( .A(n_725), .Y(n_1180) );
INVx1_ASAP7_75t_L g1258 ( .A(n_725), .Y(n_1258) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_732), .B2(n_733), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_727), .A2(n_747), .B1(n_757), .B2(n_759), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_728), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_775) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx4_ASAP7_75t_L g988 ( .A(n_729), .Y(n_988) );
INVx2_ASAP7_75t_L g1261 ( .A(n_729), .Y(n_1261) );
INVx2_ASAP7_75t_L g1443 ( .A(n_729), .Y(n_1443) );
INVx4_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
BUFx3_ASAP7_75t_L g737 ( .A(n_731), .Y(n_737) );
INVx2_ASAP7_75t_L g933 ( .A(n_731), .Y(n_933) );
BUFx2_ASAP7_75t_L g985 ( .A(n_731), .Y(n_985) );
INVx1_ASAP7_75t_L g1042 ( .A(n_731), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_733), .A2(n_911), .B1(n_915), .B2(n_932), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_733), .A2(n_906), .B1(n_922), .B2(n_932), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g1306 ( .A1(n_733), .A2(n_932), .B1(n_1307), .B2(n_1308), .Y(n_1306) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1414 ( .A1(n_735), .A2(n_1382), .B1(n_1415), .B2(n_1416), .Y(n_1414) );
INVx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_737), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_739), .A2(n_988), .B1(n_989), .B2(n_990), .Y(n_987) );
OAI33xp33_ASAP7_75t_L g1300 ( .A1(n_741), .A2(n_982), .A3(n_1301), .B1(n_1306), .B2(n_1309), .B3(n_1312), .Y(n_1300) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI33xp33_ASAP7_75t_L g770 ( .A1(n_743), .A2(n_771), .A3(n_772), .B1(n_775), .B2(n_779), .B3(n_782), .Y(n_770) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_748), .A2(n_1340), .B1(n_1346), .B2(n_1359), .Y(n_1358) );
BUFx3_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_753), .A2(n_904), .B1(n_921), .B2(n_922), .Y(n_920) );
OAI22xp33_ASAP7_75t_L g1014 ( .A1(n_753), .A2(n_1015), .B1(n_1016), .B2(n_1019), .Y(n_1014) );
OAI22xp33_ASAP7_75t_L g1316 ( .A1(n_753), .A2(n_1302), .B1(n_1310), .B2(n_1317), .Y(n_1316) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_755), .Y(n_765) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_755), .A2(n_871), .B1(n_981), .B2(n_990), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g1243 ( .A(n_755), .Y(n_1243) );
HB1xp67_ASAP7_75t_L g1254 ( .A(n_755), .Y(n_1254) );
INVx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx3_ASAP7_75t_L g761 ( .A(n_758), .Y(n_761) );
INVx2_ASAP7_75t_SL g876 ( .A(n_758), .Y(n_876) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_758), .Y(n_1005) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_758), .B(n_1144), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_759), .A2(n_776), .B1(n_783), .B2(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g1247 ( .A1(n_759), .A2(n_1248), .B1(n_1249), .B2(n_1250), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_759), .A2(n_791), .B1(n_1339), .B2(n_1340), .Y(n_1338) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_761), .A2(n_913), .B1(n_915), .B2(n_916), .Y(n_914) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_764), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_877) );
INVx1_ASAP7_75t_L g1318 ( .A(n_764), .Y(n_1318) );
OAI22xp33_ASAP7_75t_L g1323 ( .A1(n_765), .A2(n_1305), .B1(n_1311), .B2(n_1324), .Y(n_1323) );
OAI22xp33_ASAP7_75t_L g1335 ( .A1(n_765), .A2(n_1030), .B1(n_1336), .B2(n_1337), .Y(n_1335) );
OAI22xp33_ASAP7_75t_L g1347 ( .A1(n_765), .A2(n_1030), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_797), .C(n_810), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_785), .Y(n_769) );
INVx2_ASAP7_75t_SL g1409 ( .A(n_771), .Y(n_1409) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_777), .A2(n_784), .B1(n_791), .B2(n_794), .Y(n_790) );
INVx2_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
INVx5_ASAP7_75t_L g793 ( .A(n_789), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_789), .A2(n_1126), .B1(n_1127), .B2(n_1128), .Y(n_1125) );
INVx2_ASAP7_75t_SL g1154 ( .A(n_789), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_789), .Y(n_1322) );
INVx3_ASAP7_75t_L g1345 ( .A(n_789), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_791), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx8_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
BUFx3_ASAP7_75t_L g1026 ( .A(n_793), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g1029 ( .A1(n_802), .A2(n_1030), .B1(n_1032), .B2(n_1033), .Y(n_1029) );
INVxp67_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g1453 ( .A(n_803), .Y(n_1453) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g1367 ( .A(n_804), .Y(n_1367) );
OR2x6_ASAP7_75t_L g1779 ( .A(n_804), .B(n_1525), .Y(n_1779) );
OAI31xp33_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_816), .A3(n_820), .B(n_822), .Y(n_810) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_SL g1378 ( .A(n_819), .Y(n_1378) );
OAI31xp33_ASAP7_75t_L g954 ( .A1(n_822), .A2(n_955), .A3(n_960), .B(n_962), .Y(n_954) );
OAI31xp33_ASAP7_75t_L g1264 ( .A1(n_822), .A2(n_1265), .A3(n_1266), .B(n_1270), .Y(n_1264) );
OAI31xp33_ASAP7_75t_SL g1373 ( .A1(n_822), .A2(n_1374), .A3(n_1376), .B(n_1379), .Y(n_1373) );
OAI31xp33_ASAP7_75t_L g1399 ( .A1(n_822), .A2(n_1400), .A3(n_1404), .B(n_1405), .Y(n_1399) );
AO22x2_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_883), .B1(n_884), .B2(n_948), .Y(n_825) );
INVx1_ASAP7_75t_SL g948 ( .A(n_826), .Y(n_948) );
XNOR2x1_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
NOR2x1_ASAP7_75t_L g828 ( .A(n_829), .B(n_832), .Y(n_828) );
NAND3xp33_ASAP7_75t_SL g832 ( .A(n_833), .B(n_840), .C(n_865), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_836), .B1(n_837), .B2(n_838), .C(n_839), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_860), .B(n_864), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_850), .C(n_855), .Y(n_841) );
NAND2xp5_ASAP7_75t_SL g845 ( .A(n_846), .B(n_847), .Y(n_845) );
OAI22xp5_ASAP7_75t_SL g983 ( .A1(n_846), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
BUFx2_ASAP7_75t_L g1830 ( .A(n_853), .Y(n_1830) );
OAI211xp5_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .B(n_858), .C(n_859), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_856), .A2(n_869), .B1(n_870), .B2(n_872), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_857), .A2(n_1019), .B1(n_1033), .B2(n_1044), .Y(n_1043) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx4_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
BUFx4f_ASAP7_75t_SL g870 ( .A(n_871), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g1001 ( .A1(n_871), .A2(n_880), .B1(n_979), .B2(n_989), .Y(n_1001) );
OAI22xp33_ASAP7_75t_L g1431 ( .A1(n_872), .A2(n_1030), .B1(n_1413), .B2(n_1419), .Y(n_1431) );
INVx1_ASAP7_75t_L g1788 ( .A(n_872), .Y(n_1788) );
INVx2_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx2_ASAP7_75t_L g970 ( .A(n_873), .Y(n_970) );
INVx1_ASAP7_75t_L g1068 ( .A(n_873), .Y(n_1068) );
INVx1_ASAP7_75t_L g1294 ( .A(n_873), .Y(n_1294) );
INVx1_ASAP7_75t_L g1425 ( .A(n_873), .Y(n_1425) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_880), .Y(n_1393) );
OAI211xp5_ASAP7_75t_L g1541 ( .A1(n_880), .A2(n_1500), .B(n_1542), .C(n_1544), .Y(n_1541) );
BUFx3_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g1137 ( .A(n_882), .B(n_1138), .C(n_1140), .Y(n_1137) );
AOI33xp33_ASAP7_75t_L g1852 ( .A1(n_882), .A2(n_1159), .A3(n_1853), .B1(n_1854), .B2(n_1855), .B3(n_1856), .Y(n_1852) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NAND3xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_900), .C(n_936), .Y(n_886) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g961 ( .A(n_899), .Y(n_961) );
INVx1_ASAP7_75t_L g1063 ( .A(n_899), .Y(n_1063) );
NOR2xp33_ASAP7_75t_SL g900 ( .A(n_901), .B(n_923), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B1(n_906), .B2(n_907), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_903), .A2(n_921), .B1(n_925), .B2(n_928), .Y(n_924) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g1324 ( .A(n_905), .Y(n_1324) );
INVx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
HB1xp67_ASAP7_75t_L g1201 ( .A(n_909), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_912), .A2(n_916), .B1(n_925), .B2(n_928), .Y(n_935) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
BUFx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
BUFx2_ASAP7_75t_L g1430 ( .A(n_919), .Y(n_1430) );
OAI22xp5_ASAP7_75t_L g1213 ( .A1(n_925), .A2(n_1198), .B1(n_1210), .B2(n_1214), .Y(n_1213) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx2_ASAP7_75t_SL g926 ( .A(n_927), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_927), .A2(n_1204), .B1(n_1207), .B2(n_1214), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1301 ( .A1(n_928), .A2(n_1302), .B1(n_1303), .B2(n_1305), .Y(n_1301) );
OAI22xp5_ASAP7_75t_L g1312 ( .A1(n_928), .A2(n_1303), .B1(n_1313), .B2(n_1314), .Y(n_1312) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g978 ( .A1(n_930), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1882 ( .A1(n_930), .A2(n_1883), .B1(n_1884), .B2(n_1885), .Y(n_1882) );
INVx1_ASAP7_75t_L g1355 ( .A(n_932), .Y(n_1355) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_933), .Y(n_1045) );
INVx2_ASAP7_75t_L g1871 ( .A(n_933), .Y(n_1871) );
INVx2_ASAP7_75t_SL g938 ( .A(n_939), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_1191), .B1(n_1327), .B2(n_1328), .Y(n_949) );
INVx1_ASAP7_75t_L g1327 ( .A(n_950), .Y(n_1327) );
AOI22xp5_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_1074), .B1(n_1075), .B2(n_1190), .Y(n_950) );
INVx1_ASAP7_75t_L g1190 ( .A(n_951), .Y(n_1190) );
XNOR2xp5_ASAP7_75t_L g951 ( .A(n_952), .B(n_1009), .Y(n_951) );
NAND3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_965), .C(n_976), .Y(n_953) );
OAI22xp5_ASAP7_75t_SL g1040 ( .A1(n_956), .A2(n_1021), .B1(n_1025), .B2(n_1041), .Y(n_1040) );
BUFx6f_ASAP7_75t_L g980 ( .A(n_964), .Y(n_980) );
INVx2_ASAP7_75t_SL g1039 ( .A(n_964), .Y(n_1039) );
BUFx3_ASAP7_75t_L g1085 ( .A(n_964), .Y(n_1085) );
BUFx3_ASAP7_75t_L g1412 ( .A(n_964), .Y(n_1412) );
OAI31xp33_ASAP7_75t_L g965 ( .A1(n_966), .A2(n_968), .A3(n_973), .B(n_975), .Y(n_965) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g1536 ( .A1(n_970), .A2(n_1199), .B1(n_1496), .B2(n_1501), .C(n_1537), .Y(n_1536) );
NOR2xp33_ASAP7_75t_SL g976 ( .A(n_977), .B(n_999), .Y(n_976) );
OAI33xp33_ASAP7_75t_L g977 ( .A1(n_978), .A2(n_982), .A3(n_983), .B1(n_987), .B2(n_991), .B3(n_993), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_988), .A2(n_1089), .B1(n_1418), .B2(n_1419), .Y(n_1417) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_995), .B1(n_996), .B2(n_998), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_994), .A2(n_996), .B1(n_1421), .B2(n_1422), .Y(n_1420) );
OAI22xp5_ASAP7_75t_L g1821 ( .A1(n_994), .A2(n_996), .B1(n_1792), .B2(n_1822), .Y(n_1821) );
OAI22xp33_ASAP7_75t_L g1037 ( .A1(n_996), .A2(n_1015), .B1(n_1032), .B2(n_1038), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_996), .A2(n_1038), .B1(n_1449), .B2(n_1450), .Y(n_1448) );
INVx5_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx6_ASAP7_75t_L g1214 ( .A(n_997), .Y(n_1214) );
OAI33xp33_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1001), .A3(n_1002), .B1(n_1004), .B2(n_1006), .B3(n_1008), .Y(n_999) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1006), .Y(n_1159) );
INVx3_ASAP7_75t_L g1537 ( .A(n_1007), .Y(n_1537) );
NAND3xp33_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1050), .C(n_1064), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1034), .Y(n_1011) );
OAI33xp33_ASAP7_75t_L g1012 ( .A1(n_1013), .A2(n_1014), .A3(n_1020), .B1(n_1024), .B2(n_1028), .B3(n_1029), .Y(n_1012) );
OAI33xp33_ASAP7_75t_L g1239 ( .A1(n_1013), .A2(n_1028), .A3(n_1240), .B1(n_1244), .B2(n_1247), .B3(n_1251), .Y(n_1239) );
OAI33xp33_ASAP7_75t_L g1423 ( .A1(n_1013), .A2(n_1424), .A3(n_1426), .B1(n_1428), .B2(n_1429), .B3(n_1431), .Y(n_1423) );
OAI22xp33_ASAP7_75t_L g1452 ( .A1(n_1016), .A2(n_1437), .B1(n_1446), .B2(n_1453), .Y(n_1452) );
OAI22xp33_ASAP7_75t_L g1458 ( .A1(n_1016), .A2(n_1294), .B1(n_1440), .B2(n_1447), .Y(n_1458) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1018), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_1022), .A2(n_1206), .B1(n_1207), .B2(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1022), .Y(n_1787) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_1023), .A2(n_1027), .B1(n_1038), .B2(n_1049), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1424 ( .A1(n_1030), .A2(n_1411), .B1(n_1418), .B2(n_1425), .Y(n_1424) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
OAI33xp33_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1037), .A3(n_1040), .B1(n_1043), .B2(n_1046), .B3(n_1048), .Y(n_1034) );
OAI33xp33_ASAP7_75t_L g1212 ( .A1(n_1035), .A2(n_1213), .A3(n_1215), .B1(n_1216), .B2(n_1218), .B3(n_1219), .Y(n_1212) );
OAI33xp33_ASAP7_75t_L g1255 ( .A1(n_1035), .A2(n_1218), .A3(n_1256), .B1(n_1259), .B2(n_1260), .B3(n_1262), .Y(n_1255) );
OAI33xp33_ASAP7_75t_L g1435 ( .A1(n_1035), .A2(n_1046), .A3(n_1436), .B1(n_1441), .B2(n_1445), .B3(n_1448), .Y(n_1435) );
BUFx6f_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
OAI221xp5_ASAP7_75t_L g1499 ( .A1(n_1041), .A2(n_1089), .B1(n_1500), .B2(n_1501), .C(n_1502), .Y(n_1499) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_1044), .A2(n_1200), .B1(n_1211), .B2(n_1217), .Y(n_1216) );
INVx4_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
OAI33xp33_ASAP7_75t_L g1407 ( .A1(n_1046), .A2(n_1408), .A3(n_1410), .B1(n_1414), .B2(n_1417), .B3(n_1420), .Y(n_1407) );
OAI21xp5_ASAP7_75t_L g1498 ( .A1(n_1046), .A2(n_1499), .B(n_1504), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_1047), .Y(n_1046) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1047), .Y(n_1218) );
AOI322xp5_ASAP7_75t_L g1817 ( .A1(n_1047), .A2(n_1818), .A3(n_1820), .B1(n_1823), .B2(n_1825), .C1(n_1826), .C2(n_1829), .Y(n_1817) );
OAI22xp33_ASAP7_75t_L g1410 ( .A1(n_1049), .A2(n_1411), .B1(n_1412), .B2(n_1413), .Y(n_1410) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_1056), .A2(n_1057), .B1(n_1058), .B2(n_1060), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_1056), .A2(n_1058), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_1056), .A2(n_1058), .B1(n_1395), .B2(n_1403), .Y(n_1402) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
XOR2xp5_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1134), .Y(n_1076) );
XNOR2x1_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1079), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1120), .Y(n_1079) );
AOI21xp5_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B(n_1106), .Y(n_1080) );
NAND4xp25_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1091), .C(n_1095), .D(n_1101), .Y(n_1082) );
OAI21xp5_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1088), .B(n_1090), .Y(n_1083) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1085), .Y(n_1304) );
OAI22xp5_ASAP7_75t_L g1494 ( .A1(n_1085), .A2(n_1086), .B1(n_1495), .B2(n_1496), .Y(n_1494) );
BUFx6f_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
OAI211xp5_ASAP7_75t_SL g1091 ( .A1(n_1089), .A2(n_1092), .B(n_1093), .C(n_1094), .Y(n_1091) );
OAI211xp5_ASAP7_75t_SL g1095 ( .A1(n_1089), .A2(n_1096), .B(n_1097), .C(n_1099), .Y(n_1095) );
INVxp67_ASAP7_75t_L g1175 ( .A(n_1090), .Y(n_1175) );
INVx2_ASAP7_75t_SL g1108 ( .A(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1109), .Y(n_1427) );
A2O1A1Ixp33_ASAP7_75t_L g1522 ( .A1(n_1113), .A2(n_1124), .B(n_1523), .C(n_1524), .Y(n_1522) );
XNOR2x1_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1189), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1160), .Y(n_1135) );
NAND4xp25_ASAP7_75t_SL g1136 ( .A(n_1137), .B(n_1141), .C(n_1145), .D(n_1151), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1858 ( .A(n_1143), .B(n_1859), .Y(n_1858) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_1144), .B(n_1148), .Y(n_1147) );
NAND3xp33_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1157), .C(n_1159), .Y(n_1151) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
OAI221xp5_ASAP7_75t_L g1789 ( .A1(n_1156), .A2(n_1790), .B1(n_1791), .B2(n_1792), .C(n_1793), .Y(n_1789) );
NAND3xp33_ASAP7_75t_SL g1160 ( .A(n_1161), .B(n_1164), .C(n_1167), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1166), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1886 ( .A(n_1166), .B(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
OAI21xp5_ASAP7_75t_SL g1174 ( .A1(n_1175), .A2(n_1176), .B(n_1181), .Y(n_1174) );
OAI21xp33_ASAP7_75t_L g1872 ( .A1(n_1175), .A2(n_1873), .B(n_1875), .Y(n_1872) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
OAI22xp5_ASAP7_75t_L g1831 ( .A1(n_1180), .A2(n_1412), .B1(n_1790), .B2(n_1832), .Y(n_1831) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1191), .Y(n_1328) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_1192), .A2(n_1279), .B1(n_1325), .B2(n_1326), .Y(n_1191) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1192), .Y(n_1325) );
XOR2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1236), .Y(n_1192) );
AND3x1_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1220), .C(n_1227), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1212), .Y(n_1195) );
OAI22xp33_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1199), .B1(n_1200), .B2(n_1201), .Y(n_1197) );
OAI22xp33_ASAP7_75t_L g1240 ( .A1(n_1199), .A2(n_1241), .B1(n_1242), .B2(n_1243), .Y(n_1240) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_1199), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_1208), .A2(n_1342), .B1(n_1343), .B2(n_1346), .Y(n_1341) );
OAI22xp5_ASAP7_75t_L g1262 ( .A1(n_1214), .A2(n_1246), .B1(n_1250), .B2(n_1263), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1352 ( .A1(n_1214), .A2(n_1263), .B1(n_1336), .B2(n_1348), .Y(n_1352) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_1217), .A2(n_1242), .B1(n_1253), .B2(n_1261), .Y(n_1260) );
OAI33xp33_ASAP7_75t_L g1350 ( .A1(n_1218), .A2(n_1351), .A3(n_1352), .B1(n_1353), .B2(n_1356), .B3(n_1358), .Y(n_1350) );
AND3x1_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1264), .C(n_1271), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1255), .Y(n_1238) );
OAI22xp33_ASAP7_75t_L g1256 ( .A1(n_1241), .A2(n_1252), .B1(n_1257), .B2(n_1258), .Y(n_1256) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1279), .Y(n_1326) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1282), .B1(n_1291), .B2(n_1298), .C(n_1299), .Y(n_1280) );
NOR3xp33_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1286), .C(n_1287), .Y(n_1282) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
NOR3xp33_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1293), .C(n_1297), .Y(n_1291) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1315), .Y(n_1299) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1329), .Y(n_1547) );
AOI22xp5_ASAP7_75t_L g1329 ( .A1(n_1330), .A2(n_1385), .B1(n_1386), .B2(n_1546), .Y(n_1329) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1330), .Y(n_1546) );
HB1xp67_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
AND3x1_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1363), .C(n_1373), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1350), .Y(n_1333) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_1344), .A2(n_1514), .B1(n_1515), .B2(n_1528), .Y(n_1527) );
INVx2_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
OAI31xp33_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1365), .A3(n_1371), .B(n_1372), .Y(n_1363) );
INVxp67_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
OAI31xp33_ASAP7_75t_L g1459 ( .A1(n_1372), .A2(n_1460), .A3(n_1461), .B(n_1465), .Y(n_1459) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
OAI22xp5_ASAP7_75t_L g1441 ( .A1(n_1382), .A2(n_1442), .B1(n_1443), .B2(n_1444), .Y(n_1441) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
OAI22x1_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1475), .B1(n_1476), .B2(n_1545), .Y(n_1386) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1387), .Y(n_1545) );
XNOR2x1_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1432), .Y(n_1387) );
NAND3xp33_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1399), .C(n_1406), .Y(n_1389) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1423), .Y(n_1406) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
NAND3xp33_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1459), .C(n_1466), .Y(n_1433) );
NOR2xp33_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1451), .Y(n_1434) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1453), .Y(n_1801) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
INVx2_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
XNOR2x1_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1479), .Y(n_1477) );
NAND4xp75_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1489), .C(n_1513), .D(n_1516), .Y(n_1479) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
AOI211x1_ASAP7_75t_L g1489 ( .A1(n_1490), .A2(n_1497), .B(n_1498), .C(n_1508), .Y(n_1489) );
INVx2_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
NAND2x2_ASAP7_75t_L g1509 ( .A(n_1506), .B(n_1510), .Y(n_1509) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1509), .Y(n_1813) );
INVx2_ASAP7_75t_SL g1510 ( .A(n_1511), .Y(n_1510) );
INVx2_ASAP7_75t_SL g1815 ( .A(n_1512), .Y(n_1815) );
INVx4_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx2_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
AOI21xp33_ASAP7_75t_L g1526 ( .A1(n_1527), .A2(n_1529), .B(n_1532), .Y(n_1526) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
HB1xp67_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx2_ASAP7_75t_L g1782 ( .A(n_1534), .Y(n_1782) );
OAI21xp5_ASAP7_75t_SL g1535 ( .A1(n_1536), .A2(n_1538), .B(n_1541), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1802 ( .A(n_1537), .B(n_1803), .Y(n_1802) );
OAI221xp5_ASAP7_75t_L g1548 ( .A1(n_1549), .A2(n_1768), .B1(n_1771), .B2(n_1833), .C(n_1837), .Y(n_1548) );
AOI211xp5_ASAP7_75t_L g1549 ( .A1(n_1550), .A2(n_1673), .B(n_1680), .C(n_1746), .Y(n_1549) );
NAND5xp2_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1624), .C(n_1651), .D(n_1654), .E(n_1659), .Y(n_1550) );
AOI211xp5_ASAP7_75t_L g1551 ( .A1(n_1552), .A2(n_1582), .B(n_1591), .C(n_1619), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1569), .Y(n_1553) );
OAI321xp33_ASAP7_75t_L g1591 ( .A1(n_1554), .A2(n_1592), .A3(n_1599), .B1(n_1604), .B2(n_1605), .C(n_1610), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1554), .B(n_1570), .Y(n_1612) );
AND3x1_ASAP7_75t_L g1645 ( .A(n_1554), .B(n_1579), .C(n_1603), .Y(n_1645) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1554), .B(n_1637), .Y(n_1650) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1554), .B(n_1579), .Y(n_1670) );
OR2x2_ASAP7_75t_L g1697 ( .A(n_1554), .B(n_1698), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1554), .B(n_1600), .Y(n_1700) );
NAND2xp5_ASAP7_75t_L g1739 ( .A(n_1554), .B(n_1603), .Y(n_1739) );
INVx2_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1555), .B(n_1600), .Y(n_1609) );
BUFx2_ASAP7_75t_L g1615 ( .A(n_1555), .Y(n_1615) );
OR2x2_ASAP7_75t_L g1706 ( .A(n_1555), .B(n_1692), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1555), .B(n_1637), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1556), .B(n_1564), .Y(n_1555) );
AND2x4_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1559), .Y(n_1557) );
AND2x6_ASAP7_75t_L g1562 ( .A(n_1558), .B(n_1563), .Y(n_1562) );
AND2x6_ASAP7_75t_L g1565 ( .A(n_1558), .B(n_1566), .Y(n_1565) );
AND2x2_ASAP7_75t_L g1567 ( .A(n_1558), .B(n_1568), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1558), .B(n_1568), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1558), .B(n_1568), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1561), .Y(n_1559) );
INVx2_ASAP7_75t_L g1770 ( .A(n_1562), .Y(n_1770) );
HB1xp67_ASAP7_75t_L g1891 ( .A(n_1563), .Y(n_1891) );
INVx2_ASAP7_75t_L g1677 ( .A(n_1565), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1575), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1570), .B(n_1594), .Y(n_1593) );
NOR2xp33_ASAP7_75t_L g1627 ( .A(n_1570), .B(n_1628), .Y(n_1627) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1570), .Y(n_1662) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1570), .B(n_1632), .Y(n_1688) );
NOR2xp33_ASAP7_75t_L g1722 ( .A(n_1570), .B(n_1723), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1570), .B(n_1600), .Y(n_1757) );
INVx2_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1571), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1571), .B(n_1615), .Y(n_1614) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1571), .B(n_1584), .Y(n_1643) );
NAND2xp5_ASAP7_75t_L g1692 ( .A(n_1571), .B(n_1575), .Y(n_1692) );
NOR2xp33_ASAP7_75t_L g1694 ( .A(n_1571), .B(n_1695), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1571), .B(n_1595), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1573), .Y(n_1571) );
INVxp67_ASAP7_75t_L g1679 ( .A(n_1574), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1575), .B(n_1614), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1579), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1576), .B(n_1601), .Y(n_1600) );
INVx2_ASAP7_75t_L g1603 ( .A(n_1576), .Y(n_1603) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1576), .B(n_1615), .Y(n_1628) );
NAND3xp33_ASAP7_75t_L g1701 ( .A(n_1576), .B(n_1606), .C(n_1674), .Y(n_1701) );
OR2x2_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1578), .Y(n_1576) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1579), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1579), .B(n_1603), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1579), .B(n_1615), .Y(n_1687) );
OR2x2_ASAP7_75t_L g1723 ( .A(n_1579), .B(n_1615), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1581), .Y(n_1579) );
A2O1A1Ixp33_ASAP7_75t_L g1690 ( .A1(n_1582), .A2(n_1674), .B(n_1691), .C(n_1693), .Y(n_1690) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_1584), .B(n_1588), .Y(n_1583) );
CKINVDCx6p67_ASAP7_75t_R g1617 ( .A(n_1584), .Y(n_1617) );
OR2x2_ASAP7_75t_L g1621 ( .A(n_1584), .B(n_1622), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1584), .B(n_1632), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1584), .B(n_1588), .Y(n_1672) );
NAND2xp5_ASAP7_75t_L g1754 ( .A(n_1584), .B(n_1674), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1584), .B(n_1762), .Y(n_1761) );
OR2x6_ASAP7_75t_L g1584 ( .A(n_1585), .B(n_1587), .Y(n_1584) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1588), .Y(n_1598) );
INVx3_ASAP7_75t_L g1604 ( .A(n_1588), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1623 ( .A(n_1588), .B(n_1618), .Y(n_1623) );
OR2x2_ASAP7_75t_L g1626 ( .A(n_1588), .B(n_1595), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1588), .B(n_1617), .Y(n_1638) );
AND2x2_ASAP7_75t_L g1641 ( .A(n_1588), .B(n_1595), .Y(n_1641) );
OR2x2_ASAP7_75t_L g1656 ( .A(n_1588), .B(n_1617), .Y(n_1656) );
OAI221xp5_ASAP7_75t_L g1715 ( .A1(n_1588), .A2(n_1716), .B1(n_1717), .B2(n_1719), .C(n_1720), .Y(n_1715) );
OAI32xp33_ASAP7_75t_L g1742 ( .A1(n_1588), .A2(n_1604), .A3(n_1606), .B1(n_1697), .B2(n_1743), .Y(n_1742) );
AND2x4_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1590), .Y(n_1588) );
OAI32xp33_ASAP7_75t_L g1759 ( .A1(n_1592), .A2(n_1606), .A3(n_1646), .B1(n_1760), .B2(n_1761), .Y(n_1759) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1594), .Y(n_1646) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1594), .B(n_1617), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1598), .Y(n_1594) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1595), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1597), .Y(n_1595) );
OR2x2_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1602), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1600), .B(n_1614), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1601), .B(n_1603), .Y(n_1637) );
O2A1O1Ixp33_ASAP7_75t_L g1710 ( .A1(n_1601), .A2(n_1711), .B(n_1712), .C(n_1713), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1602), .B(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1602), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1602), .B(n_1615), .Y(n_1658) );
OAI322xp33_ASAP7_75t_L g1639 ( .A1(n_1603), .A2(n_1640), .A3(n_1642), .B1(n_1644), .B2(n_1646), .C1(n_1647), .C2(n_1649), .Y(n_1639) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1603), .B(n_1615), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1603), .B(n_1615), .Y(n_1744) );
CKINVDCx14_ASAP7_75t_R g1735 ( .A(n_1604), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1609), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_1606), .B(n_1700), .Y(n_1732) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1607), .B(n_1650), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1711 ( .A(n_1607), .B(n_1648), .Y(n_1711) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1607), .B(n_1700), .Y(n_1729) );
INVx2_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1657 ( .A(n_1608), .B(n_1658), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1608), .B(n_1637), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1608), .B(n_1648), .Y(n_1748) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1609), .B(n_1632), .Y(n_1765) );
OAI21xp5_ASAP7_75t_L g1610 ( .A1(n_1611), .A2(n_1613), .B(n_1616), .Y(n_1610) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1611), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1667 ( .A(n_1612), .B(n_1637), .Y(n_1667) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1613), .Y(n_1752) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1614), .Y(n_1635) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1616), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1717 ( .A(n_1616), .B(n_1718), .Y(n_1717) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1618), .Y(n_1616) );
NOR2xp33_ASAP7_75t_L g1625 ( .A(n_1617), .B(n_1626), .Y(n_1625) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1617), .B(n_1648), .Y(n_1647) );
NOR2xp33_ASAP7_75t_SL g1709 ( .A(n_1617), .B(n_1646), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1713 ( .A(n_1617), .B(n_1674), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1617), .B(n_1632), .Y(n_1727) );
INVx2_ASAP7_75t_L g1632 ( .A(n_1618), .Y(n_1632) );
NOR2xp33_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1621), .Y(n_1758) );
OAI22xp5_ASAP7_75t_L g1725 ( .A1(n_1622), .A2(n_1697), .B1(n_1726), .B2(n_1728), .Y(n_1725) );
OAI211xp5_ASAP7_75t_L g1733 ( .A1(n_1622), .A2(n_1699), .B(n_1734), .C(n_1740), .Y(n_1733) );
CKINVDCx6p67_ASAP7_75t_R g1622 ( .A(n_1623), .Y(n_1622) );
NAND2xp5_ASAP7_75t_L g1661 ( .A(n_1623), .B(n_1662), .Y(n_1661) );
AOI221xp5_ASAP7_75t_L g1624 ( .A1(n_1625), .A2(n_1627), .B1(n_1629), .B2(n_1638), .C(n_1639), .Y(n_1624) );
INVx2_ASAP7_75t_L g1648 ( .A(n_1626), .Y(n_1648) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1633), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1630), .B(n_1722), .Y(n_1721) );
A2O1A1Ixp33_ASAP7_75t_L g1749 ( .A1(n_1630), .A2(n_1698), .B(n_1699), .C(n_1750), .Y(n_1749) );
INVx2_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1631), .B(n_1652), .Y(n_1651) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1631), .B(n_1672), .Y(n_1671) );
NOR2xp33_ASAP7_75t_L g1751 ( .A(n_1631), .B(n_1752), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1631), .B(n_1729), .Y(n_1767) );
INVx2_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
OR2x2_ASAP7_75t_L g1716 ( .A(n_1632), .B(n_1634), .Y(n_1716) );
INVx1_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
OR2x2_ASAP7_75t_L g1634 ( .A(n_1635), .B(n_1636), .Y(n_1634) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1638), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1638), .B(n_1694), .Y(n_1693) );
OAI22xp5_ASAP7_75t_L g1665 ( .A1(n_1640), .A2(n_1666), .B1(n_1668), .B2(n_1671), .Y(n_1665) );
NOR2xp33_ASAP7_75t_L g1741 ( .A(n_1640), .B(n_1644), .Y(n_1741) );
INVx2_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
AOI22xp33_ASAP7_75t_L g1707 ( .A1(n_1641), .A2(n_1645), .B1(n_1708), .B2(n_1709), .Y(n_1707) );
CKINVDCx14_ASAP7_75t_R g1642 ( .A(n_1643), .Y(n_1642) );
INVx2_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
O2A1O1Ixp33_ASAP7_75t_L g1755 ( .A1(n_1652), .A2(n_1756), .B(n_1758), .C(n_1759), .Y(n_1755) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
NAND2xp5_ASAP7_75t_L g1654 ( .A(n_1655), .B(n_1657), .Y(n_1654) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
O2A1O1Ixp33_ASAP7_75t_L g1659 ( .A1(n_1658), .A2(n_1660), .B(n_1663), .C(n_1665), .Y(n_1659) );
NOR2xp33_ASAP7_75t_L g1760 ( .A(n_1658), .B(n_1700), .Y(n_1760) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
NOR2xp33_ASAP7_75t_L g1669 ( .A(n_1662), .B(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
OAI221xp5_ASAP7_75t_L g1682 ( .A1(n_1664), .A2(n_1683), .B1(n_1684), .B2(n_1689), .C(n_1690), .Y(n_1682) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
OAI31xp33_ASAP7_75t_L g1763 ( .A1(n_1672), .A2(n_1764), .A3(n_1765), .B(n_1766), .Y(n_1763) );
INVx2_ASAP7_75t_SL g1673 ( .A(n_1674), .Y(n_1673) );
INVx2_ASAP7_75t_SL g1719 ( .A(n_1674), .Y(n_1719) );
OAI22xp5_ASAP7_75t_SL g1675 ( .A1(n_1676), .A2(n_1677), .B1(n_1678), .B2(n_1679), .Y(n_1675) );
NAND3xp33_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1714), .C(n_1730), .Y(n_1680) );
NOR4xp25_ASAP7_75t_L g1681 ( .A(n_1682), .B(n_1696), .C(n_1704), .D(n_1710), .Y(n_1681) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
OAI21xp5_ASAP7_75t_L g1720 ( .A1(n_1685), .A2(n_1721), .B(n_1724), .Y(n_1720) );
NOR2xp33_ASAP7_75t_L g1685 ( .A(n_1686), .B(n_1688), .Y(n_1685) );
A2O1A1Ixp33_ASAP7_75t_L g1747 ( .A1(n_1686), .A2(n_1748), .B(n_1749), .C(n_1753), .Y(n_1747) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
AOI31xp33_ASAP7_75t_L g1696 ( .A1(n_1697), .A2(n_1699), .A3(n_1701), .B(n_1702), .Y(n_1696) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1697), .Y(n_1764) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
OAI21xp33_ASAP7_75t_L g1704 ( .A1(n_1705), .A2(n_1706), .B(n_1707), .Y(n_1704) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1708), .Y(n_1712) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1713), .Y(n_1724) );
NOR2xp33_ASAP7_75t_L g1714 ( .A(n_1715), .B(n_1725), .Y(n_1714) );
INVx3_ASAP7_75t_L g1745 ( .A(n_1719), .Y(n_1745) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
OAI31xp33_ASAP7_75t_L g1730 ( .A1(n_1731), .A2(n_1733), .A3(n_1742), .B(n_1745), .Y(n_1730) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1735), .B(n_1736), .Y(n_1734) );
NOR2xp33_ASAP7_75t_L g1736 ( .A(n_1737), .B(n_1739), .Y(n_1736) );
CKINVDCx14_ASAP7_75t_R g1737 ( .A(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1739), .Y(n_1762) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
CKINVDCx14_ASAP7_75t_R g1743 ( .A(n_1744), .Y(n_1743) );
NAND3xp33_ASAP7_75t_L g1746 ( .A(n_1747), .B(n_1755), .C(n_1763), .Y(n_1746) );
INVxp67_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
CKINVDCx20_ASAP7_75t_R g1768 ( .A(n_1769), .Y(n_1768) );
CKINVDCx20_ASAP7_75t_R g1769 ( .A(n_1770), .Y(n_1769) );
INVx2_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
NOR2x1_ASAP7_75t_L g1773 ( .A(n_1774), .B(n_1807), .Y(n_1773) );
A2O1A1Ixp33_ASAP7_75t_L g1774 ( .A1(n_1775), .A2(n_1785), .B(n_1804), .C(n_1805), .Y(n_1774) );
AOI211xp5_ASAP7_75t_SL g1775 ( .A1(n_1776), .A2(n_1777), .B(n_1778), .C(n_1780), .Y(n_1775) );
INVx3_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
NOR3xp33_ASAP7_75t_SL g1785 ( .A(n_1786), .B(n_1794), .C(n_1800), .Y(n_1785) );
INVx2_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1799), .Y(n_1798) );
NAND2xp5_ASAP7_75t_L g1807 ( .A(n_1808), .B(n_1817), .Y(n_1807) );
AOI22xp5_ASAP7_75t_L g1811 ( .A1(n_1812), .A2(n_1813), .B1(n_1814), .B2(n_1815), .Y(n_1811) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
AND2x4_ASAP7_75t_L g1826 ( .A(n_1827), .B(n_1828), .Y(n_1826) );
INVx2_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
BUFx3_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
BUFx2_ASAP7_75t_SL g1838 ( .A(n_1839), .Y(n_1838) );
BUFx3_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
INVxp33_ASAP7_75t_SL g1841 ( .A(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
HB1xp67_ASAP7_75t_L g1845 ( .A(n_1846), .Y(n_1845) );
OR2x2_ASAP7_75t_L g1846 ( .A(n_1847), .B(n_1860), .Y(n_1846) );
NAND3xp33_ASAP7_75t_L g1847 ( .A(n_1848), .B(n_1852), .C(n_1858), .Y(n_1847) );
NAND3xp33_ASAP7_75t_SL g1860 ( .A(n_1861), .B(n_1864), .C(n_1886), .Y(n_1860) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx2_ASAP7_75t_SL g1888 ( .A(n_1889), .Y(n_1888) );
INVx1_ASAP7_75t_L g1889 ( .A(n_1890), .Y(n_1889) );
OAI21xp5_ASAP7_75t_L g1890 ( .A1(n_1891), .A2(n_1892), .B(n_1893), .Y(n_1890) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1894), .Y(n_1893) );
endmodule