module fake_jpeg_31775_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_55),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_57),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g114 ( 
.A(n_59),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_19),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_89),
.Y(n_139)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g163 ( 
.A(n_85),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_1),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_2),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_96),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g126 ( 
.A(n_98),
.Y(n_126)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_25),
.B(n_2),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_103),
.Y(n_152)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_2),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_22),
.B1(n_23),
.B2(n_20),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_116),
.A2(n_148),
.B1(n_155),
.B2(n_66),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_52),
.A2(n_46),
.B1(n_23),
.B2(n_20),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g169 ( 
.A1(n_117),
.A2(n_154),
.B1(n_161),
.B2(n_63),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_46),
.B(n_23),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_122),
.A2(n_117),
.B(n_154),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_95),
.A2(n_20),
.B1(n_48),
.B2(n_40),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_53),
.A2(n_48),
.B1(n_40),
.B2(n_30),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_51),
.B1(n_43),
.B2(n_42),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_38),
.B1(n_37),
.B2(n_43),
.Y(n_173)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_56),
.A2(n_30),
.B1(n_51),
.B2(n_42),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_168),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_169),
.B(n_173),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_114),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_171),
.B(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_114),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_37),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_175),
.B(n_177),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_176),
.A2(n_204),
.B1(n_217),
.B2(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_33),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_178),
.B(n_199),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_191),
.Y(n_244)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_182),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_68),
.B1(n_61),
.B2(n_94),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_184),
.A2(n_186),
.B1(n_167),
.B2(n_130),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_107),
.A2(n_64),
.B1(n_72),
.B2(n_74),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_118),
.B(n_70),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_187),
.B(n_108),
.C(n_130),
.Y(n_241)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_148),
.A2(n_59),
.B1(n_97),
.B2(n_89),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_190),
.B(n_222),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_76),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_195),
.Y(n_238)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_205),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_32),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_202),
.Y(n_265)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_138),
.A2(n_38),
.B1(n_32),
.B2(n_39),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_119),
.B(n_39),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_206),
.Y(n_274)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_85),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_215),
.Y(n_247)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_211),
.Y(n_269)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_143),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_138),
.B(n_34),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_227),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_31),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_140),
.A2(n_29),
.B1(n_83),
.B2(n_27),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_125),
.B(n_102),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_219),
.B(n_8),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_125),
.B(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_223),
.B(n_224),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_111),
.B(n_98),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_126),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_142),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_226),
.A2(n_229),
.B1(n_3),
.B2(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_105),
.B(n_27),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_228),
.B(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_145),
.B1(n_128),
.B2(n_159),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_231),
.A2(n_232),
.B1(n_245),
.B2(n_250),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_193),
.A2(n_167),
.B1(n_129),
.B2(n_159),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_190),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_169),
.A2(n_136),
.B1(n_146),
.B2(n_166),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_256),
.B1(n_206),
.B2(n_228),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_193),
.A2(n_146),
.B1(n_27),
.B2(n_113),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_27),
.B1(n_113),
.B2(n_35),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_259),
.B1(n_277),
.B2(n_179),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_187),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_187),
.A2(n_27),
.B1(n_35),
.B2(n_6),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

OAI32xp33_ASAP7_75t_L g262 ( 
.A1(n_175),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_275),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_178),
.B(n_18),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_279),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_227),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_177),
.A2(n_10),
.B(n_11),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_12),
.B(n_13),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_173),
.Y(n_295)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_284),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_285),
.A2(n_289),
.B1(n_291),
.B2(n_296),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_252),
.A2(n_190),
.B(n_213),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_286),
.B(n_310),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_292),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_170),
.B1(n_199),
.B2(n_172),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_293),
.B(n_318),
.Y(n_358)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_295),
.B(n_303),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_173),
.B1(n_207),
.B2(n_181),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_248),
.B(n_244),
.C(n_272),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_298),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_240),
.A2(n_173),
.B1(n_188),
.B2(n_189),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_305),
.B1(n_306),
.B2(n_321),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_307),
.Y(n_342)
);

INVx11_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_201),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_302),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_239),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_261),
.B(n_192),
.C(n_185),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_309),
.C(n_323),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_253),
.A2(n_183),
.B1(n_182),
.B2(n_196),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_282),
.A2(n_206),
.B1(n_221),
.B2(n_220),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_281),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_251),
.B(n_180),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_314),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_234),
.B(n_194),
.C(n_195),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_282),
.A2(n_263),
.B(n_244),
.Y(n_310)
);

INVx5_ASAP7_75t_SL g311 ( 
.A(n_274),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_311),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_234),
.B(n_225),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_276),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_241),
.B(n_200),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_251),
.B(n_202),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_203),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_315),
.B(n_242),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_266),
.A2(n_216),
.B1(n_211),
.B2(n_210),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_316),
.A2(n_270),
.B1(n_269),
.B2(n_246),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_281),
.A2(n_218),
.B(n_212),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_317),
.A2(n_328),
.B(n_265),
.Y(n_341)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_271),
.B(n_222),
.C(n_13),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_230),
.B(n_168),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_324),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_320),
.B(n_326),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_248),
.A2(n_209),
.B1(n_13),
.B2(n_14),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_237),
.Y(n_322)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_12),
.C(n_14),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_15),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_258),
.B(n_15),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_329),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_275),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_256),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_277),
.B1(n_259),
.B2(n_245),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_232),
.A2(n_15),
.B(n_16),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_262),
.B(n_16),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_246),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_269),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_337),
.A2(n_340),
.B1(n_353),
.B2(n_354),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_365),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_296),
.A2(n_231),
.B1(n_258),
.B2(n_238),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_341),
.A2(n_362),
.B(n_315),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_343),
.A2(n_291),
.B1(n_306),
.B2(n_299),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_297),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_347),
.A2(n_351),
.B1(n_363),
.B2(n_366),
.Y(n_383)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_290),
.Y(n_349)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_297),
.A2(n_236),
.B1(n_267),
.B2(n_243),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_285),
.A2(n_265),
.B1(n_273),
.B2(n_264),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_289),
.A2(n_273),
.B1(n_243),
.B2(n_257),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_284),
.Y(n_355)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_264),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_359),
.B(n_361),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_287),
.B(n_280),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_295),
.A2(n_268),
.B1(n_257),
.B2(n_233),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_368),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_242),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_329),
.A2(n_268),
.B1(n_233),
.B2(n_255),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_312),
.B(n_276),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_283),
.A2(n_235),
.B1(n_255),
.B2(n_276),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_370),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_338),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_376),
.B(n_377),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_339),
.Y(n_377)
);

AND2x2_ASAP7_75t_SL g425 ( 
.A(n_379),
.B(n_402),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_304),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_382),
.C(n_387),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_308),
.Y(n_381)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_381),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_313),
.C(n_304),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_300),
.Y(n_384)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_309),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_313),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_408),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_341),
.A2(n_298),
.B(n_288),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_391),
.A2(n_395),
.B(n_399),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_313),
.C(n_288),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_331),
.C(n_363),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_332),
.A2(n_287),
.B1(n_298),
.B2(n_288),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_394),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_367),
.A2(n_328),
.B(n_286),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_335),
.A2(n_324),
.B(n_292),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_332),
.A2(n_315),
.B1(n_314),
.B2(n_317),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_396),
.B(n_404),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_330),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_397),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_319),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_403),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_352),
.A2(n_310),
.B(n_315),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_348),
.Y(n_400)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_400),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_365),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_401),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_358),
.A2(n_305),
.B(n_316),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_348),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_355),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_405),
.A2(n_354),
.B1(n_370),
.B2(n_323),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_336),
.A2(n_337),
.B1(n_340),
.B2(n_360),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_406),
.B(n_321),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_356),
.A2(n_318),
.B(n_325),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_407),
.B(n_360),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_368),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_410),
.B(n_432),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_331),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_422),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_374),
.A2(n_389),
.B1(n_396),
.B2(n_406),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_414),
.A2(n_429),
.B1(n_405),
.B2(n_383),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_420),
.C(n_375),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_417),
.Y(n_445)
);

OAI32xp33_ASAP7_75t_L g418 ( 
.A1(n_376),
.A2(n_350),
.A3(n_356),
.B1(n_351),
.B2(n_336),
.Y(n_418)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_427),
.B1(n_434),
.B2(n_389),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_333),
.C(n_371),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_382),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_391),
.A2(n_366),
.B1(n_323),
.B2(n_333),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_381),
.B(n_322),
.Y(n_431)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_431),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_373),
.Y(n_432)
);

OAI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_374),
.A2(n_357),
.B1(n_311),
.B2(n_334),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_386),
.Y(n_435)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_357),
.Y(n_436)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_384),
.B(n_346),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_438),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_377),
.B(n_346),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_375),
.B(n_327),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_439),
.B(n_408),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g442 ( 
.A(n_413),
.B(n_393),
.CI(n_392),
.CON(n_442),
.SN(n_442)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_453),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_443),
.A2(n_430),
.B1(n_410),
.B2(n_425),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_421),
.A2(n_412),
.B(n_399),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_444),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_446),
.A2(n_452),
.B1(n_456),
.B2(n_459),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_411),
.A2(n_388),
.B1(n_383),
.B2(n_407),
.Y(n_447)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_448),
.B(n_460),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_415),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_394),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_448),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_394),
.B1(n_379),
.B2(n_404),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_426),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_454),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_427),
.A2(n_403),
.B1(n_402),
.B2(n_400),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_395),
.C(n_386),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_462),
.C(n_464),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_378),
.B1(n_385),
.B2(n_349),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_433),
.B(n_311),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_426),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_432),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_409),
.B(n_385),
.C(n_294),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_409),
.B(n_378),
.C(n_301),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_414),
.A2(n_301),
.B1(n_369),
.B2(n_17),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_469),
.B(n_481),
.C(n_482),
.Y(n_502)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_421),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_473),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_474),
.A2(n_416),
.B1(n_465),
.B2(n_429),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_463),
.Y(n_479)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_479),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_420),
.C(n_439),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_412),
.C(n_423),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_440),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_483),
.B(n_438),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_425),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_485),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_423),
.C(n_436),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_417),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_SL g504 ( 
.A(n_486),
.B(n_489),
.Y(n_504)
);

INVx11_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_488),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_425),
.C(n_437),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_476),
.A2(n_455),
.B1(n_443),
.B2(n_457),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_490),
.A2(n_488),
.B1(n_485),
.B2(n_424),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_472),
.A2(n_455),
.B(n_463),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_492),
.Y(n_515)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_493),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_474),
.A2(n_444),
.B(n_452),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_494),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_487),
.A2(n_456),
.B(n_451),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_495),
.B(n_497),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_468),
.A2(n_446),
.B(n_457),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_471),
.A2(n_442),
.B1(n_441),
.B2(n_416),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_499),
.Y(n_519)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_505),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_482),
.A2(n_425),
.B(n_465),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_507),
.Y(n_512)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_478),
.C(n_469),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_508),
.A2(n_517),
.B(n_521),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_491),
.A2(n_442),
.B1(n_486),
.B2(n_489),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_498),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_516),
.B(n_518),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_478),
.C(n_481),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_484),
.Y(n_518)
);

OAI31xp67_ASAP7_75t_L g520 ( 
.A1(n_492),
.A2(n_418),
.A3(n_424),
.B(n_431),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_520),
.A2(n_499),
.B1(n_454),
.B2(n_467),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_501),
.B(n_473),
.C(n_475),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_515),
.A2(n_500),
.B1(n_496),
.B2(n_494),
.Y(n_522)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_522),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_490),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_523),
.B(n_525),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_495),
.B(n_497),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_524),
.A2(n_532),
.B(n_510),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_493),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_527),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_503),
.C(n_506),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_528),
.B(n_529),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_519),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_435),
.Y(n_532)
);

O2A1O1Ixp33_ASAP7_75t_SL g534 ( 
.A1(n_522),
.A2(n_510),
.B(n_520),
.C(n_511),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_534),
.A2(n_536),
.B(n_527),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_SL g536 ( 
.A(n_531),
.B(n_504),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_538),
.A2(n_524),
.B(n_475),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_540),
.A2(n_541),
.B(n_543),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_539),
.B(n_530),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_533),
.B(n_521),
.C(n_503),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_542),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_537),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_547),
.C(n_369),
.Y(n_548)
);

OAI31xp33_ASAP7_75t_SL g547 ( 
.A1(n_544),
.A2(n_524),
.A3(n_535),
.B(n_428),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_548),
.Y(n_549)
);

O2A1O1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_17),
.B(n_18),
.C(n_545),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_550),
.B(n_17),
.Y(n_551)
);


endmodule