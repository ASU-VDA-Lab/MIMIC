module real_aes_2445_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_798, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_798;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g212 ( .A(n_0), .B(n_134), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_1), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_2), .B(n_140), .Y(n_493) );
XOR2xp5_ASAP7_75t_L g108 ( .A(n_3), .B(n_31), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_4), .B(n_130), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_5), .B(n_140), .Y(n_153) );
INVx1_ASAP7_75t_L g127 ( .A(n_6), .Y(n_127) );
NAND2xp33_ASAP7_75t_SL g204 ( .A(n_7), .B(n_138), .Y(n_204) );
INVx1_ASAP7_75t_L g185 ( .A(n_8), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_9), .A2(n_45), .B1(n_468), .B2(n_469), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_9), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g794 ( .A(n_10), .Y(n_794) );
AND2x2_ASAP7_75t_L g151 ( .A(n_11), .B(n_144), .Y(n_151) );
AND2x2_ASAP7_75t_L g525 ( .A(n_12), .B(n_178), .Y(n_525) );
AND2x2_ASAP7_75t_L g533 ( .A(n_13), .B(n_201), .Y(n_533) );
INVx2_ASAP7_75t_L g145 ( .A(n_14), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_15), .B(n_130), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_16), .Y(n_446) );
AOI221x1_ASAP7_75t_L g198 ( .A1(n_17), .A2(n_122), .B1(n_199), .B2(n_201), .C(n_203), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_18), .B(n_140), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_19), .B(n_140), .Y(n_506) );
INVx1_ASAP7_75t_L g450 ( .A(n_20), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_21), .A2(n_91), .B1(n_140), .B2(n_186), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_22), .A2(n_122), .B(n_155), .Y(n_154) );
AOI221xp5_ASAP7_75t_SL g165 ( .A1(n_23), .A2(n_38), .B1(n_122), .B2(n_140), .C(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_24), .B(n_134), .Y(n_156) );
AOI22xp5_ASAP7_75t_SL g438 ( .A1(n_25), .A2(n_79), .B1(n_439), .B2(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_25), .Y(n_440) );
OR2x2_ASAP7_75t_L g146 ( .A(n_26), .B(n_90), .Y(n_146) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_26), .A2(n_90), .B(n_145), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_27), .B(n_130), .Y(n_177) );
INVxp67_ASAP7_75t_L g197 ( .A(n_28), .Y(n_197) );
AND2x2_ASAP7_75t_L g228 ( .A(n_29), .B(n_143), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_30), .A2(n_122), .B(n_211), .Y(n_210) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_31), .A2(n_201), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_32), .B(n_130), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_33), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_34), .A2(n_122), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_35), .B(n_130), .Y(n_492) );
AND2x2_ASAP7_75t_L g123 ( .A(n_36), .B(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g138 ( .A(n_36), .B(n_127), .Y(n_138) );
INVx1_ASAP7_75t_L g193 ( .A(n_36), .Y(n_193) );
OR2x6_ASAP7_75t_L g448 ( .A(n_37), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_39), .B(n_140), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_40), .A2(n_83), .B1(n_122), .B2(n_191), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_41), .B(n_130), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_42), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_43), .B(n_140), .Y(n_558) );
XOR2xp5_ASAP7_75t_L g463 ( .A(n_44), .B(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_45), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_46), .B(n_134), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_47), .A2(n_122), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g215 ( .A(n_48), .B(n_143), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_49), .B(n_134), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_50), .B(n_143), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_51), .B(n_140), .Y(n_481) );
INVx1_ASAP7_75t_L g126 ( .A(n_52), .Y(n_126) );
INVx1_ASAP7_75t_L g136 ( .A(n_52), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_53), .B(n_130), .Y(n_531) );
AND2x2_ASAP7_75t_L g497 ( .A(n_54), .B(n_143), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_55), .B(n_140), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_56), .B(n_134), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_57), .B(n_134), .Y(n_491) );
AND2x2_ASAP7_75t_L g147 ( .A(n_58), .B(n_143), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_59), .B(n_140), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_60), .B(n_130), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_61), .B(n_140), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_62), .A2(n_122), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_63), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_64), .B(n_144), .Y(n_180) );
AND2x2_ASAP7_75t_L g512 ( .A(n_65), .B(n_144), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_66), .A2(n_122), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_67), .B(n_130), .Y(n_157) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_68), .B(n_178), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_69), .B(n_134), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_70), .B(n_134), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_71), .A2(n_95), .B1(n_122), .B2(n_191), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_72), .B(n_130), .Y(n_509) );
INVx1_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
INVx1_ASAP7_75t_L g132 ( .A(n_73), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_74), .B(n_134), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_75), .A2(n_122), .B(n_501), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_76), .A2(n_122), .B(n_560), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_77), .A2(n_122), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g494 ( .A(n_78), .B(n_144), .Y(n_494) );
INVx1_ASAP7_75t_L g439 ( .A(n_79), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_80), .B(n_143), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_81), .B(n_140), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_82), .A2(n_85), .B1(n_140), .B2(n_186), .Y(n_263) );
INVx1_ASAP7_75t_L g451 ( .A(n_84), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_86), .B(n_134), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_87), .B(n_134), .Y(n_168) );
AND2x2_ASAP7_75t_L g563 ( .A(n_88), .B(n_178), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g121 ( .A1(n_89), .A2(n_122), .B(n_128), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_92), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_93), .B(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_94), .A2(n_122), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_96), .B(n_130), .Y(n_561) );
INVxp67_ASAP7_75t_L g200 ( .A(n_97), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_98), .B(n_140), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_99), .B(n_130), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_100), .A2(n_122), .B(n_175), .Y(n_174) );
BUFx2_ASAP7_75t_L g511 ( .A(n_101), .Y(n_511) );
BUFx2_ASAP7_75t_SL g460 ( .A(n_102), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_102), .B(n_452), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_103), .A2(n_465), .B1(n_466), .B2(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_103), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_787), .B(n_795), .Y(n_104) );
OA22x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_456), .B1(n_461), .B2(n_462), .Y(n_105) );
OAI21xp5_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_441), .B(n_452), .Y(n_106) );
XNOR2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AOI22x1_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_111), .B1(n_437), .B2(n_438), .Y(n_109) );
INVx4_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_111), .A2(n_471), .B1(n_473), .B2(n_773), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_111), .B(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_376), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_269), .C(n_320), .Y(n_112) );
OAI211xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_159), .B(n_216), .C(n_247), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_148), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_118), .B(n_221), .Y(n_384) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g229 ( .A(n_119), .B(n_150), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_119), .B(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g246 ( .A(n_119), .B(n_236), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_119), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g283 ( .A(n_119), .B(n_259), .Y(n_283) );
INVx2_ASAP7_75t_L g309 ( .A(n_119), .Y(n_309) );
AND2x4_ASAP7_75t_L g318 ( .A(n_119), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g423 ( .A(n_119), .B(n_290), .Y(n_423) );
AO21x2_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_142), .B(n_147), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_139), .Y(n_120) );
AND2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
BUFx3_ASAP7_75t_L g190 ( .A(n_123), .Y(n_190) );
AND2x6_ASAP7_75t_L g134 ( .A(n_124), .B(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g195 ( .A(n_124), .Y(n_195) );
AND2x4_ASAP7_75t_L g191 ( .A(n_125), .B(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x4_ASAP7_75t_L g130 ( .A(n_126), .B(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g188 ( .A(n_126), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_127), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B(n_137), .Y(n_128) );
AND2x4_ASAP7_75t_L g141 ( .A(n_131), .B(n_135), .Y(n_141) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_134), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_137), .A2(n_156), .B(n_157), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_137), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_137), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_137), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_137), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_137), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_137), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_137), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_137), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_137), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_137), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_137), .A2(n_561), .B(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g140 ( .A(n_138), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g205 ( .A(n_141), .Y(n_205) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_142), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_142), .A2(n_222), .B(n_228), .Y(n_236) );
AOI21x1_ASAP7_75t_L g518 ( .A1(n_142), .A2(n_519), .B(n_525), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_143), .Y(n_142) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_143), .A2(n_165), .B(n_169), .Y(n_164) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_143), .A2(n_540), .B(n_541), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_143), .A2(n_558), .B(n_559), .Y(n_557) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g158 ( .A(n_145), .B(n_146), .Y(n_158) );
AND2x2_ASAP7_75t_L g307 ( .A(n_148), .B(n_308), .Y(n_307) );
OAI32xp33_ASAP7_75t_L g390 ( .A1(n_148), .A2(n_312), .A3(n_316), .B1(n_323), .B2(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_148), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g244 ( .A(n_149), .B(n_245), .Y(n_244) );
NAND3xp33_ASAP7_75t_L g317 ( .A(n_149), .B(n_239), .C(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g343 ( .A(n_149), .B(n_246), .Y(n_343) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_150), .Y(n_233) );
INVx5_ASAP7_75t_L g268 ( .A(n_150), .Y(n_268) );
AND2x4_ASAP7_75t_L g324 ( .A(n_150), .B(n_236), .Y(n_324) );
OR2x2_ASAP7_75t_L g339 ( .A(n_150), .B(n_259), .Y(n_339) );
OR2x2_ASAP7_75t_L g365 ( .A(n_150), .B(n_221), .Y(n_365) );
AND2x2_ASAP7_75t_L g373 ( .A(n_150), .B(n_319), .Y(n_373) );
AND2x4_ASAP7_75t_SL g398 ( .A(n_150), .B(n_318), .Y(n_398) );
OR2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_158), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_158), .B(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_158), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_158), .B(n_200), .Y(n_199) );
NOR3xp33_ASAP7_75t_L g203 ( .A(n_158), .B(n_204), .C(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_158), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_158), .A2(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_160), .B(n_318), .Y(n_394) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_170), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_161), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OR2x6_ASAP7_75t_SL g218 ( .A(n_162), .B(n_219), .Y(n_218) );
INVxp67_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g243 ( .A(n_163), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_163), .B(n_278), .Y(n_296) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_163), .Y(n_434) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g251 ( .A(n_164), .Y(n_251) );
AND2x2_ASAP7_75t_L g276 ( .A(n_164), .B(n_207), .Y(n_276) );
INVx2_ASAP7_75t_L g304 ( .A(n_164), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_164), .B(n_171), .Y(n_345) );
BUFx3_ASAP7_75t_L g369 ( .A(n_164), .Y(n_369) );
OR2x2_ASAP7_75t_L g381 ( .A(n_164), .B(n_171), .Y(n_381) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_164), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_170), .A2(n_412), .B1(n_415), .B2(n_416), .Y(n_411) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_181), .Y(n_170) );
INVx1_ASAP7_75t_L g239 ( .A(n_171), .Y(n_239) );
OR2x2_ASAP7_75t_L g250 ( .A(n_171), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
AND2x4_ASAP7_75t_SL g274 ( .A(n_171), .B(n_182), .Y(n_274) );
AND2x4_ASAP7_75t_L g279 ( .A(n_171), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g288 ( .A(n_171), .Y(n_288) );
OR2x2_ASAP7_75t_L g294 ( .A(n_171), .B(n_182), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_171), .B(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_171), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_171), .B(n_276), .Y(n_410) );
OR2x2_ASAP7_75t_L g426 ( .A(n_171), .B(n_329), .Y(n_426) );
OR2x6_ASAP7_75t_L g171 ( .A(n_172), .B(n_180), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_178), .Y(n_172) );
INVx2_ASAP7_75t_SL g261 ( .A(n_178), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_178), .A2(n_506), .B(n_507), .Y(n_505) );
BUFx4f_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_181), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g252 ( .A(n_181), .Y(n_252) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_181), .B(n_243), .Y(n_359) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_206), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_182), .B(n_207), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_182), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_182), .B(n_251), .Y(n_255) );
INVx3_ASAP7_75t_L g280 ( .A(n_182), .Y(n_280) );
INVx1_ASAP7_75t_L g313 ( .A(n_182), .Y(n_313) );
AND2x2_ASAP7_75t_L g393 ( .A(n_182), .B(n_257), .Y(n_393) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_198), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_186), .B1(n_191), .B2(n_196), .Y(n_183) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_190), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2x1p5_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g487 ( .A(n_201), .Y(n_487) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI21x1_ASAP7_75t_L g208 ( .A1(n_202), .A2(n_209), .B(n_215), .Y(n_208) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_202), .A2(n_527), .B(n_533), .Y(n_526) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_207), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g278 ( .A(n_207), .Y(n_278) );
AND2x2_ASAP7_75t_L g303 ( .A(n_207), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g329 ( .A(n_207), .B(n_251), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_207), .B(n_280), .Y(n_346) );
INVx1_ASAP7_75t_L g352 ( .A(n_207), .Y(n_352) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_214), .Y(n_209) );
AOI222xp33_ASAP7_75t_SL g216 ( .A1(n_217), .A2(n_220), .B1(n_230), .B2(n_237), .C1(n_240), .C2(n_244), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_229), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_221), .B(n_290), .Y(n_341) );
AND2x4_ASAP7_75t_L g357 ( .A(n_221), .B(n_268), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_227), .Y(n_222) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_232), .B(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g282 ( .A(n_233), .B(n_283), .Y(n_282) );
AOI222xp33_ASAP7_75t_L g247 ( .A1(n_234), .A2(n_248), .B1(n_253), .B2(n_258), .C1(n_266), .C2(n_798), .Y(n_247) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g386 ( .A(n_235), .B(n_290), .Y(n_386) );
OR2x2_ASAP7_75t_L g429 ( .A(n_235), .B(n_335), .Y(n_429) );
AND2x2_ASAP7_75t_L g258 ( .A(n_236), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g319 ( .A(n_236), .Y(n_319) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_236), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_237), .A2(n_348), .B(n_353), .C(n_354), .Y(n_347) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g375 ( .A(n_239), .Y(n_375) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
AND2x2_ASAP7_75t_L g289 ( .A(n_245), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g298 ( .A(n_245), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OAI31xp33_ASAP7_75t_L g340 ( .A1(n_248), .A2(n_266), .A3(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g342 ( .A1(n_249), .A2(n_299), .B(n_343), .C(n_344), .Y(n_342) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
OR2x2_ASAP7_75t_L g331 ( .A(n_250), .B(n_280), .Y(n_331) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
BUFx2_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
AND2x2_ASAP7_75t_L g308 ( .A(n_259), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_260), .Y(n_290) );
AOI21x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_265), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_268), .B(n_325), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_281), .B(n_284), .C(n_306), .Y(n_269) );
INVxp33_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_272), .B(n_277), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g310 ( .A(n_274), .B(n_303), .Y(n_310) );
OR2x2_ASAP7_75t_L g286 ( .A(n_275), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g316 ( .A(n_275), .B(n_290), .Y(n_316) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g392 ( .A(n_276), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g415 ( .A(n_277), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_279), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_279), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g427 ( .A(n_279), .B(n_303), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_279), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g370 ( .A(n_280), .B(n_352), .Y(n_370) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AOI322xp5_ASAP7_75t_L g424 ( .A1(n_283), .A2(n_303), .A3(n_357), .B1(n_382), .B2(n_425), .C1(n_427), .C2(n_428), .Y(n_424) );
AOI211xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_289), .B(n_291), .C(n_300), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_287), .B(n_315), .Y(n_337) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g302 ( .A(n_288), .B(n_303), .Y(n_302) );
NOR2x1p5_ASAP7_75t_L g368 ( .A(n_288), .B(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_288), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_289), .A2(n_307), .B(n_310), .C(n_311), .Y(n_306) );
AND2x4_ASAP7_75t_L g325 ( .A(n_290), .B(n_309), .Y(n_325) );
INVx2_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_290), .B(n_324), .Y(n_355) );
AND2x2_ASAP7_75t_L g397 ( .A(n_290), .B(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_290), .B(n_414), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_290), .B(n_318), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B(n_297), .Y(n_291) );
AND2x2_ASAP7_75t_L g387 ( .A(n_293), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g315 ( .A(n_296), .Y(n_315) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_308), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g402 ( .A(n_308), .Y(n_402) );
O2A1O1Ixp33_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_314), .B(n_316), .C(n_317), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_315), .Y(n_399) );
INVx3_ASAP7_75t_SL g414 ( .A(n_318), .Y(n_414) );
NAND5xp2_ASAP7_75t_L g320 ( .A(n_321), .B(n_340), .C(n_347), .D(n_360), .E(n_371), .Y(n_320) );
AOI222xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_326), .B1(n_330), .B2(n_332), .C1(n_336), .C2(n_338), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_323), .A2(n_404), .B1(n_408), .B2(n_409), .Y(n_403) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g353 ( .A(n_324), .B(n_325), .Y(n_353) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_334), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_335), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g372 ( .A(n_335), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g383 ( .A(n_335), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g413 ( .A(n_339), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g361 ( .A(n_346), .Y(n_361) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B(n_358), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_357), .A2(n_361), .B1(n_362), .B2(n_366), .Y(n_360) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_357), .Y(n_408) );
INVx2_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g374 ( .A(n_359), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g379 ( .A(n_361), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_SL g407 ( .A(n_370), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
NOR3xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_395), .C(n_418), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_378), .B(n_394), .Y(n_377) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_382), .B1(n_385), .B2(n_387), .C(n_390), .Y(n_378) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g419 ( .A(n_381), .B(n_407), .Y(n_419) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
OAI321xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_399), .A3(n_400), .B1(n_402), .B2(n_403), .C(n_411), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_409), .A2(n_431), .B1(n_435), .B2(n_436), .Y(n_430) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_420), .B(n_424), .C(n_430), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp33_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
CKINVDCx11_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g455 ( .A(n_445), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
AND2x6_ASAP7_75t_SL g472 ( .A(n_446), .B(n_448), .Y(n_472) );
OR2x6_ASAP7_75t_SL g773 ( .A(n_446), .B(n_447), .Y(n_773) );
OR2x2_ASAP7_75t_L g786 ( .A(n_446), .B(n_448), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
CKINVDCx11_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
CKINVDCx8_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
AO221x1_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_470), .B1(n_774), .B2(n_782), .C(n_783), .Y(n_462) );
INVx1_ASAP7_75t_L g782 ( .A(n_463), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
CKINVDCx11_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_472), .Y(n_781) );
INVx4_ASAP7_75t_L g778 ( .A(n_473), .Y(n_778) );
AND3x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_651), .C(n_747), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_593), .C(n_620), .Y(n_474) );
OAI211xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_513), .B(n_542), .C(n_566), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_495), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_477), .A2(n_544), .B(n_548), .C(n_554), .Y(n_543) );
OR2x2_ASAP7_75t_L g666 ( .A(n_477), .B(n_603), .Y(n_666) );
INVx2_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g633 ( .A(n_478), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_478), .B(n_604), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_478), .B(n_749), .Y(n_764) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_486), .Y(n_478) );
AND2x2_ASAP7_75t_L g550 ( .A(n_479), .B(n_496), .Y(n_550) );
INVx1_ASAP7_75t_L g570 ( .A(n_479), .Y(n_570) );
OR2x2_ASAP7_75t_L g585 ( .A(n_479), .B(n_504), .Y(n_585) );
INVx2_ASAP7_75t_L g591 ( .A(n_479), .Y(n_591) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_479), .Y(n_646) );
INVx1_ASAP7_75t_L g723 ( .A(n_479), .Y(n_723) );
NOR2x1_ASAP7_75t_SL g572 ( .A(n_486), .B(n_504), .Y(n_572) );
AND2x2_ASAP7_75t_L g602 ( .A(n_486), .B(n_591), .Y(n_602) );
AO21x1_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_488), .B(n_494), .Y(n_486) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_487), .A2(n_488), .B(n_494), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_493), .Y(n_488) );
OR2x2_ASAP7_75t_L g596 ( .A(n_495), .B(n_597), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_495), .B(n_703), .Y(n_702) );
INVx3_ASAP7_75t_L g724 ( .A(n_495), .Y(n_724) );
NAND2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .Y(n_495) );
OR2x2_ASAP7_75t_SL g584 ( .A(n_496), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g588 ( .A(n_496), .Y(n_588) );
INVx4_ASAP7_75t_L g604 ( .A(n_496), .Y(n_604) );
OR2x2_ASAP7_75t_L g619 ( .A(n_496), .B(n_552), .Y(n_619) );
AND2x2_ASAP7_75t_L g658 ( .A(n_496), .B(n_572), .Y(n_658) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_496), .Y(n_670) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AND2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g603 ( .A(n_504), .B(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g618 ( .A(n_504), .Y(n_618) );
AND2x2_ASAP7_75t_L g634 ( .A(n_504), .B(n_604), .Y(n_634) );
AND2x2_ASAP7_75t_L g647 ( .A(n_504), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g679 ( .A(n_504), .B(n_591), .Y(n_679) );
INVx2_ASAP7_75t_SL g749 ( .A(n_504), .Y(n_749) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_512), .Y(n_504) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NOR2xp67_ASAP7_75t_L g514 ( .A(n_515), .B(n_534), .Y(n_514) );
OAI211xp5_ASAP7_75t_L g620 ( .A1(n_515), .A2(n_621), .B(n_625), .C(n_641), .Y(n_620) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g716 ( .A(n_516), .B(n_555), .Y(n_716) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
INVx2_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
AND2x4_ASAP7_75t_SL g576 ( .A(n_517), .B(n_556), .Y(n_576) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_517), .Y(n_580) );
AND2x2_ASAP7_75t_L g638 ( .A(n_517), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g712 ( .A(n_517), .Y(n_712) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_518), .Y(n_614) );
AND2x2_ASAP7_75t_L g657 ( .A(n_518), .B(n_526), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_524), .Y(n_519) );
INVx2_ASAP7_75t_L g547 ( .A(n_526), .Y(n_547) );
AND2x2_ASAP7_75t_L g607 ( .A(n_526), .B(n_556), .Y(n_607) );
INVx2_ASAP7_75t_L g639 ( .A(n_526), .Y(n_639) );
OR2x2_ASAP7_75t_L g662 ( .A(n_526), .B(n_537), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_534), .B(n_579), .Y(n_686) );
AND2x2_ASAP7_75t_L g720 ( .A(n_534), .B(n_656), .Y(n_720) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI31xp33_ASAP7_75t_SL g641 ( .A1(n_535), .A2(n_622), .A3(n_642), .B(n_649), .Y(n_641) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_536), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx3_ASAP7_75t_L g575 ( .A(n_537), .Y(n_575) );
AND2x2_ASAP7_75t_L g592 ( .A(n_537), .B(n_555), .Y(n_592) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AND2x4_ASAP7_75t_L g582 ( .A(n_538), .B(n_539), .Y(n_582) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g727 ( .A(n_545), .Y(n_727) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_547), .B(n_556), .Y(n_609) );
AND2x2_ASAP7_75t_L g650 ( .A(n_547), .B(n_565), .Y(n_650) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g630 ( .A(n_551), .B(n_588), .Y(n_630) );
AND2x2_ASAP7_75t_L g589 ( .A(n_552), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_552), .Y(n_598) );
INVx2_ASAP7_75t_L g648 ( .A(n_552), .Y(n_648) );
AND2x2_ASAP7_75t_L g738 ( .A(n_552), .B(n_723), .Y(n_738) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g744 ( .A(n_554), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_555), .B(n_564), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_555), .B(n_614), .Y(n_683) );
AND2x2_ASAP7_75t_L g731 ( .A(n_555), .B(n_657), .Y(n_731) );
INVx4_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g640 ( .A(n_556), .B(n_612), .Y(n_640) );
AND2x2_ASAP7_75t_L g649 ( .A(n_556), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g661 ( .A(n_556), .Y(n_661) );
BUFx2_ASAP7_75t_L g677 ( .A(n_556), .Y(n_677) );
AND2x4_ASAP7_75t_L g711 ( .A(n_556), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g756 ( .A(n_556), .B(n_657), .Y(n_756) );
OR2x6_ASAP7_75t_L g556 ( .A(n_557), .B(n_563), .Y(n_556) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_573), .B1(n_577), .B2(n_583), .C1(n_586), .C2(n_592), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_568), .A2(n_632), .B1(n_635), .B2(n_640), .Y(n_631) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g615 ( .A(n_569), .B(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_SL g629 ( .A(n_569), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_569), .B(n_634), .Y(n_767) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g728 ( .A(n_570), .B(n_634), .Y(n_728) );
OR2x2_ASAP7_75t_L g705 ( .A(n_571), .B(n_587), .Y(n_705) );
OR2x2_ASAP7_75t_L g713 ( .A(n_571), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g697 ( .A(n_572), .B(n_590), .Y(n_697) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
OR2x2_ASAP7_75t_L g605 ( .A(n_575), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g755 ( .A(n_575), .B(n_756), .Y(n_755) );
AND2x2_ASAP7_75t_L g706 ( .A(n_576), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_576), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_SL g741 ( .A(n_576), .Y(n_741) );
INVxp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx2_ASAP7_75t_L g726 ( .A(n_579), .Y(n_726) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g628 ( .A(n_580), .B(n_607), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_581), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g627 ( .A(n_581), .Y(n_627) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_581), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g730 ( .A(n_581), .B(n_602), .Y(n_730) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g664 ( .A(n_582), .B(n_650), .Y(n_664) );
AND2x2_ASAP7_75t_L g707 ( .A(n_582), .B(n_639), .Y(n_707) );
AND2x4_ASAP7_75t_L g622 ( .A(n_583), .B(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g763 ( .A(n_585), .B(n_619), .Y(n_763) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_587), .B(n_602), .Y(n_746) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_588), .B(n_602), .Y(n_668) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_588), .A2(n_629), .B(n_730), .C(n_731), .Y(n_729) );
AND2x2_ASAP7_75t_L g760 ( .A(n_588), .B(n_738), .Y(n_760) );
INVx1_ASAP7_75t_L g671 ( .A(n_589), .Y(n_671) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_592), .B(n_656), .Y(n_655) );
OAI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_605), .B(n_608), .Y(n_593) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_595), .B(n_599), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_596), .A2(n_749), .B1(n_750), .B2(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g624 ( .A(n_598), .Y(n_624) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g645 ( .A(n_604), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g696 ( .A(n_604), .Y(n_696) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_615), .Y(n_608) );
INVx1_ASAP7_75t_L g687 ( .A(n_609), .Y(n_687) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_629), .B(n_631), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OR2x2_ASAP7_75t_L g672 ( .A(n_627), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g709 ( .A(n_627), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_627), .B(n_657), .Y(n_745) );
INVx1_ASAP7_75t_L g765 ( .A(n_628), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_630), .A2(n_733), .B1(n_736), .B2(n_739), .C(n_742), .Y(n_732) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI321xp33_ASAP7_75t_L g753 ( .A1(n_635), .A2(n_670), .A3(n_754), .B1(n_757), .B2(n_759), .C(n_761), .Y(n_753) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g694 ( .A(n_639), .Y(n_694) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g688 ( .A(n_644), .Y(n_688) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g714 ( .A(n_645), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_647), .A2(n_675), .B1(n_679), .B2(n_680), .C(n_685), .Y(n_674) );
INVxp67_ASAP7_75t_L g703 ( .A(n_648), .Y(n_703) );
INVx1_ASAP7_75t_L g673 ( .A(n_650), .Y(n_673) );
NOR2xp67_ASAP7_75t_L g651 ( .A(n_652), .B(n_698), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_674), .C(n_689), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_658), .B1(n_659), .B2(n_665), .C(n_667), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g772 ( .A(n_657), .Y(n_772) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_660), .B(n_663), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_661), .B(n_707), .Y(n_752) );
INVx2_ASAP7_75t_SL g684 ( .A(n_662), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_663), .A2(n_668), .B1(n_669), .B2(n_672), .Y(n_667) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_671), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_672), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g678 ( .A(n_673), .Y(n_678) );
AOI222xp33_ASAP7_75t_L g717 ( .A1(n_675), .A2(n_718), .B1(n_720), .B2(n_721), .C1(n_725), .C2(n_728), .Y(n_717) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_676), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g751 ( .A(n_676), .B(n_730), .Y(n_751) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_684), .B(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_684), .B(n_744), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B(n_688), .Y(n_685) );
NAND2xp33_ASAP7_75t_SL g689 ( .A(n_690), .B(n_695), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_695), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
NAND4xp25_ASAP7_75t_SL g698 ( .A(n_699), .B(n_717), .C(n_729), .D(n_732), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_704), .B(n_706), .C(n_708), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_705), .A2(n_709), .B1(n_713), .B2(n_715), .Y(n_708) );
INVx1_ASAP7_75t_L g735 ( .A(n_707), .Y(n_735) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_724), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_724), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_741), .A2(n_763), .B1(n_764), .B2(n_765), .Y(n_762) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_745), .B(n_746), .Y(n_742) );
NOR4xp25_ASAP7_75t_L g747 ( .A(n_748), .B(n_753), .C(n_766), .D(n_768), .Y(n_747) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
CKINVDCx11_ASAP7_75t_R g777 ( .A(n_773), .Y(n_777) );
OAI21x1_ASAP7_75t_SL g774 ( .A1(n_775), .A2(n_778), .B(n_779), .Y(n_774) );
BUFx4f_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
INVx3_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
BUFx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx3_ASAP7_75t_L g791 ( .A(n_786), .Y(n_791) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
BUFx3_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_789), .B(n_796), .Y(n_795) );
INVx2_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_791), .B(n_792), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
endmodule