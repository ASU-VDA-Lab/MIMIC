module fake_jpeg_28927_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_8),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_1),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_23),
.Y(n_29)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_24),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_11),
.B1(n_17),
.B2(n_4),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_9),
.C(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_11),
.B1(n_3),
.B2(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_15),
.B1(n_18),
.B2(n_14),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_30),
.A2(n_34),
.B1(n_38),
.B2(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_35),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_27),
.A2(n_18),
.B1(n_19),
.B2(n_14),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_5),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_2),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_45),
.B(n_33),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_36),
.C(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_5),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_35),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_50),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_44),
.C(n_37),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_40),
.B(n_45),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_43),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_54),
.B(n_55),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_49),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_48),
.A3(n_45),
.B1(n_42),
.B2(n_43),
.C1(n_30),
.C2(n_32),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_58),
.B(n_33),
.Y(n_61)
);

AOI222xp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_58),
.B1(n_31),
.B2(n_41),
.C1(n_8),
.C2(n_32),
.Y(n_62)
);


endmodule