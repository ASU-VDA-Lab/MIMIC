module fake_jpeg_17969_n_111 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_111);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_111;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_11),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_13),
.A2(n_19),
.B1(n_23),
.B2(n_12),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_13),
.B1(n_21),
.B2(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_21),
.Y(n_42)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_13),
.B1(n_17),
.B2(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_43),
.B1(n_30),
.B2(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_25),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_72),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_22),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_57),
.B(n_53),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_76),
.A2(n_71),
.B1(n_66),
.B2(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_87),
.B1(n_14),
.B2(n_18),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_59),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_1),
.C(n_2),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_4),
.B(n_6),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_75),
.B1(n_68),
.B2(n_18),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_90),
.A2(n_86),
.B1(n_14),
.B2(n_25),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_22),
.B(n_24),
.Y(n_94)
);

AOI21x1_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_79),
.B(n_81),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_88),
.C(n_93),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_92),
.C(n_90),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_99),
.C(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_4),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_25),
.CI(n_7),
.CON(n_102),
.SN(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

OA21x2_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_97),
.B(n_10),
.Y(n_105)
);

AOI21x1_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_108),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);


endmodule