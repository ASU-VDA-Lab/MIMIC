module fake_jpeg_11842_n_183 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_183);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_13),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_4),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_44),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_81),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_55),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_77),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_0),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_69),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_73),
.B1(n_55),
.B2(n_65),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_99),
.B1(n_100),
.B2(n_63),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_50),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_71),
.B1(n_64),
.B2(n_55),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_71),
.B1(n_68),
.B2(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_53),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_103),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_74),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_106),
.B(n_107),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_46),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_121),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_116),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_66),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_122),
.C(n_24),
.Y(n_133)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_72),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_56),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_48),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_128),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_122),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_143),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_2),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_12),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_7),
.B(n_8),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_7),
.B(n_9),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_148),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_34),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_134),
.B(n_137),
.Y(n_149)
);

AO221x1_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_160),
.B1(n_161),
.B2(n_126),
.C(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NOR4xp25_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_133),
.C(n_130),
.D(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_9),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_10),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_153),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_141),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C1(n_21),
.C2(n_22),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_152),
.C(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_150),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_163),
.B(n_159),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_168),
.B1(n_160),
.B2(n_161),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_165),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_173),
.B(n_169),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_168),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_14),
.B(n_26),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_40),
.Y(n_183)
);


endmodule