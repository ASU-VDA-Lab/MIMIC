module fake_jpeg_31934_n_55 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_55);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_SL g17 ( 
.A1(n_0),
.A2(n_15),
.B(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_25),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx12f_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_38),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_45),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_39),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_46),
.B(n_44),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OAI321xp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_37),
.A3(n_20),
.B1(n_29),
.B2(n_30),
.C(n_41),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_43),
.Y(n_55)
);


endmodule