module fake_jpeg_24386_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_13),
.B(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_43),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_48),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_1),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_56),
.Y(n_94)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_35),
.B1(n_24),
.B2(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_64),
.B1(n_65),
.B2(n_79),
.Y(n_93)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_62),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_35),
.B1(n_24),
.B2(n_28),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_32),
.B1(n_28),
.B2(n_24),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_70),
.B(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_16),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_38),
.A2(n_35),
.B1(n_32),
.B2(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_88),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_32),
.B1(n_20),
.B2(n_44),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_82),
.A2(n_85),
.B1(n_98),
.B2(n_102),
.Y(n_141)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_44),
.B1(n_37),
.B2(n_47),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_36),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_103),
.B1(n_43),
.B2(n_55),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_92),
.B(n_99),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_63),
.B(n_80),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_96),
.A2(n_99),
.A3(n_107),
.B1(n_81),
.B2(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_108),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_29),
.B1(n_16),
.B2(n_23),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_101),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_29),
.B1(n_16),
.B2(n_23),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_29),
.B1(n_40),
.B2(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_105),
.A2(n_34),
.B1(n_30),
.B2(n_21),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_46),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_46),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_113),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_52),
.B(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_41),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_66),
.B(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_128),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_122),
.A2(n_130),
.B(n_140),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_93),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_40),
.C(n_21),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_134),
.B1(n_147),
.B2(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_29),
.B(n_31),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_137),
.B(n_114),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_72),
.C(n_71),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_104),
.C(n_90),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_62),
.B1(n_29),
.B2(n_31),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_136),
.A2(n_25),
.B1(n_91),
.B2(n_83),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_29),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_115),
.B(n_95),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_93),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_103),
.B1(n_110),
.B2(n_87),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_146),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_34),
.B1(n_25),
.B2(n_27),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_3),
.B(n_4),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_175),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_109),
.B(n_113),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_157),
.B(n_160),
.Y(n_198)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_159),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_104),
.B(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_164),
.Y(n_189)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_172),
.C(n_84),
.Y(n_215)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_106),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_169),
.A2(n_22),
.B1(n_18),
.B2(n_4),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_86),
.C(n_89),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_179),
.B1(n_142),
.B2(n_140),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_112),
.B1(n_90),
.B2(n_106),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_174),
.A2(n_119),
.B1(n_132),
.B2(n_130),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_86),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_116),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_22),
.Y(n_204)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_112),
.B1(n_116),
.B2(n_92),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_132),
.B1(n_124),
.B2(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_185),
.A2(n_192),
.B1(n_193),
.B2(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_203),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_149),
.B1(n_138),
.B2(n_119),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_146),
.B1(n_121),
.B2(n_125),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_131),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_196),
.Y(n_219)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_138),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_120),
.B1(n_123),
.B2(n_86),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_120),
.B1(n_123),
.B2(n_27),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_210),
.B1(n_7),
.B2(n_8),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_162),
.B1(n_184),
.B2(n_179),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_22),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_212),
.B(n_5),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_1),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_3),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_167),
.B(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_15),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_3),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_215),
.C(n_216),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_160),
.A2(n_84),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_4),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_84),
.C(n_6),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_150),
.A2(n_174),
.A3(n_157),
.B1(n_153),
.B2(n_158),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_151),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_220),
.A2(n_226),
.B(n_228),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_167),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_235),
.B1(n_210),
.B2(n_200),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_156),
.B(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_187),
.B(n_5),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_6),
.C(n_7),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_243),
.C(n_244),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_190),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_235)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_7),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_202),
.B1(n_217),
.B2(n_214),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_194),
.B(n_8),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_15),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_9),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_9),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_251),
.Y(n_276)
);

AOI311xp33_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_218),
.A3(n_208),
.B(n_192),
.C(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_256),
.Y(n_280)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_257),
.A2(n_258),
.B1(n_269),
.B2(n_11),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_188),
.B1(n_204),
.B2(n_206),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_224),
.C(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_262),
.C(n_224),
.Y(n_271)
);

OA21x2_ASAP7_75t_L g260 ( 
.A1(n_220),
.A2(n_212),
.B(n_207),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_270),
.B(n_232),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_261),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_209),
.C(n_205),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_212),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_233),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_199),
.B1(n_197),
.B2(n_203),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_229),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_282),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_243),
.C(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_275),
.C(n_278),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_229),
.C(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_254),
.C(n_252),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_247),
.B(n_221),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_279),
.B(n_281),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_236),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_246),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_222),
.C(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_264),
.C(n_255),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_222),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_236),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_287),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_242),
.B1(n_235),
.B2(n_13),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_260),
.B(n_250),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_11),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_289),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_288),
.B1(n_272),
.B2(n_247),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_292),
.A2(n_303),
.B1(n_11),
.B2(n_12),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_301),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_251),
.B(n_260),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_275),
.B(n_284),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_248),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_304),
.B(n_263),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_250),
.B1(n_270),
.B2(n_253),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_276),
.A2(n_264),
.B(n_253),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_283),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_249),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_311),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_276),
.B(n_273),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g326 ( 
.A(n_308),
.B(n_310),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_285),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_306),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_313),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_282),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_278),
.B1(n_249),
.B2(n_263),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_296),
.B1(n_295),
.B2(n_298),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_317),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_12),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_301),
.Y(n_328)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_308),
.B1(n_315),
.B2(n_298),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_322),
.A2(n_329),
.B1(n_13),
.B2(n_14),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_305),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_319),
.B(n_291),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_316),
.C(n_294),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_330),
.B(n_331),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_318),
.C(n_14),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_13),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_334),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_14),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_15),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_333),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_321),
.B(n_331),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_339),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_335),
.B(n_337),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_336),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_342),
.B(n_326),
.C(n_327),
.D(n_322),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_330),
.B(n_326),
.Y(n_347)
);


endmodule