module fake_netlist_6_1922_n_782 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_782);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_782;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

BUFx2_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_43),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_36),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_58),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_38),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_57),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_60),
.B(n_143),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_12),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_33),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_22),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_120),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_89),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_92),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_64),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_72),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_135),
.Y(n_174)
);

BUFx2_ASAP7_75t_SL g175 ( 
.A(n_65),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_114),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_91),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_51),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_28),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_11),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_2),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_66),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_100),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_142),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_42),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_L g194 ( 
.A(n_123),
.B(n_93),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_20),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_140),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_133),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_73),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_4),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_59),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_14),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

OAI22x1_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_195),
.B1(n_169),
.B2(n_158),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_145),
.B(n_0),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_1),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_2),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_3),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_3),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_4),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

AOI22x1_ASAP7_75t_SL g226 ( 
.A1(n_186),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_5),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_6),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_15),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_147),
.B(n_7),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_8),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_173),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_152),
.B(n_12),
.Y(n_238)
);

BUFx8_ASAP7_75t_SL g239 ( 
.A(n_163),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_13),
.B(n_16),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_83),
.B(n_17),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_239),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_239),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_215),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_243),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_R g254 ( 
.A(n_242),
.B(n_165),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_243),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_204),
.B(n_156),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_236),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_199),
.B1(n_198),
.B2(n_193),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_204),
.B(n_159),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_160),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_244),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_204),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_241),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_R g283 ( 
.A(n_240),
.B(n_13),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_241),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_212),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_212),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_R g288 ( 
.A(n_240),
.B(n_164),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_223),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_229),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_241),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_241),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_205),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_231),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_233),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_238),
.C(n_232),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_210),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_219),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_247),
.B(n_216),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_230),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_226),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_253),
.B(n_217),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_262),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_295),
.B(n_217),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_265),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_232),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_270),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_264),
.B(n_230),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_238),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_257),
.B(n_218),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_261),
.B(n_216),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

AOI221xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_235),
.B1(n_228),
.B2(n_224),
.C(n_218),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_254),
.B(n_221),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_268),
.B(n_221),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_258),
.B(n_225),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_248),
.B(n_170),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_271),
.B(n_225),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_279),
.B(n_225),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_280),
.B(n_171),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_284),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_225),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_172),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_259),
.B(n_224),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_220),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_285),
.B(n_228),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_288),
.B(n_220),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_286),
.B(n_220),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_249),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_247),
.B(n_222),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_247),
.B(n_222),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_253),
.B(n_222),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_263),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_253),
.B(n_174),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_L g360 ( 
.A(n_253),
.B(n_230),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_304),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_353),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_180),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_230),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_302),
.Y(n_367)
);

OR2x6_ASAP7_75t_L g368 ( 
.A(n_314),
.B(n_245),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_327),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

OR2x6_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_206),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_326),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_355),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_230),
.B1(n_187),
.B2(n_188),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_324),
.B(n_182),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_183),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_296),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_202),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_202),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_327),
.Y(n_384)
);

BUFx12f_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_318),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_337),
.B(n_184),
.Y(n_389)
);

BUFx4f_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_202),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

BUFx8_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_329),
.B(n_202),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_337),
.B(n_206),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_356),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_18),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_19),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_337),
.B(n_21),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_306),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_336),
.B(n_330),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_336),
.B(n_23),
.Y(n_406)
);

OR2x6_ASAP7_75t_L g407 ( 
.A(n_325),
.B(n_24),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_306),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

AO22x1_ASAP7_75t_L g410 ( 
.A1(n_299),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_316),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_315),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

OR2x6_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_29),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_330),
.B(n_30),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_320),
.B(n_32),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_297),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_347),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_300),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_357),
.B(n_34),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_359),
.B(n_35),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_301),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_303),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_322),
.B(n_37),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_298),
.B(n_39),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_350),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_317),
.B(n_40),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_405),
.A2(n_396),
.B(n_381),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_392),
.A2(n_360),
.B(n_334),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_383),
.B(n_322),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_364),
.B(n_346),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_374),
.B(n_340),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_342),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_338),
.Y(n_436)
);

O2A1O1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_365),
.A2(n_425),
.B(n_389),
.C(n_391),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_375),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_SL g439 ( 
.A1(n_401),
.A2(n_308),
.B(n_332),
.C(n_344),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_372),
.B(n_376),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_345),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_339),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_362),
.B(n_309),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_412),
.B(n_390),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_408),
.A2(n_339),
.B1(n_44),
.B2(n_45),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_379),
.A2(n_41),
.B(n_46),
.C(n_47),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_385),
.A2(n_417),
.B1(n_428),
.B2(n_412),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_R g448 ( 
.A(n_363),
.B(n_48),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_390),
.B(n_49),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_399),
.A2(n_50),
.B(n_53),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_367),
.B(n_54),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_369),
.B(n_414),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_R g455 ( 
.A(n_403),
.B(n_55),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_361),
.B(n_62),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_399),
.A2(n_63),
.B(n_67),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_366),
.B(n_68),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_399),
.B(n_69),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_414),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_393),
.B(n_70),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_371),
.B(n_71),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g466 ( 
.A1(n_402),
.A2(n_406),
.B(n_416),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_384),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_407),
.B(n_74),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_373),
.A2(n_75),
.B(n_76),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_409),
.B(n_413),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_373),
.B(n_78),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_422),
.A2(n_377),
.B1(n_421),
.B2(n_368),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_386),
.A2(n_79),
.B(n_80),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_368),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_407),
.B(n_86),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_386),
.B(n_88),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_SL g479 ( 
.A(n_378),
.B(n_90),
.C(n_94),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_388),
.B(n_95),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_400),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_423),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_430),
.A2(n_426),
.B(n_388),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

BUFx4_ASAP7_75t_SL g488 ( 
.A(n_436),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_394),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_443),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_472),
.Y(n_491)
);

INVx8_ASAP7_75t_L g492 ( 
.A(n_454),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_458),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_448),
.Y(n_494)
);

AO21x2_ASAP7_75t_L g495 ( 
.A1(n_466),
.A2(n_382),
.B(n_400),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_454),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_453),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_455),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_440),
.B(n_382),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_429),
.A2(n_395),
.B(n_415),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_435),
.B(n_394),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_442),
.B(n_410),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_470),
.Y(n_504)
);

NAND2x1p5_ASAP7_75t_L g505 ( 
.A(n_461),
.B(n_371),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_431),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_432),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_454),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_477),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_456),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_444),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_433),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_437),
.A2(n_481),
.B(n_452),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_467),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_456),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_484),
.A2(n_415),
.B(n_102),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_457),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_456),
.B(n_101),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_471),
.Y(n_522)
);

OA21x2_ASAP7_75t_L g523 ( 
.A1(n_469),
.A2(n_103),
.B(n_104),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_461),
.B(n_105),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_478),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_474),
.A2(n_473),
.B(n_459),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_497),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_487),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_491),
.A2(n_447),
.B1(n_469),
.B2(n_433),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_492),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_492),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_516),
.A2(n_439),
.B(n_441),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_503),
.A2(n_450),
.B(n_464),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_479),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_493),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_512),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_524),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_530),
.A2(n_446),
.B(n_445),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_509),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_526),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_465),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_517),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_515),
.A2(n_503),
.B1(n_520),
.B2(n_508),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_491),
.A2(n_482),
.B1(n_475),
.B2(n_460),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_486),
.A2(n_451),
.B(n_482),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_504),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_528),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_489),
.Y(n_554)
);

BUFx8_ASAP7_75t_SL g555 ( 
.A(n_490),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_502),
.A2(n_462),
.B1(n_107),
.B2(n_108),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_529),
.B(n_106),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_500),
.Y(n_558)
);

NAND2x1p5_ASAP7_75t_L g559 ( 
.A(n_529),
.B(n_109),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_490),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

CKINVDCx11_ASAP7_75t_R g562 ( 
.A(n_494),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_518),
.Y(n_563)
);

AO21x1_ASAP7_75t_L g564 ( 
.A1(n_501),
.A2(n_110),
.B(n_111),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_115),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_495),
.Y(n_566)
);

CKINVDCx8_ASAP7_75t_R g567 ( 
.A(n_499),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_519),
.A2(n_116),
.B(n_117),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_502),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_489),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_560),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_555),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_552),
.B(n_511),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_535),
.Y(n_574)
);

AOI221xp5_ASAP7_75t_SL g575 ( 
.A1(n_549),
.A2(n_514),
.B1(n_496),
.B2(n_510),
.C(n_513),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_539),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_552),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_565),
.A2(n_523),
.B1(n_521),
.B2(n_529),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_565),
.A2(n_523),
.B1(n_521),
.B2(n_529),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_548),
.B(n_518),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_540),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_514),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_535),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_525),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_561),
.B(n_528),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_538),
.B(n_513),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_531),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_555),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_547),
.B(n_513),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_547),
.B(n_513),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_553),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_538),
.B(n_510),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_541),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_567),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_561),
.B(n_496),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_560),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_510),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_541),
.Y(n_600)
);

OA21x2_ASAP7_75t_L g601 ( 
.A1(n_551),
.A2(n_495),
.B(n_521),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_562),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_554),
.B(n_510),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_563),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_567),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_570),
.B(n_492),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_R g607 ( 
.A(n_543),
.B(n_488),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_563),
.B(n_496),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_533),
.B(n_496),
.Y(n_609)
);

OAI21x1_ASAP7_75t_SL g610 ( 
.A1(n_564),
.A2(n_527),
.B(n_521),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_542),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_557),
.B(n_527),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_545),
.B(n_521),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_R g614 ( 
.A(n_562),
.B(n_488),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_125),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_566),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_566),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_546),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_532),
.B(n_505),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_557),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_583),
.B(n_537),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_617),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_597),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_585),
.B(n_556),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_615),
.A2(n_569),
.B1(n_564),
.B2(n_550),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_616),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_577),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_577),
.B(n_536),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_617),
.B(n_536),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_536),
.Y(n_630)
);

NOR2x1_ASAP7_75t_L g631 ( 
.A(n_596),
.B(n_553),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_581),
.B(n_553),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_580),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_580),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_595),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_595),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_604),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_590),
.B(n_534),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_573),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_599),
.B(n_559),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_618),
.B(n_543),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_600),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_588),
.B(n_543),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_598),
.B(n_559),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_576),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_600),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_597),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_574),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_603),
.B(n_568),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_608),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_594),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_587),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_593),
.B(n_534),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_609),
.B(n_505),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_611),
.B(n_126),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_586),
.B(n_141),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_597),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_601),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_601),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_625),
.A2(n_596),
.B1(n_605),
.B2(n_579),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_645),
.B(n_590),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_645),
.B(n_578),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_639),
.B(n_575),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_621),
.B(n_607),
.C(n_613),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_647),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_652),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_622),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_651),
.B(n_571),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_652),
.Y(n_670)
);

NAND4xp25_ASAP7_75t_L g671 ( 
.A(n_637),
.B(n_606),
.C(n_605),
.D(n_619),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_647),
.B(n_591),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_622),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_633),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_633),
.Y(n_675)
);

AND2x4_ASAP7_75t_SL g676 ( 
.A(n_623),
.B(n_612),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_626),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_653),
.B(n_591),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_650),
.B(n_615),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_650),
.B(n_637),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_632),
.B(n_574),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_630),
.B(n_578),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_640),
.B(n_654),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_626),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_624),
.B(n_620),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_623),
.B(n_612),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_659),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_687),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_683),
.B(n_680),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_685),
.B(n_644),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_681),
.B(n_641),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_687),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_668),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_667),
.B(n_630),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_668),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_682),
.B(n_629),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_669),
.B(n_641),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_673),
.B(n_629),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_643),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_666),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_678),
.B(n_643),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_679),
.B(n_649),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_663),
.B(n_649),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_693),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_694),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_693),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_690),
.A2(n_661),
.B1(n_665),
.B2(n_607),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_R g708 ( 
.A(n_700),
.B(n_623),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_690),
.A2(n_685),
.B1(n_671),
.B2(n_686),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_703),
.A2(n_686),
.B1(n_664),
.B2(n_663),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_697),
.B(n_667),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_695),
.B(n_694),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_688),
.Y(n_713)
);

OAI32xp33_ASAP7_75t_L g714 ( 
.A1(n_698),
.A2(n_657),
.A3(n_655),
.B1(n_675),
.B2(n_674),
.Y(n_714)
);

AOI21xp33_ASAP7_75t_L g715 ( 
.A1(n_707),
.A2(n_657),
.B(n_631),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_L g716 ( 
.A(n_709),
.B(n_602),
.C(n_655),
.Y(n_716)
);

OAI21xp33_ASAP7_75t_L g717 ( 
.A1(n_710),
.A2(n_689),
.B(n_662),
.Y(n_717)
);

OA22x2_ASAP7_75t_L g718 ( 
.A1(n_705),
.A2(n_696),
.B1(n_702),
.B2(n_699),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_711),
.B(n_696),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_708),
.A2(n_686),
.B(n_676),
.Y(n_720)
);

NOR2x1_ASAP7_75t_L g721 ( 
.A(n_720),
.B(n_706),
.Y(n_721)
);

AOI322xp5_ASAP7_75t_L g722 ( 
.A1(n_716),
.A2(n_704),
.A3(n_701),
.B1(n_712),
.B2(n_691),
.C1(n_589),
.C2(n_694),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_719),
.Y(n_723)
);

XOR2x2_ASAP7_75t_L g724 ( 
.A(n_718),
.B(n_589),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_717),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_715),
.B(n_712),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_725),
.B(n_713),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_724),
.A2(n_714),
.B(n_572),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_726),
.B(n_584),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_723),
.B(n_672),
.Y(n_730)
);

AO22x2_ASAP7_75t_L g731 ( 
.A1(n_728),
.A2(n_721),
.B1(n_722),
.B2(n_692),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_727),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_731),
.A2(n_729),
.B(n_730),
.Y(n_733)
);

AOI221xp5_ASAP7_75t_L g734 ( 
.A1(n_732),
.A2(n_614),
.B1(n_672),
.B2(n_662),
.C(n_610),
.Y(n_734)
);

AOI211xp5_ASAP7_75t_L g735 ( 
.A1(n_732),
.A2(n_614),
.B(n_656),
.C(n_574),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_735),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_734),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_733),
.A2(n_662),
.B1(n_672),
.B2(n_676),
.Y(n_738)
);

NOR2x1_ASAP7_75t_L g739 ( 
.A(n_733),
.B(n_584),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_734),
.A2(n_638),
.B1(n_658),
.B2(n_574),
.Y(n_740)
);

NOR2x1_ASAP7_75t_L g741 ( 
.A(n_733),
.B(n_656),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_741),
.A2(n_612),
.B(n_638),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_736),
.B(n_638),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_692),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_739),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_738),
.B(n_688),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_740),
.A2(n_648),
.B1(n_670),
.B2(n_684),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_739),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_748),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_745),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_743),
.Y(n_751)
);

XNOR2xp5_ASAP7_75t_L g752 ( 
.A(n_744),
.B(n_579),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_746),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_747),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_742),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_751),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_749),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_750),
.A2(n_755),
.B1(n_754),
.B2(n_753),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_752),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_751),
.Y(n_761)
);

XOR2x1_ASAP7_75t_L g762 ( 
.A(n_751),
.B(n_129),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_751),
.B(n_670),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_750),
.A2(n_648),
.B1(n_597),
.B2(n_592),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_SL g765 ( 
.A1(n_756),
.A2(n_648),
.B1(n_592),
.B2(n_601),
.Y(n_765)
);

AOI31xp33_ASAP7_75t_L g766 ( 
.A1(n_761),
.A2(n_677),
.A3(n_627),
.B(n_132),
.Y(n_766)
);

OAI31xp33_ASAP7_75t_L g767 ( 
.A1(n_762),
.A2(n_659),
.A3(n_677),
.B(n_627),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_759),
.Y(n_768)
);

OAI31xp33_ASAP7_75t_L g769 ( 
.A1(n_757),
.A2(n_646),
.A3(n_642),
.B(n_636),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_758),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_760),
.B(n_646),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_763),
.B(n_597),
.Y(n_772)
);

AO22x1_ASAP7_75t_L g773 ( 
.A1(n_770),
.A2(n_764),
.B1(n_642),
.B2(n_636),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_768),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_771),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_772),
.Y(n_776)
);

OAI22x1_ASAP7_75t_L g777 ( 
.A1(n_774),
.A2(n_766),
.B1(n_767),
.B2(n_769),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_775),
.A2(n_765),
.B1(n_635),
.B2(n_634),
.C(n_660),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_777),
.B(n_776),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_779),
.A2(n_778),
.B1(n_773),
.B2(n_660),
.Y(n_780)
);

OR2x6_ASAP7_75t_L g781 ( 
.A(n_780),
.B(n_131),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_781),
.A2(n_635),
.B1(n_634),
.B2(n_628),
.Y(n_782)
);


endmodule