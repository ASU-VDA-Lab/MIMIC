module real_aes_9627_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_2043;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_2003;
wire n_1279;
wire n_2014;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_2029;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_2006;
wire n_551;
wire n_884;
wire n_2035;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_2031;
wire n_1160;
wire n_1849;
wire n_2040;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1994;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1583;
wire n_1095;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_1926;
wire n_898;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_2004;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_2038;
wire n_1214;
wire n_806;
wire n_1940;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_2041;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_1945;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_2012;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_2045;
wire n_1401;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_2036;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_2033;
wire n_1769;
wire n_1812;
wire n_1985;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2039;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1580;
wire n_1000;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_2023;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_2019;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_2042;
wire n_1066;
wire n_2046;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1800;
wire n_1435;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_2048;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_2032;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_2027;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_2034;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_2028;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_2011;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_2037;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_2030;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_1969;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_2044;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_2047;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_2010;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_1484;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1003 ( .A1(n_0), .A2(n_711), .B1(n_1004), .B2(n_1006), .C(n_1013), .Y(n_1003) );
AOI21xp33_ASAP7_75t_L g1045 ( .A1(n_0), .A2(n_862), .B(n_1046), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_1), .A2(n_371), .B1(n_770), .B2(n_1041), .Y(n_1391) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1), .Y(n_1414) );
INVx1_ASAP7_75t_L g1424 ( .A(n_2), .Y(n_1424) );
OAI221xp5_ASAP7_75t_L g1453 ( .A1(n_2), .A2(n_209), .B1(n_884), .B2(n_1454), .C(n_1455), .Y(n_1453) );
INVxp67_ASAP7_75t_L g716 ( .A(n_3), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g763 ( .A1(n_3), .A2(n_221), .B1(n_751), .B2(n_764), .C(n_766), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g1243 ( .A(n_4), .Y(n_1243) );
OAI221xp5_ASAP7_75t_L g1288 ( .A1(n_5), .A2(n_547), .B1(n_649), .B2(n_1289), .C(n_1294), .Y(n_1288) );
INVx1_ASAP7_75t_L g1307 ( .A(n_5), .Y(n_1307) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_6), .A2(n_88), .B1(n_493), .B2(n_500), .Y(n_492) );
INVx1_ASAP7_75t_L g537 ( .A(n_6), .Y(n_537) );
INVx1_ASAP7_75t_L g980 ( .A(n_7), .Y(n_980) );
INVxp33_ASAP7_75t_L g1638 ( .A(n_8), .Y(n_1638) );
AOI221xp5_ASAP7_75t_L g1663 ( .A1(n_8), .A2(n_121), .B1(n_1482), .B2(n_1664), .C(n_1665), .Y(n_1663) );
AOI22xp5_ASAP7_75t_L g1722 ( .A1(n_9), .A2(n_360), .B1(n_1708), .B2(n_1711), .Y(n_1722) );
CKINVDCx5p33_ASAP7_75t_R g1938 ( .A(n_10), .Y(n_1938) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_11), .A2(n_275), .B1(n_681), .B2(n_685), .C(n_688), .Y(n_680) );
INVx1_ASAP7_75t_L g757 ( .A(n_11), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g1286 ( .A1(n_12), .A2(n_136), .B1(n_528), .B2(n_529), .C(n_658), .Y(n_1286) );
INVx1_ASAP7_75t_L g1312 ( .A(n_12), .Y(n_1312) );
INVx1_ASAP7_75t_L g1649 ( .A(n_13), .Y(n_1649) );
OAI221xp5_ASAP7_75t_L g1018 ( .A1(n_14), .A2(n_204), .B1(n_701), .B2(n_706), .C(n_708), .Y(n_1018) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_14), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_15), .A2(n_347), .B1(n_1077), .B2(n_1078), .C(n_1080), .Y(n_1076) );
INVx1_ASAP7_75t_L g1090 ( .A(n_15), .Y(n_1090) );
AO22x1_ASAP7_75t_L g1277 ( .A1(n_16), .A2(n_1278), .B1(n_1314), .B2(n_1315), .Y(n_1277) );
INVx1_ASAP7_75t_L g1315 ( .A(n_16), .Y(n_1315) );
AOI22xp33_ASAP7_75t_SL g1185 ( .A1(n_17), .A2(n_337), .B1(n_1130), .B2(n_1131), .Y(n_1185) );
INVxp33_ASAP7_75t_SL g1211 ( .A(n_17), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_18), .Y(n_730) );
INVx1_ASAP7_75t_L g525 ( .A(n_19), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_19), .A2(n_110), .B1(n_592), .B2(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g1061 ( .A(n_20), .Y(n_1061) );
INVxp33_ASAP7_75t_SL g1179 ( .A(n_21), .Y(n_1179) );
AOI221xp5_ASAP7_75t_L g1195 ( .A1(n_21), .A2(n_187), .B1(n_946), .B2(n_952), .C(n_1196), .Y(n_1195) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_22), .Y(n_1332) );
AOI22xp33_ASAP7_75t_SL g1128 ( .A1(n_23), .A2(n_179), .B1(n_832), .B2(n_833), .Y(n_1128) );
AOI221xp5_ASAP7_75t_L g1149 ( .A1(n_23), .A2(n_272), .B1(n_952), .B2(n_1150), .C(n_1152), .Y(n_1149) );
INVx1_ASAP7_75t_L g482 ( .A(n_24), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g546 ( .A1(n_24), .A2(n_547), .B1(n_549), .B2(n_561), .C(n_572), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g698 ( .A1(n_25), .A2(n_143), .B1(n_699), .B2(n_704), .C(n_708), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_25), .A2(n_143), .B1(n_745), .B2(n_748), .Y(n_744) );
OAI221xp5_ASAP7_75t_L g1360 ( .A1(n_26), .A2(n_93), .B1(n_748), .B2(n_1361), .C(n_1362), .Y(n_1360) );
INVx1_ASAP7_75t_L g1365 ( .A(n_26), .Y(n_1365) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_27), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g1723 ( .A1(n_28), .A2(n_312), .B1(n_1701), .B2(n_1719), .Y(n_1723) );
OAI22xp5_ASAP7_75t_L g1220 ( .A1(n_29), .A2(n_350), .B1(n_576), .B2(n_581), .Y(n_1220) );
AOI22xp33_ASAP7_75t_SL g1266 ( .A1(n_29), .A2(n_350), .B1(n_1267), .B2(n_1268), .Y(n_1266) );
AOI221xp5_ASAP7_75t_L g1064 ( .A1(n_30), .A2(n_56), .B1(n_652), .B2(n_977), .C(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_30), .A2(n_314), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
CKINVDCx16_ASAP7_75t_R g1699 ( .A(n_31), .Y(n_1699) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_32), .Y(n_1010) );
INVx1_ASAP7_75t_L g1067 ( .A(n_33), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_33), .A2(n_56), .B1(n_1093), .B2(n_1094), .C(n_1096), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_34), .A2(n_356), .B1(n_827), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g867 ( .A(n_34), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_35), .A2(n_366), .B1(n_621), .B2(n_864), .Y(n_1526) );
INVx1_ASAP7_75t_L g1560 ( .A(n_35), .Y(n_1560) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_36), .A2(n_119), .B1(n_621), .B2(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g659 ( .A(n_36), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_37), .A2(n_89), .B1(n_1021), .B2(n_1023), .Y(n_1020) );
INVx1_ASAP7_75t_L g1043 ( .A(n_37), .Y(n_1043) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_38), .A2(n_68), .B1(n_616), .B2(n_618), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g640 ( .A1(n_38), .A2(n_433), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g1082 ( .A(n_39), .Y(n_1082) );
INVxp33_ASAP7_75t_L g1921 ( .A(n_40), .Y(n_1921) );
AOI221xp5_ASAP7_75t_L g1943 ( .A1(n_40), .A2(n_120), .B1(n_469), .B2(n_1944), .C(n_1945), .Y(n_1943) );
AOI221xp5_ASAP7_75t_L g887 ( .A1(n_41), .A2(n_264), .B1(n_767), .B2(n_875), .C(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g920 ( .A(n_41), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g1928 ( .A1(n_42), .A2(n_194), .B1(n_1929), .B2(n_1930), .Y(n_1928) );
AOI22xp33_ASAP7_75t_L g1952 ( .A1(n_42), .A2(n_194), .B1(n_1953), .B2(n_1954), .Y(n_1952) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_43), .A2(n_50), .B1(n_653), .B2(n_1077), .Y(n_1285) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_43), .A2(n_136), .B1(n_592), .B2(n_595), .Y(n_1313) );
AOI22xp33_ASAP7_75t_SL g1186 ( .A1(n_44), .A2(n_328), .B1(n_832), .B2(n_1187), .Y(n_1186) );
INVxp33_ASAP7_75t_L g1210 ( .A(n_44), .Y(n_1210) );
INVx1_ASAP7_75t_L g381 ( .A(n_45), .Y(n_381) );
INVx1_ASAP7_75t_L g1585 ( .A(n_46), .Y(n_1585) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_46), .A2(n_302), .B1(n_473), .B2(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1628 ( .A(n_47), .Y(n_1628) );
INVx1_ASAP7_75t_L g1518 ( .A(n_48), .Y(n_1518) );
CKINVDCx5p33_ASAP7_75t_R g1669 ( .A(n_49), .Y(n_1669) );
INVx1_ASAP7_75t_L g1311 ( .A(n_50), .Y(n_1311) );
INVx1_ASAP7_75t_L g1575 ( .A(n_51), .Y(n_1575) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_52), .A2(n_142), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_52), .A2(n_234), .B1(n_860), .B2(n_863), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_53), .A2(n_208), .B1(n_469), .B2(n_472), .Y(n_468) );
INVx1_ASAP7_75t_L g571 ( .A(n_53), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g1707 ( .A1(n_54), .A2(n_190), .B1(n_1708), .B2(n_1711), .Y(n_1707) );
AOI22xp33_ASAP7_75t_L g1801 ( .A1(n_55), .A2(n_240), .B1(n_1695), .B2(n_1761), .Y(n_1801) );
INVx1_ASAP7_75t_L g1176 ( .A(n_57), .Y(n_1176) );
CKINVDCx5p33_ASAP7_75t_R g1443 ( .A(n_58), .Y(n_1443) );
AOI22xp33_ASAP7_75t_SL g1932 ( .A1(n_59), .A2(n_333), .B1(n_1130), .B2(n_1933), .Y(n_1932) );
AOI221xp5_ASAP7_75t_L g1949 ( .A1(n_59), .A2(n_333), .B1(n_888), .B2(n_1389), .C(n_1950), .Y(n_1949) );
INVx1_ASAP7_75t_L g836 ( .A(n_60), .Y(n_836) );
CKINVDCx5p33_ASAP7_75t_R g1495 ( .A(n_61), .Y(n_1495) );
INVxp33_ASAP7_75t_L g1578 ( .A(n_62), .Y(n_1578) );
AOI221xp5_ASAP7_75t_L g1608 ( .A1(n_62), .A2(n_320), .B1(n_878), .B2(n_1609), .C(n_1611), .Y(n_1608) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_63), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g1136 ( .A(n_64), .Y(n_1136) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_65), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_66), .A2(n_132), .B1(n_544), .B2(n_661), .Y(n_1287) );
OAI22xp5_ASAP7_75t_SL g1300 ( .A1(n_66), .A2(n_132), .B1(n_495), .B2(n_630), .Y(n_1300) );
XOR2x2_ASAP7_75t_L g1113 ( .A(n_67), .B(n_1114), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g1717 ( .A1(n_67), .A2(n_166), .B1(n_1708), .B2(n_1711), .Y(n_1717) );
INVx1_ASAP7_75t_L g639 ( .A(n_68), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_69), .A2(n_370), .B1(n_769), .B2(n_948), .Y(n_950) );
OAI22xp33_ASAP7_75t_L g989 ( .A1(n_69), .A2(n_353), .B1(n_547), .B2(n_990), .Y(n_989) );
CKINVDCx16_ASAP7_75t_R g1702 ( .A(n_70), .Y(n_1702) );
AO221x2_ASAP7_75t_L g1725 ( .A1(n_71), .A2(n_273), .B1(n_1701), .B2(n_1719), .C(n_1726), .Y(n_1725) );
AOI22xp33_ASAP7_75t_SL g1934 ( .A1(n_72), .A2(n_163), .B1(n_1130), .B2(n_1930), .Y(n_1934) );
INVxp67_ASAP7_75t_SL g1941 ( .A(n_72), .Y(n_1941) );
AOI22xp5_ASAP7_75t_SL g1738 ( .A1(n_73), .A2(n_258), .B1(n_1695), .B2(n_1701), .Y(n_1738) );
INVx1_ASAP7_75t_L g1598 ( .A(n_74), .Y(n_1598) );
INVxp33_ASAP7_75t_L g1627 ( .A(n_75), .Y(n_1627) );
AOI221xp5_ASAP7_75t_L g1655 ( .A1(n_75), .A2(n_150), .B1(n_1656), .B2(n_1658), .C(n_1660), .Y(n_1655) );
CKINVDCx5p33_ASAP7_75t_R g1123 ( .A(n_76), .Y(n_1123) );
INVx1_ASAP7_75t_L g1060 ( .A(n_77), .Y(n_1060) );
INVxp33_ASAP7_75t_SL g1124 ( .A(n_78), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1142 ( .A1(n_78), .A2(n_268), .B1(n_846), .B2(n_1143), .C(n_1145), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_79), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_80), .A2(n_198), .B1(n_433), .B2(n_1012), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_80), .A2(n_198), .B1(n_782), .B2(n_1032), .Y(n_1031) );
INVxp67_ASAP7_75t_SL g1986 ( .A(n_81), .Y(n_1986) );
AOI22xp33_ASAP7_75t_L g2009 ( .A1(n_81), .A2(n_244), .B1(n_830), .B2(n_2010), .Y(n_2009) );
INVxp33_ASAP7_75t_L g1637 ( .A(n_82), .Y(n_1637) );
AOI22xp33_ASAP7_75t_L g1666 ( .A1(n_82), .A2(n_301), .B1(n_613), .B2(n_1667), .Y(n_1666) );
OAI221xp5_ASAP7_75t_L g1632 ( .A1(n_83), .A2(n_257), .B1(n_909), .B2(n_1549), .C(n_1580), .Y(n_1632) );
OAI22xp5_ASAP7_75t_L g1654 ( .A1(n_83), .A2(n_257), .B1(n_748), .B2(n_1607), .Y(n_1654) );
INVx1_ASAP7_75t_L g1596 ( .A(n_84), .Y(n_1596) );
CKINVDCx14_ASAP7_75t_R g1765 ( .A(n_85), .Y(n_1765) );
INVx1_ASAP7_75t_L g1298 ( .A(n_86), .Y(n_1298) );
AOI22xp33_ASAP7_75t_SL g1129 ( .A1(n_87), .A2(n_272), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_87), .A2(n_179), .B1(n_864), .B2(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g542 ( .A(n_88), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_89), .A2(n_152), .B1(n_471), .B2(n_1041), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_90), .A2(n_340), .B1(n_790), .B2(n_1026), .Y(n_1340) );
INVx1_ASAP7_75t_L g1363 ( .A(n_90), .Y(n_1363) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_91), .Y(n_1529) );
INVxp67_ASAP7_75t_SL g1118 ( .A(n_92), .Y(n_1118) );
OAI22xp33_ASAP7_75t_L g1140 ( .A1(n_92), .A2(n_315), .B1(n_841), .B2(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1366 ( .A(n_93), .Y(n_1366) );
XOR2xp5_ASAP7_75t_L g938 ( .A(n_94), .B(n_939), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_95), .Y(n_880) );
INVx1_ASAP7_75t_L g1121 ( .A(n_96), .Y(n_1121) );
INVx1_ASAP7_75t_L g978 ( .A(n_97), .Y(n_978) );
CKINVDCx5p33_ASAP7_75t_R g1394 ( .A(n_98), .Y(n_1394) );
AOI22xp33_ASAP7_75t_SL g1935 ( .A1(n_99), .A2(n_147), .B1(n_1929), .B2(n_1933), .Y(n_1935) );
INVxp67_ASAP7_75t_L g1948 ( .A(n_99), .Y(n_1948) );
INVx1_ASAP7_75t_L g1446 ( .A(n_100), .Y(n_1446) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_100), .A2(n_334), .B1(n_471), .B2(n_614), .Y(n_1456) );
CKINVDCx5p33_ASAP7_75t_R g728 ( .A(n_101), .Y(n_728) );
INVx1_ASAP7_75t_L g1227 ( .A(n_102), .Y(n_1227) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_102), .A2(n_123), .B1(n_878), .B2(n_944), .Y(n_1260) );
AOI22xp33_ASAP7_75t_SL g1427 ( .A1(n_103), .A2(n_205), .B1(n_667), .B2(n_1187), .Y(n_1427) );
AOI22xp33_ASAP7_75t_L g1463 ( .A1(n_103), .A2(n_206), .B1(n_1464), .B2(n_1465), .Y(n_1463) );
INVx1_ASAP7_75t_L g1532 ( .A(n_104), .Y(n_1532) );
OAI221xp5_ASAP7_75t_L g1548 ( .A1(n_104), .A2(n_170), .B1(n_706), .B2(n_1549), .C(n_1550), .Y(n_1548) );
INVx1_ASAP7_75t_L g1541 ( .A(n_105), .Y(n_1541) );
CKINVDCx5p33_ASAP7_75t_R g1603 ( .A(n_106), .Y(n_1603) );
AOI22xp33_ASAP7_75t_L g1799 ( .A1(n_107), .A2(n_230), .B1(n_1708), .B2(n_1800), .Y(n_1799) );
CKINVDCx5p33_ASAP7_75t_R g1537 ( .A(n_108), .Y(n_1537) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_109), .A2(n_332), .B1(n_944), .B2(n_946), .Y(n_943) );
INVx1_ASAP7_75t_L g965 ( .A(n_109), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_110), .A2(n_362), .B1(n_527), .B2(n_529), .C(n_531), .Y(n_526) );
INVx1_ASAP7_75t_L g801 ( .A(n_111), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_111), .A2(n_193), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g486 ( .A(n_112), .Y(n_486) );
OAI211xp5_ASAP7_75t_L g505 ( .A1(n_112), .A2(n_506), .B(n_516), .C(n_536), .Y(n_505) );
INVx1_ASAP7_75t_L g1497 ( .A(n_113), .Y(n_1497) );
AOI221xp5_ASAP7_75t_L g1538 ( .A1(n_114), .A2(n_242), .B1(n_1104), .B2(n_1355), .C(n_1480), .Y(n_1538) );
INVx1_ASAP7_75t_L g1547 ( .A(n_114), .Y(n_1547) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_115), .A2(n_250), .B1(n_488), .B2(n_490), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_115), .A2(n_250), .B1(n_576), .B2(n_581), .Y(n_575) );
INVx1_ASAP7_75t_L g1384 ( .A(n_116), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g1406 ( .A1(n_116), .A2(n_144), .B1(n_705), .B2(n_908), .C(n_909), .Y(n_1406) );
AO22x2_ASAP7_75t_L g1316 ( .A1(n_117), .A2(n_1317), .B1(n_1367), .B2(n_1368), .Y(n_1316) );
CKINVDCx14_ASAP7_75t_R g1367 ( .A(n_117), .Y(n_1367) );
INVx1_ASAP7_75t_L g1600 ( .A(n_118), .Y(n_1600) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_119), .A2(n_125), .B1(n_430), .B2(n_509), .Y(n_666) );
INVxp33_ASAP7_75t_SL g1925 ( .A(n_120), .Y(n_1925) );
INVxp67_ASAP7_75t_L g1641 ( .A(n_121), .Y(n_1641) );
AOI221xp5_ASAP7_75t_L g1479 ( .A1(n_122), .A2(n_265), .B1(n_875), .B2(n_1355), .C(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1504 ( .A(n_122), .Y(n_1504) );
INVx1_ASAP7_75t_L g1225 ( .A(n_123), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_124), .A2(n_139), .B1(n_469), .B2(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g648 ( .A(n_124), .Y(n_648) );
OAI222xp33_ASAP7_75t_L g669 ( .A1(n_125), .A2(n_171), .B1(n_251), .B2(n_597), .C1(n_599), .C2(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g412 ( .A(n_126), .Y(n_412) );
BUFx2_ASAP7_75t_L g427 ( .A(n_126), .Y(n_427) );
INVx1_ASAP7_75t_L g446 ( .A(n_126), .Y(n_446) );
OR2x2_ASAP7_75t_L g703 ( .A(n_126), .B(n_432), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_127), .A2(n_174), .B1(n_433), .B2(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1039 ( .A(n_127), .Y(n_1039) );
CKINVDCx5p33_ASAP7_75t_R g1393 ( .A(n_128), .Y(n_1393) );
INVx1_ASAP7_75t_L g1601 ( .A(n_129), .Y(n_1601) );
INVx1_ASAP7_75t_L g1293 ( .A(n_130), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_130), .A2(n_246), .B1(n_847), .B2(n_945), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_131), .A2(n_135), .B1(n_1437), .B2(n_1439), .Y(n_1436) );
INVx1_ASAP7_75t_L g1467 ( .A(n_131), .Y(n_1467) );
INVx1_ASAP7_75t_L g631 ( .A(n_133), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_133), .A2(n_224), .B1(n_544), .B2(n_661), .C(n_665), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g1133 ( .A1(n_134), .A2(n_227), .B1(n_1130), .B2(n_1131), .Y(n_1133) );
INVxp33_ASAP7_75t_SL g1158 ( .A(n_134), .Y(n_1158) );
INVx1_ASAP7_75t_L g1461 ( .A(n_135), .Y(n_1461) );
INVx1_ASAP7_75t_L g1283 ( .A(n_137), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_137), .A2(n_288), .B1(n_742), .B2(n_847), .Y(n_1309) );
INVx1_ASAP7_75t_L g1577 ( .A(n_138), .Y(n_1577) );
INVx1_ASAP7_75t_L g646 ( .A(n_139), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_140), .Y(n_1246) );
OAI221xp5_ASAP7_75t_L g1579 ( .A1(n_141), .A2(n_357), .B1(n_1549), .B2(n_1580), .C(n_1581), .Y(n_1579) );
OAI22xp5_ASAP7_75t_L g1606 ( .A1(n_141), .A2(n_357), .B1(n_748), .B2(n_1607), .Y(n_1606) );
AOI221xp5_ASAP7_75t_L g855 ( .A1(n_142), .A2(n_297), .B1(n_767), .B2(n_856), .C(n_858), .Y(n_855) );
INVx1_ASAP7_75t_L g1385 ( .A(n_144), .Y(n_1385) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_145), .A2(n_282), .B1(n_832), .B2(n_833), .Y(n_1134) );
INVxp33_ASAP7_75t_L g1157 ( .A(n_145), .Y(n_1157) );
INVx1_ASAP7_75t_L g814 ( .A(n_146), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_146), .A2(n_154), .B1(n_845), .B2(n_846), .C(n_848), .Y(n_844) );
INVxp33_ASAP7_75t_L g1956 ( .A(n_147), .Y(n_1956) );
INVx1_ASAP7_75t_L g1081 ( .A(n_148), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_148), .A2(n_347), .B1(n_1086), .B2(n_1088), .C(n_1089), .Y(n_1085) );
NAND2xp33_ASAP7_75t_SL g1382 ( .A(n_149), .B(n_623), .Y(n_1382) );
INVx1_ASAP7_75t_L g1402 ( .A(n_149), .Y(n_1402) );
INVxp33_ASAP7_75t_L g1631 ( .A(n_150), .Y(n_1631) );
OAI221xp5_ASAP7_75t_L g1234 ( .A1(n_151), .A2(n_506), .B1(n_1235), .B2(n_1240), .C(n_1245), .Y(n_1234) );
AOI22xp33_ASAP7_75t_SL g1264 ( .A1(n_151), .A2(n_237), .B1(n_860), .B2(n_1265), .Y(n_1264) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_152), .A2(n_172), .B1(n_790), .B2(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g793 ( .A(n_153), .Y(n_793) );
INVx1_ASAP7_75t_L g809 ( .A(n_154), .Y(n_809) );
INVx1_ASAP7_75t_L g1924 ( .A(n_155), .Y(n_1924) );
INVx1_ASAP7_75t_L g1178 ( .A(n_156), .Y(n_1178) );
INVx1_ASAP7_75t_L g689 ( .A(n_157), .Y(n_689) );
INVx1_ASAP7_75t_L g406 ( .A(n_158), .Y(n_406) );
INVx1_ASAP7_75t_L g1232 ( .A(n_159), .Y(n_1232) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_159), .A2(n_164), .B1(n_1262), .B2(n_1263), .Y(n_1261) );
INVxp67_ASAP7_75t_L g1590 ( .A(n_160), .Y(n_1590) );
AOI221xp5_ASAP7_75t_L g1613 ( .A1(n_160), .A2(n_228), .B1(n_767), .B2(n_1614), .C(n_1616), .Y(n_1613) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_161), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g1496 ( .A(n_162), .Y(n_1496) );
INVxp33_ASAP7_75t_L g1957 ( .A(n_163), .Y(n_1957) );
INVx1_ASAP7_75t_L g1231 ( .A(n_164), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g2018 ( .A1(n_165), .A2(n_278), .B1(n_1618), .B2(n_1664), .Y(n_2018) );
INVxp67_ASAP7_75t_SL g2022 ( .A(n_165), .Y(n_2022) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_167), .Y(n_895) );
INVx1_ASAP7_75t_L g1471 ( .A(n_168), .Y(n_1471) );
INVx1_ASAP7_75t_L g1991 ( .A(n_169), .Y(n_1991) );
OAI22xp5_ASAP7_75t_L g2026 ( .A1(n_169), .A2(n_321), .B1(n_2027), .B2(n_2029), .Y(n_2026) );
INVx1_ASAP7_75t_L g1531 ( .A(n_170), .Y(n_1531) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_171), .A2(n_293), .B1(n_656), .B2(n_657), .C(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g1048 ( .A(n_172), .Y(n_1048) );
INVxp67_ASAP7_75t_SL g1918 ( .A(n_173), .Y(n_1918) );
OAI22xp33_ASAP7_75t_L g1942 ( .A1(n_173), .A2(n_197), .B1(n_745), .B2(n_748), .Y(n_1942) );
INVx1_ASAP7_75t_L g1035 ( .A(n_174), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1488 ( .A1(n_175), .A2(n_267), .B1(n_1489), .B2(n_1491), .C(n_1492), .Y(n_1488) );
INVx1_ASAP7_75t_L g1513 ( .A(n_175), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g1330 ( .A(n_176), .Y(n_1330) );
AOI22xp5_ASAP7_75t_SL g1737 ( .A1(n_177), .A2(n_195), .B1(n_1708), .B2(n_1711), .Y(n_1737) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_178), .Y(n_890) );
INVx1_ASAP7_75t_L g1685 ( .A(n_180), .Y(n_1685) );
INVx1_ASAP7_75t_L g1325 ( .A(n_181), .Y(n_1325) );
AOI22xp33_ASAP7_75t_SL g1358 ( .A1(n_181), .A2(n_335), .B1(n_847), .B2(n_1207), .Y(n_1358) );
INVxp33_ASAP7_75t_SL g1972 ( .A(n_182), .Y(n_1972) );
AOI22xp33_ASAP7_75t_L g2011 ( .A1(n_182), .A2(n_218), .B1(n_1929), .B2(n_2012), .Y(n_2011) );
CKINVDCx5p33_ASAP7_75t_R g1478 ( .A(n_183), .Y(n_1478) );
INVx1_ASAP7_75t_L g1630 ( .A(n_184), .Y(n_1630) );
AOI22xp33_ASAP7_75t_SL g1184 ( .A1(n_185), .A2(n_225), .B1(n_820), .B2(n_1130), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_185), .A2(n_286), .B1(n_846), .B2(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1445 ( .A(n_186), .Y(n_1445) );
AOI21xp33_ASAP7_75t_L g1457 ( .A1(n_186), .A2(n_1046), .B(n_1458), .Y(n_1457) );
INVxp33_ASAP7_75t_SL g1174 ( .A(n_187), .Y(n_1174) );
CKINVDCx16_ASAP7_75t_R g1692 ( .A(n_188), .Y(n_1692) );
AOI22xp33_ASAP7_75t_L g1962 ( .A1(n_188), .A2(n_1963), .B1(n_1968), .B2(n_2045), .Y(n_1962) );
AO22x2_ASAP7_75t_SL g1968 ( .A1(n_188), .A2(n_1692), .B1(n_1969), .B2(n_2044), .Y(n_1968) );
AOI22xp33_ASAP7_75t_SL g1381 ( .A1(n_189), .A2(n_327), .B1(n_489), .B2(n_490), .Y(n_1381) );
INVx1_ASAP7_75t_L g1401 ( .A(n_189), .Y(n_1401) );
INVx1_ASAP7_75t_L g1686 ( .A(n_191), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1691 ( .A(n_191), .B(n_1684), .Y(n_1691) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_192), .A2(n_222), .B1(n_601), .B2(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g901 ( .A(n_192), .Y(n_901) );
INVx1_ASAP7_75t_L g805 ( .A(n_193), .Y(n_805) );
INVx1_ASAP7_75t_L g1620 ( .A(n_195), .Y(n_1620) );
INVx2_ASAP7_75t_L g393 ( .A(n_196), .Y(n_393) );
INVxp67_ASAP7_75t_SL g1919 ( .A(n_197), .Y(n_1919) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_199), .Y(n_811) );
BUFx3_ASAP7_75t_L g421 ( .A(n_200), .Y(n_421) );
INVx1_ASAP7_75t_L g459 ( .A(n_200), .Y(n_459) );
XNOR2x2_ASAP7_75t_L g677 ( .A(n_201), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g975 ( .A(n_202), .Y(n_975) );
INVxp67_ASAP7_75t_L g723 ( .A(n_203), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_203), .A2(n_281), .B1(n_769), .B2(n_772), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g1053 ( .A(n_204), .Y(n_1053) );
AOI221xp5_ASAP7_75t_L g1462 ( .A1(n_205), .A2(n_304), .B1(n_875), .B2(n_1037), .C(n_1096), .Y(n_1462) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_206), .A2(n_304), .B1(n_1429), .B2(n_1431), .Y(n_1428) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_207), .A2(n_286), .B1(n_832), .B2(n_1183), .Y(n_1182) );
AOI221xp5_ASAP7_75t_L g1201 ( .A1(n_207), .A2(n_225), .B1(n_1093), .B2(n_1202), .C(n_1204), .Y(n_1201) );
INVx1_ASAP7_75t_L g565 ( .A(n_208), .Y(n_565) );
INVx1_ASAP7_75t_L g1423 ( .A(n_209), .Y(n_1423) );
INVx1_ASAP7_75t_L g1320 ( .A(n_210), .Y(n_1320) );
AOI21xp33_ASAP7_75t_L g1359 ( .A1(n_210), .A2(n_742), .B(n_1204), .Y(n_1359) );
CKINVDCx5p33_ASAP7_75t_R g1239 ( .A(n_211), .Y(n_1239) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_212), .A2(n_291), .B1(n_1037), .B2(n_1345), .C(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1409 ( .A(n_212), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g2007 ( .A1(n_213), .A2(n_262), .B1(n_827), .B2(n_2008), .Y(n_2007) );
AOI22xp33_ASAP7_75t_L g2015 ( .A1(n_213), .A2(n_262), .B1(n_1954), .B2(n_2016), .Y(n_2015) );
OAI22xp5_ASAP7_75t_L g1483 ( .A1(n_214), .A2(n_305), .B1(n_882), .B2(n_1484), .Y(n_1483) );
OAI221xp5_ASAP7_75t_L g1506 ( .A1(n_214), .A2(n_305), .B1(n_705), .B2(n_708), .C(n_908), .Y(n_1506) );
INVx1_ASAP7_75t_L g1646 ( .A(n_215), .Y(n_1646) );
INVx1_ASAP7_75t_L g1068 ( .A(n_216), .Y(n_1068) );
AOI22xp33_ASAP7_75t_SL g2006 ( .A1(n_217), .A2(n_364), .B1(n_821), .B2(n_1929), .Y(n_2006) );
AOI22xp33_ASAP7_75t_SL g2017 ( .A1(n_217), .A2(n_364), .B1(n_1345), .B2(n_1667), .Y(n_2017) );
INVx1_ASAP7_75t_L g1989 ( .A(n_218), .Y(n_1989) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_219), .A2(n_353), .B1(n_952), .B2(n_953), .Y(n_951) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_219), .A2(n_370), .B1(n_506), .B2(n_962), .Y(n_961) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_220), .Y(n_959) );
INVxp67_ASAP7_75t_L g719 ( .A(n_221), .Y(n_719) );
INVx1_ASAP7_75t_L g905 ( .A(n_222), .Y(n_905) );
INVx1_ASAP7_75t_L g416 ( .A(n_223), .Y(n_416) );
INVx1_ASAP7_75t_L g453 ( .A(n_223), .Y(n_453) );
INVx1_ASAP7_75t_L g628 ( .A(n_224), .Y(n_628) );
INVx1_ASAP7_75t_L g1922 ( .A(n_226), .Y(n_1922) );
INVxp67_ASAP7_75t_SL g1139 ( .A(n_227), .Y(n_1139) );
INVxp67_ASAP7_75t_L g1588 ( .A(n_228), .Y(n_1588) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_229), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_230), .A2(n_1164), .B1(n_1165), .B2(n_1215), .Y(n_1163) );
INVx1_ASAP7_75t_L g1215 ( .A(n_230), .Y(n_1215) );
CKINVDCx20_ASAP7_75t_R g1376 ( .A(n_231), .Y(n_1376) );
OAI21xp33_ASAP7_75t_L g1057 ( .A1(n_232), .A2(n_1058), .B(n_1083), .Y(n_1057) );
INVx1_ASAP7_75t_L g1112 ( .A(n_232), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_233), .Y(n_1190) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_234), .A2(n_297), .B1(n_825), .B2(n_827), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g1329 ( .A(n_235), .Y(n_1329) );
OA22x2_ASAP7_75t_L g869 ( .A1(n_236), .A2(n_870), .B1(n_930), .B2(n_931), .Y(n_869) );
INVx1_ASAP7_75t_L g931 ( .A(n_236), .Y(n_931) );
OAI221xp5_ASAP7_75t_L g1221 ( .A1(n_237), .A2(n_547), .B1(n_649), .B2(n_1222), .C(n_1228), .Y(n_1221) );
XOR2xp5_ASAP7_75t_L g1000 ( .A(n_238), .B(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1622 ( .A(n_239), .Y(n_1622) );
CKINVDCx14_ASAP7_75t_R g1727 ( .A(n_241), .Y(n_1727) );
INVx1_ASAP7_75t_L g1545 ( .A(n_242), .Y(n_1545) );
XNOR2xp5_ASAP7_75t_L g605 ( .A(n_243), .B(n_606), .Y(n_605) );
INVxp33_ASAP7_75t_SL g1977 ( .A(n_244), .Y(n_1977) );
INVx1_ASAP7_75t_L g1075 ( .A(n_245), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1102 ( .A1(n_245), .A2(n_316), .B1(n_1046), .B2(n_1103), .C(n_1104), .Y(n_1102) );
INVx1_ASAP7_75t_L g1291 ( .A(n_246), .Y(n_1291) );
INVx1_ASAP7_75t_L g521 ( .A(n_247), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_247), .A2(n_362), .B1(n_597), .B2(n_599), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g1524 ( .A(n_248), .Y(n_1524) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_249), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_251), .A2(n_359), .B1(n_652), .B2(n_653), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g1250 ( .A(n_252), .Y(n_1250) );
INVx1_ASAP7_75t_L g1982 ( .A(n_253), .Y(n_1982) );
INVx1_ASAP7_75t_L g1650 ( .A(n_254), .Y(n_1650) );
OAI22xp5_ASAP7_75t_L g1337 ( .A1(n_255), .A2(n_259), .B1(n_1338), .B2(n_1339), .Y(n_1337) );
INVx1_ASAP7_75t_L g1349 ( .A(n_255), .Y(n_1349) );
OA332x1_ASAP7_75t_L g1318 ( .A1(n_256), .A2(n_711), .A3(n_1004), .B1(n_1319), .B2(n_1324), .B3(n_1327), .C1(n_1331), .C2(n_1335), .Y(n_1318) );
AOI21xp5_ASAP7_75t_L g1353 ( .A1(n_256), .A2(n_1354), .B(n_1355), .Y(n_1353) );
AOI22xp33_ASAP7_75t_SL g1352 ( .A1(n_259), .A2(n_340), .B1(n_742), .B2(n_847), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_260), .A2(n_270), .B1(n_769), .B2(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g973 ( .A(n_260), .Y(n_973) );
CKINVDCx5p33_ASAP7_75t_R g1469 ( .A(n_261), .Y(n_1469) );
CKINVDCx5p33_ASAP7_75t_R g1528 ( .A(n_263), .Y(n_1528) );
INVx1_ASAP7_75t_L g916 ( .A(n_264), .Y(n_916) );
INVx1_ASAP7_75t_L g1502 ( .A(n_265), .Y(n_1502) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_266), .A2(n_269), .B1(n_882), .B2(n_884), .Y(n_881) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_266), .A2(n_269), .B1(n_705), .B2(n_908), .C(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g1510 ( .A(n_267), .Y(n_1510) );
INVxp33_ASAP7_75t_SL g1120 ( .A(n_268), .Y(n_1120) );
INVx1_ASAP7_75t_L g971 ( .A(n_270), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_271), .Y(n_1296) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_274), .A2(n_290), .B1(n_616), .B2(n_875), .C(n_876), .Y(n_874) );
INVx1_ASAP7_75t_L g902 ( .A(n_274), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_275), .A2(n_368), .B1(n_751), .B2(n_752), .C(n_754), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_276), .A2(n_306), .B1(n_1041), .B2(n_1464), .Y(n_1493) );
INVx1_ASAP7_75t_L g1514 ( .A(n_276), .Y(n_1514) );
CKINVDCx20_ASAP7_75t_R g1687 ( .A(n_277), .Y(n_1687) );
INVxp33_ASAP7_75t_L g2040 ( .A(n_278), .Y(n_2040) );
BUFx3_ASAP7_75t_L g423 ( .A(n_279), .Y(n_423) );
INVx1_ASAP7_75t_L g461 ( .A(n_279), .Y(n_461) );
AO221x2_ASAP7_75t_L g1760 ( .A1(n_280), .A2(n_352), .B1(n_1761), .B2(n_1762), .C(n_1763), .Y(n_1760) );
INVxp67_ASAP7_75t_L g713 ( .A(n_281), .Y(n_713) );
INVxp67_ASAP7_75t_SL g1148 ( .A(n_282), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1718 ( .A1(n_283), .A2(n_284), .B1(n_1701), .B2(n_1719), .Y(n_1718) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_285), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_285), .B(n_354), .Y(n_432) );
AND2x2_ASAP7_75t_L g510 ( .A(n_285), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g535 ( .A(n_285), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_287), .A2(n_338), .B1(n_945), .B2(n_1104), .C(n_1389), .Y(n_1525) );
INVx1_ASAP7_75t_L g1555 ( .A(n_287), .Y(n_1555) );
INVx1_ASAP7_75t_L g1282 ( .A(n_288), .Y(n_1282) );
CKINVDCx5p33_ASAP7_75t_R g1244 ( .A(n_289), .Y(n_1244) );
INVx1_ASAP7_75t_L g904 ( .A(n_290), .Y(n_904) );
INVx1_ASAP7_75t_L g1415 ( .A(n_291), .Y(n_1415) );
CKINVDCx5p33_ASAP7_75t_R g1295 ( .A(n_292), .Y(n_1295) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_293), .A2(n_359), .B1(n_595), .B2(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g418 ( .A(n_294), .Y(n_418) );
OR2x2_ASAP7_75t_L g594 ( .A(n_294), .B(n_416), .Y(n_594) );
INVx1_ASAP7_75t_L g1565 ( .A(n_295), .Y(n_1565) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_296), .A2(n_313), .B1(n_578), .B2(n_1015), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_296), .A2(n_313), .B1(n_784), .B2(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1008 ( .A(n_298), .Y(n_1008) );
AOI21xp33_ASAP7_75t_L g1036 ( .A1(n_298), .A2(n_767), .B(n_1037), .Y(n_1036) );
CKINVDCx5p33_ASAP7_75t_R g1535 ( .A(n_299), .Y(n_1535) );
AO22x2_ASAP7_75t_L g1216 ( .A1(n_300), .A2(n_1217), .B1(n_1218), .B2(n_1274), .Y(n_1216) );
INVx1_ASAP7_75t_L g1274 ( .A(n_300), .Y(n_1274) );
INVxp67_ASAP7_75t_L g1642 ( .A(n_301), .Y(n_1642) );
INVxp67_ASAP7_75t_L g1593 ( .A(n_302), .Y(n_1593) );
AOI22xp5_ASAP7_75t_SL g1713 ( .A1(n_303), .A2(n_309), .B1(n_1695), .B2(n_1701), .Y(n_1713) );
INVx1_ASAP7_75t_L g1509 ( .A(n_306), .Y(n_1509) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_307), .Y(n_1237) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_308), .A2(n_311), .B1(n_832), .B2(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g854 ( .A(n_308), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g1248 ( .A(n_310), .Y(n_1248) );
INVx1_ASAP7_75t_L g866 ( .A(n_311), .Y(n_866) );
INVxp67_ASAP7_75t_SL g1066 ( .A(n_314), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g1117 ( .A(n_315), .Y(n_1117) );
INVx1_ASAP7_75t_L g1074 ( .A(n_316), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g1911 ( .A1(n_317), .A2(n_1912), .B1(n_1913), .B2(n_1914), .Y(n_1911) );
CKINVDCx5p33_ASAP7_75t_R g1912 ( .A(n_317), .Y(n_1912) );
CKINVDCx5p33_ASAP7_75t_R g1396 ( .A(n_318), .Y(n_1396) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_319), .Y(n_785) );
INVxp33_ASAP7_75t_L g1574 ( .A(n_320), .Y(n_1574) );
INVx1_ASAP7_75t_L g1996 ( .A(n_321), .Y(n_1996) );
INVx1_ASAP7_75t_L g1397 ( .A(n_322), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_323), .A2(n_348), .B1(n_1433), .B2(n_1435), .Y(n_1432) );
INVx1_ASAP7_75t_L g1468 ( .A(n_323), .Y(n_1468) );
INVxp67_ASAP7_75t_SL g1170 ( .A(n_324), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_324), .A2(n_374), .B1(n_841), .B2(n_1141), .Y(n_1194) );
OAI221xp5_ASAP7_75t_SL g1071 ( .A1(n_325), .A2(n_361), .B1(n_644), .B2(n_1072), .C(n_1073), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_325), .A2(n_361), .B1(n_864), .B2(n_945), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_326), .A2(n_351), .B1(n_1465), .B2(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1501 ( .A(n_326), .Y(n_1501) );
INVx1_ASAP7_75t_L g1405 ( .A(n_327), .Y(n_1405) );
INVxp67_ASAP7_75t_SL g1208 ( .A(n_328), .Y(n_1208) );
CKINVDCx5p33_ASAP7_75t_R g1540 ( .A(n_329), .Y(n_1540) );
CKINVDCx5p33_ASAP7_75t_R g1334 ( .A(n_330), .Y(n_1334) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_331), .Y(n_1387) );
INVx1_ASAP7_75t_L g967 ( .A(n_332), .Y(n_967) );
INVx1_ASAP7_75t_L g1441 ( .A(n_334), .Y(n_1441) );
INVx1_ASAP7_75t_L g1321 ( .A(n_335), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g1487 ( .A(n_336), .Y(n_1487) );
INVxp67_ASAP7_75t_SL g1193 ( .A(n_337), .Y(n_1193) );
INVx1_ASAP7_75t_L g1557 ( .A(n_338), .Y(n_1557) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_339), .A2(n_341), .B1(n_489), .B2(n_490), .Y(n_625) );
INVx1_ASAP7_75t_L g634 ( .A(n_339), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_341), .Y(n_635) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_342), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_342), .B(n_381), .Y(n_1682) );
AND3x2_ASAP7_75t_L g1698 ( .A(n_342), .B(n_381), .C(n_1685), .Y(n_1698) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_343), .Y(n_409) );
INVx2_ASAP7_75t_L g394 ( .A(n_344), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_345), .A2(n_363), .B1(n_616), .B2(n_752), .Y(n_889) );
INVx1_ASAP7_75t_L g915 ( .A(n_345), .Y(n_915) );
OAI211xp5_ASAP7_75t_L g1280 ( .A1(n_346), .A2(n_506), .B(n_1281), .C(n_1284), .Y(n_1280) );
INVx1_ASAP7_75t_L g1308 ( .A(n_346), .Y(n_1308) );
INVx1_ASAP7_75t_L g1452 ( .A(n_348), .Y(n_1452) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_349), .Y(n_467) );
INVx1_ASAP7_75t_L g1505 ( .A(n_351), .Y(n_1505) );
INVx1_ASAP7_75t_L g396 ( .A(n_354), .Y(n_396) );
INVx2_ASAP7_75t_L g511 ( .A(n_354), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_355), .Y(n_462) );
INVx1_ASAP7_75t_L g839 ( .A(n_356), .Y(n_839) );
INVx1_ASAP7_75t_L g986 ( .A(n_358), .Y(n_986) );
INVx1_ASAP7_75t_L g922 ( .A(n_363), .Y(n_922) );
AOI21xp33_ASAP7_75t_L g1383 ( .A1(n_365), .A2(n_770), .B(n_1046), .Y(n_1383) );
INVx1_ASAP7_75t_L g1404 ( .A(n_365), .Y(n_1404) );
INVx1_ASAP7_75t_L g1553 ( .A(n_366), .Y(n_1553) );
CKINVDCx5p33_ASAP7_75t_R g1326 ( .A(n_367), .Y(n_1326) );
INVxp33_ASAP7_75t_SL g693 ( .A(n_368), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g2019 ( .A1(n_369), .A2(n_373), .B1(n_952), .B2(n_1041), .Y(n_2019) );
INVxp33_ASAP7_75t_L g2033 ( .A(n_369), .Y(n_2033) );
INVx1_ASAP7_75t_L g1411 ( .A(n_371), .Y(n_1411) );
INVx1_ASAP7_75t_L g1647 ( .A(n_372), .Y(n_1647) );
INVxp67_ASAP7_75t_SL g2037 ( .A(n_373), .Y(n_2037) );
INVxp67_ASAP7_75t_SL g1171 ( .A(n_374), .Y(n_1171) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_397), .B(n_1672), .Y(n_375) );
BUFx12f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1967 ( .A(n_379), .B(n_385), .Y(n_1967) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g1961 ( .A(n_380), .Y(n_1961) );
NAND2xp5_ASAP7_75t_L g2048 ( .A(n_380), .B(n_382), .Y(n_2048) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1960 ( .A(n_382), .B(n_1961), .Y(n_1960) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x6_ASAP7_75t_L g2043 ( .A(n_387), .B(n_412), .Y(n_2043) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g560 ( .A(n_388), .B(n_396), .Y(n_560) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g641 ( .A(n_389), .B(n_642), .Y(n_641) );
INVx8_ASAP7_75t_L g2039 ( .A(n_390), .Y(n_2039) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
INVx2_ASAP7_75t_SL g557 ( .A(n_391), .Y(n_557) );
INVx1_ASAP7_75t_L g715 ( .A(n_391), .Y(n_715) );
OR2x2_ASAP7_75t_L g790 ( .A(n_391), .B(n_703), .Y(n_790) );
BUFx2_ASAP7_75t_L g914 ( .A(n_391), .Y(n_914) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_391), .A2(n_552), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_391), .A2(n_552), .B1(n_1081), .B2(n_1082), .Y(n_1080) );
BUFx6f_ASAP7_75t_L g1328 ( .A(n_391), .Y(n_1328) );
OR2x6_ASAP7_75t_L g2042 ( .A(n_391), .B(n_2032), .Y(n_2042) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g435 ( .A(n_393), .B(n_394), .Y(n_435) );
INVx1_ASAP7_75t_L g514 ( .A(n_393), .Y(n_514) );
INVx2_ASAP7_75t_L g520 ( .A(n_393), .Y(n_520) );
AND2x4_ASAP7_75t_L g524 ( .A(n_393), .B(n_515), .Y(n_524) );
INVx1_ASAP7_75t_L g555 ( .A(n_393), .Y(n_555) );
INVx2_ASAP7_75t_L g515 ( .A(n_394), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_394), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g541 ( .A(n_394), .Y(n_541) );
INVx1_ASAP7_75t_L g554 ( .A(n_394), .Y(n_554) );
INVx1_ASAP7_75t_L g580 ( .A(n_394), .Y(n_580) );
AND2x4_ASAP7_75t_L g2028 ( .A(n_395), .B(n_541), .Y(n_2028) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g2029 ( .A(n_396), .B(n_800), .Y(n_2029) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_1371), .B2(n_1372), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_934), .B2(n_935), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_676), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_602), .B1(n_673), .B2(n_674), .Y(n_402) );
INVx1_ASAP7_75t_L g673 ( .A(n_403), .Y(n_673) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
XNOR2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
AND4x1_ASAP7_75t_L g407 ( .A(n_408), .B(n_436), .C(n_504), .D(n_590), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_410), .B(n_1250), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_410), .B(n_1298), .Y(n_1297) );
OR2x6_ASAP7_75t_L g410 ( .A(n_411), .B(n_424), .Y(n_410) );
INVx2_ASAP7_75t_L g670 ( .A(n_411), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g991 ( .A1(n_411), .A2(n_978), .B1(n_982), .B2(n_986), .C1(n_992), .C2(n_994), .Y(n_991) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
AND2x4_ASAP7_75t_L g478 ( .A(n_412), .B(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g626 ( .A(n_412), .B(n_479), .Y(n_626) );
INVx2_ASAP7_75t_L g1107 ( .A(n_413), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_413), .B(n_1363), .Y(n_1362) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_419), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g444 ( .A(n_414), .B(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g746 ( .A(n_414), .B(n_747), .Y(n_746) );
AND2x2_ASAP7_75t_L g749 ( .A(n_414), .B(n_502), .Y(n_749) );
INVx1_ASAP7_75t_L g778 ( .A(n_414), .Y(n_778) );
AND2x2_ASAP7_75t_L g843 ( .A(n_414), .B(n_502), .Y(n_843) );
AND2x4_ASAP7_75t_L g883 ( .A(n_414), .B(n_747), .Y(n_883) );
AND2x4_ASAP7_75t_L g885 ( .A(n_414), .B(n_502), .Y(n_885) );
BUFx2_ASAP7_75t_L g892 ( .A(n_414), .Y(n_892) );
AND2x4_ASAP7_75t_L g414 ( .A(n_415), .B(n_417), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g479 ( .A(n_417), .B(n_453), .Y(n_479) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g452 ( .A(n_418), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g1975 ( .A(n_418), .Y(n_1975) );
INVx1_ASAP7_75t_L g1980 ( .A(n_418), .Y(n_1980) );
HB1xp67_ASAP7_75t_L g1985 ( .A(n_418), .Y(n_1985) );
INVx6_ASAP7_75t_L g617 ( .A(n_419), .Y(n_617) );
INVx2_ASAP7_75t_L g771 ( .A(n_419), .Y(n_771) );
BUFx2_ASAP7_75t_L g1464 ( .A(n_419), .Y(n_1464) );
AND2x4_ASAP7_75t_L g1983 ( .A(n_419), .B(n_1984), .Y(n_1983) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g503 ( .A(n_420), .Y(n_503) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g442 ( .A(n_421), .B(n_423), .Y(n_442) );
AND2x4_ASAP7_75t_L g471 ( .A(n_421), .B(n_461), .Y(n_471) );
INVx1_ASAP7_75t_L g498 ( .A(n_422), .Y(n_498) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g476 ( .A(n_423), .B(n_459), .Y(n_476) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_425), .A2(n_872), .B1(n_896), .B2(n_897), .Y(n_871) );
INVx2_ASAP7_75t_L g1108 ( .A(n_425), .Y(n_1108) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x6_ASAP7_75t_L g450 ( .A(n_426), .B(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g610 ( .A(n_426), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g818 ( .A(n_426), .B(n_560), .Y(n_818) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_426), .B(n_532), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_426), .B(n_560), .Y(n_1063) );
BUFx2_ASAP7_75t_L g1214 ( .A(n_426), .Y(n_1214) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g589 ( .A(n_427), .Y(n_589) );
OR2x6_ASAP7_75t_L g711 ( .A(n_427), .B(n_641), .Y(n_711) );
INVx1_ASAP7_75t_L g985 ( .A(n_428), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_433), .Y(n_428) );
AND2x2_ASAP7_75t_L g539 ( .A(n_429), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_429), .B(n_540), .Y(n_1247) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x6_ASAP7_75t_L g544 ( .A(n_430), .B(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g572 ( .A(n_430), .B(n_573), .Y(n_572) );
OR2x6_ASAP7_75t_L g649 ( .A(n_430), .B(n_573), .Y(n_649) );
INVx1_ASAP7_75t_L g664 ( .A(n_430), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g987 ( .A1(n_430), .A2(n_638), .B(n_988), .Y(n_987) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_433), .B(n_684), .Y(n_1005) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g667 ( .A(n_434), .Y(n_667) );
INVx2_ASAP7_75t_SL g692 ( .A(n_434), .Y(n_692) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_435), .Y(n_530) );
NOR3xp33_ASAP7_75t_SL g436 ( .A(n_437), .B(n_447), .C(n_492), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_438), .A2(n_494), .B1(n_628), .B2(n_629), .C(n_631), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g956 ( .A1(n_438), .A2(n_629), .B1(n_957), .B2(n_958), .C(n_959), .Y(n_956) );
NOR3xp33_ASAP7_75t_L g1299 ( .A(n_438), .B(n_1300), .C(n_1301), .Y(n_1299) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_443), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g624 ( .A(n_441), .Y(n_624) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_441), .Y(n_779) );
BUFx6f_ASAP7_75t_L g1104 ( .A(n_441), .Y(n_1104) );
AND2x4_ASAP7_75t_L g1999 ( .A(n_441), .B(n_2000), .Y(n_1999) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_442), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_443), .B(n_618), .Y(n_1273) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g499 ( .A(n_444), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_444), .B(n_501), .Y(n_500) );
OR2x6_ASAP7_75t_L g630 ( .A(n_444), .B(n_501), .Y(n_630) );
OR2x6_ASAP7_75t_L g736 ( .A(n_445), .B(n_533), .Y(n_736) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g593 ( .A(n_446), .B(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g684 ( .A(n_446), .B(n_510), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_454), .B1(n_477), .B2(n_480), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g942 ( .A(n_450), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g1259 ( .A(n_450), .Y(n_1259) );
INVx1_ASAP7_75t_L g1390 ( .A(n_451), .Y(n_1390) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g611 ( .A(n_452), .Y(n_611) );
INVx2_ASAP7_75t_SL g767 ( .A(n_452), .Y(n_767) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_452), .Y(n_1097) );
INVx1_ASAP7_75t_L g1204 ( .A(n_452), .Y(n_1204) );
INVx1_ASAP7_75t_L g2003 ( .A(n_453), .Y(n_2003) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_462), .B1(n_463), .B2(n_467), .C(n_468), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g754 ( .A1(n_455), .A2(n_479), .B1(n_689), .B2(n_755), .C(n_757), .Y(n_754) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g598 ( .A(n_456), .Y(n_598) );
INVx2_ASAP7_75t_L g1146 ( .A(n_456), .Y(n_1146) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g481 ( .A(n_457), .Y(n_481) );
OR2x2_ASAP7_75t_L g782 ( .A(n_457), .B(n_594), .Y(n_782) );
INVx1_ASAP7_75t_L g851 ( .A(n_457), .Y(n_851) );
INVx1_ASAP7_75t_L g1087 ( .A(n_457), .Y(n_1087) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
AND2x2_ASAP7_75t_L g466 ( .A(n_458), .B(n_460), .Y(n_466) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_462), .A2(n_467), .B1(n_550), .B2(n_556), .C(n_558), .Y(n_549) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g485 ( .A(n_466), .Y(n_485) );
BUFx2_ASAP7_75t_L g756 ( .A(n_466), .Y(n_756) );
INVx1_ASAP7_75t_L g849 ( .A(n_466), .Y(n_849) );
INVx1_ASAP7_75t_L g1050 ( .A(n_466), .Y(n_1050) );
BUFx4f_ASAP7_75t_L g1304 ( .A(n_466), .Y(n_1304) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g997 ( .A(n_470), .Y(n_997) );
INVx1_ASAP7_75t_L g1093 ( .A(n_470), .Y(n_1093) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
BUFx3_ASAP7_75t_L g489 ( .A(n_471), .Y(n_489) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_471), .Y(n_601) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_471), .Y(n_742) );
BUFx2_ASAP7_75t_L g888 ( .A(n_471), .Y(n_888) );
BUFx6f_ASAP7_75t_L g945 ( .A(n_471), .Y(n_945) );
BUFx6f_ASAP7_75t_L g1037 ( .A(n_471), .Y(n_1037) );
BUFx2_ASAP7_75t_L g1482 ( .A(n_471), .Y(n_1482) );
AND2x6_ASAP7_75t_L g1978 ( .A(n_471), .B(n_1979), .Y(n_1978) );
HB1xp67_ASAP7_75t_L g2016 ( .A(n_471), .Y(n_2016) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g753 ( .A(n_474), .Y(n_753) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g784 ( .A(n_475), .B(n_594), .Y(n_784) );
INVx1_ASAP7_75t_L g1041 ( .A(n_475), .Y(n_1041) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g491 ( .A(n_476), .Y(n_491) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_476), .Y(n_614) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_476), .Y(n_847) );
INVx1_ASAP7_75t_L g1659 ( .A(n_476), .Y(n_1659) );
INVx1_ASAP7_75t_L g955 ( .A(n_477), .Y(n_955) );
OAI22xp5_ASAP7_75t_SL g1301 ( .A1(n_477), .A2(n_610), .B1(n_1302), .B2(n_1306), .Y(n_1301) );
INVx4_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx4f_ASAP7_75t_L g1270 ( .A(n_478), .Y(n_1270) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_479), .Y(n_852) );
INVx1_ASAP7_75t_L g876 ( .A(n_479), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_479), .Y(n_1046) );
INVx2_ASAP7_75t_L g1199 ( .A(n_479), .Y(n_1199) );
INVx2_ASAP7_75t_SL g1355 ( .A(n_479), .Y(n_1355) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B1(n_483), .B2(n_486), .C(n_487), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g1945 ( .A1(n_481), .A2(n_1350), .B1(n_1922), .B2(n_1924), .C(n_1946), .Y(n_1945) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x6_ASAP7_75t_L g595 ( .A(n_485), .B(n_593), .Y(n_595) );
OAI21xp33_ASAP7_75t_L g1034 ( .A1(n_485), .A2(n_1035), .B(n_1036), .Y(n_1034) );
OAI221xp5_ASAP7_75t_L g1145 ( .A1(n_485), .A2(n_852), .B1(n_1121), .B2(n_1123), .C(n_1146), .Y(n_1145) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_488), .Y(n_751) );
BUFx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g946 ( .A(n_490), .Y(n_946) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x6_ASAP7_75t_L g592 ( .A(n_491), .B(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g672 ( .A(n_491), .B(n_593), .Y(n_672) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g958 ( .A(n_495), .Y(n_958) );
INVx2_ASAP7_75t_L g1257 ( .A(n_495), .Y(n_1257) );
NAND2x1p5_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g747 ( .A(n_497), .Y(n_747) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g1995 ( .A(n_498), .Y(n_1995) );
OR2x2_ASAP7_75t_L g1141 ( .A(n_501), .B(n_778), .Y(n_1141) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_502), .A2(n_747), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x6_ASAP7_75t_L g1997 ( .A(n_503), .B(n_1980), .Y(n_1997) );
OAI31xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_546), .A3(n_575), .B(n_585), .Y(n_504) );
INVx8_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AOI221xp5_ASAP7_75t_SL g650 ( .A1(n_507), .A2(n_651), .B1(n_655), .B2(n_659), .C(n_660), .Y(n_650) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
AND2x4_ASAP7_75t_L g582 ( .A(n_508), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g548 ( .A(n_510), .B(n_530), .Y(n_548) );
AND2x2_ASAP7_75t_L g577 ( .A(n_510), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g534 ( .A(n_511), .Y(n_534) );
INVx1_ASAP7_75t_L g642 ( .A(n_511), .Y(n_642) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_512), .Y(n_657) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g528 ( .A(n_513), .Y(n_528) );
BUFx2_ASAP7_75t_L g807 ( .A(n_513), .Y(n_807) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_513), .Y(n_823) );
BUFx6f_ASAP7_75t_L g1012 ( .A(n_513), .Y(n_1012) );
AND2x4_ASAP7_75t_L g2023 ( .A(n_513), .B(n_2024), .Y(n_2023) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OAI221xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_521), .B1(n_522), .B2(n_525), .C(n_526), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g919 ( .A(n_518), .Y(n_919) );
INVx1_ASAP7_75t_L g1007 ( .A(n_518), .Y(n_1007) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g564 ( .A(n_519), .Y(n_564) );
INVx1_ASAP7_75t_L g645 ( .A(n_519), .Y(n_645) );
INVx1_ASAP7_75t_L g545 ( .A(n_520), .Y(n_545) );
AND2x4_ASAP7_75t_L g578 ( .A(n_520), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_SL g820 ( .A(n_522), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g1599 ( .A1(n_522), .A2(n_981), .B1(n_1600), .B2(n_1601), .Y(n_1599) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g830 ( .A(n_523), .Y(n_830) );
INVx2_ASAP7_75t_SL g968 ( .A(n_523), .Y(n_968) );
INVx2_ASAP7_75t_SL g1132 ( .A(n_523), .Y(n_1132) );
INVx2_ASAP7_75t_SL g1226 ( .A(n_523), .Y(n_1226) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g570 ( .A(n_524), .Y(n_570) );
INVx1_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
INVx1_ASAP7_75t_L g2036 ( .A(n_524), .Y(n_2036) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x6_ASAP7_75t_L g687 ( .A(n_528), .B(n_684), .Y(n_687) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_528), .B(n_702), .Y(n_708) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g656 ( .A(n_530), .Y(n_656) );
INVx3_ASAP7_75t_L g826 ( .A(n_530), .Y(n_826) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_SL g658 ( .A(n_532), .Y(n_658) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g2025 ( .A(n_534), .Y(n_2025) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B1(n_542), .B2(n_543), .Y(n_536) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g804 ( .A(n_540), .B(n_702), .Y(n_804) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g663 ( .A(n_541), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_543), .A2(n_1246), .B1(n_1247), .B2(n_1248), .Y(n_1245) );
CKINVDCx11_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g707 ( .A(n_545), .Y(n_707) );
CKINVDCx6p67_ASAP7_75t_R g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g717 ( .A(n_551), .Y(n_717) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx3_ASAP7_75t_L g732 ( .A(n_552), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g979 ( .A1(n_552), .A2(n_980), .B1(n_981), .B2(n_982), .C(n_983), .Y(n_979) );
OAI22xp33_ASAP7_75t_L g1327 ( .A1(n_552), .A2(n_1328), .B1(n_1329), .B2(n_1330), .Y(n_1327) );
BUFx3_ASAP7_75t_L g1639 ( .A(n_552), .Y(n_1639) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g574 ( .A(n_554), .B(n_555), .Y(n_574) );
INVx1_ASAP7_75t_L g800 ( .A(n_555), .Y(n_800) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_556), .A2(n_1229), .B1(n_1231), .B2(n_1232), .C(n_1233), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1294 ( .A1(n_556), .A2(n_638), .B1(n_1233), .B2(n_1295), .C(n_1296), .Y(n_1294) );
OAI22xp33_ASAP7_75t_L g1324 ( .A1(n_556), .A2(n_732), .B1(n_1325), .B2(n_1326), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g1636 ( .A1(n_556), .A2(n_1637), .B1(n_1638), .B2(n_1639), .Y(n_1636) );
OAI22xp33_ASAP7_75t_L g1648 ( .A1(n_556), .A2(n_1639), .B1(n_1649), .B2(n_1650), .Y(n_1648) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_558), .A2(n_970), .B1(n_971), .B2(n_972), .C(n_973), .Y(n_969) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_SL g1233 ( .A(n_560), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B1(n_566), .B2(n_571), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g1290 ( .A(n_564), .Y(n_1290) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g921 ( .A(n_569), .Y(n_921) );
INVx2_ASAP7_75t_L g926 ( .A(n_569), .Y(n_926) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_569), .B(n_684), .Y(n_1027) );
INVx2_ASAP7_75t_L g1079 ( .A(n_569), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1323 ( .A(n_569), .Y(n_1323) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_570), .Y(n_654) );
INVx3_ASAP7_75t_L g697 ( .A(n_570), .Y(n_697) );
INVx1_ASAP7_75t_L g929 ( .A(n_573), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g1517 ( .A1(n_573), .A2(n_912), .B1(n_1487), .B2(n_1495), .Y(n_1517) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g638 ( .A(n_574), .Y(n_638) );
INVx2_ASAP7_75t_L g970 ( .A(n_574), .Y(n_970) );
BUFx2_ASAP7_75t_L g1230 ( .A(n_574), .Y(n_1230) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI221x1_ASAP7_75t_L g633 ( .A1(n_577), .A2(n_582), .B1(n_634), .B2(n_635), .C(n_636), .Y(n_633) );
INVx3_ASAP7_75t_L g990 ( .A(n_577), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g1281 ( .A1(n_577), .A2(n_582), .B1(n_1282), .B2(n_1283), .Y(n_1281) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_578), .Y(n_652) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_578), .Y(n_683) );
BUFx6f_ASAP7_75t_L g1077 ( .A(n_578), .Y(n_1077) );
INVx1_ASAP7_75t_L g1430 ( .A(n_578), .Y(n_1430) );
INVx1_ASAP7_75t_L g1434 ( .A(n_578), .Y(n_1434) );
BUFx2_ASAP7_75t_L g2010 ( .A(n_578), .Y(n_2010) );
AND2x4_ASAP7_75t_L g2031 ( .A(n_578), .B(n_2032), .Y(n_2031) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g962 ( .A(n_582), .Y(n_962) );
INVx1_ASAP7_75t_L g647 ( .A(n_583), .Y(n_647) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g1015 ( .A(n_584), .Y(n_1015) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_586), .A2(n_738), .B1(n_785), .B2(n_786), .Y(n_737) );
INVx5_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g1279 ( .A1(n_587), .A2(n_1280), .B(n_1288), .Y(n_1279) );
BUFx8_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OAI31xp33_ASAP7_75t_L g960 ( .A1(n_588), .A2(n_961), .A3(n_963), .B(n_989), .Y(n_960) );
INVx2_ASAP7_75t_L g1055 ( .A(n_588), .Y(n_1055) );
AOI31xp33_ASAP7_75t_L g1939 ( .A1(n_588), .A2(n_1940), .A3(n_1947), .B(n_1955), .Y(n_1939) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g668 ( .A(n_589), .Y(n_668) );
AND2x4_ASAP7_75t_L g2002 ( .A(n_589), .B(n_2003), .Y(n_2002) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_596), .Y(n_590) );
CKINVDCx6p67_ASAP7_75t_R g994 ( .A(n_592), .Y(n_994) );
OR2x2_ASAP7_75t_L g597 ( .A(n_593), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g599 ( .A(n_593), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g993 ( .A(n_593), .Y(n_993) );
INVx2_ASAP7_75t_L g743 ( .A(n_594), .Y(n_743) );
A2O1A1Ixp33_ASAP7_75t_L g1342 ( .A1(n_594), .A2(n_1343), .B(n_1344), .C(n_1346), .Y(n_1342) );
CKINVDCx6p67_ASAP7_75t_R g998 ( .A(n_595), .Y(n_998) );
INVx1_ASAP7_75t_L g845 ( .A(n_600), .Y(n_845) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g857 ( .A(n_601), .Y(n_857) );
AND2x2_ASAP7_75t_L g879 ( .A(n_601), .B(n_743), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_601), .A2(n_619), .B1(n_1082), .B2(n_1090), .Y(n_1089) );
BUFx4f_ASAP7_75t_L g1491 ( .A(n_601), .Y(n_1491) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g675 ( .A(n_603), .Y(n_675) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR4xp75_ASAP7_75t_L g606 ( .A(n_607), .B(n_632), .C(n_669), .D(n_671), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_627), .Y(n_607) );
AOI33xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .A3(n_615), .B1(n_620), .B2(n_625), .B3(n_626), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_613), .A2(n_1103), .B1(n_1329), .B2(n_1334), .Y(n_1343) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g773 ( .A(n_614), .Y(n_773) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_614), .Y(n_864) );
INVx2_ASAP7_75t_L g954 ( .A(n_614), .Y(n_954) );
INVx1_ASAP7_75t_L g1088 ( .A(n_614), .Y(n_1088) );
AND2x6_ASAP7_75t_L g1987 ( .A(n_614), .B(n_1974), .Y(n_1987) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_617), .Y(n_622) );
INVx2_ASAP7_75t_L g862 ( .A(n_617), .Y(n_862) );
INVx2_ASAP7_75t_L g1103 ( .A(n_617), .Y(n_1103) );
INVx1_ASAP7_75t_L g1207 ( .A(n_617), .Y(n_1207) );
INVx2_ASAP7_75t_SL g1458 ( .A(n_617), .Y(n_1458) );
INVx2_ASAP7_75t_L g1976 ( .A(n_617), .Y(n_1976) );
BUFx2_ASAP7_75t_SL g858 ( .A(n_618), .Y(n_858) );
INVx1_ASAP7_75t_L g1151 ( .A(n_618), .Y(n_1151) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g762 ( .A(n_619), .B(n_743), .Y(n_762) );
AND2x4_ASAP7_75t_L g891 ( .A(n_619), .B(n_892), .Y(n_891) );
INVx2_ASAP7_75t_SL g1095 ( .A(n_619), .Y(n_1095) );
INVx1_ASAP7_75t_L g1203 ( .A(n_619), .Y(n_1203) );
BUFx3_ASAP7_75t_L g1265 ( .A(n_619), .Y(n_1265) );
BUFx4f_ASAP7_75t_L g1345 ( .A(n_619), .Y(n_1345) );
INVx1_ASAP7_75t_L g1490 ( .A(n_619), .Y(n_1490) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g1480 ( .A(n_622), .Y(n_1480) );
INVx4_ASAP7_75t_L g1667 ( .A(n_622), .Y(n_1667) );
INVx1_ASAP7_75t_L g765 ( .A(n_623), .Y(n_765) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g875 ( .A(n_624), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g1256 ( .A1(n_629), .A2(n_1246), .B1(n_1248), .B2(n_1257), .Y(n_1256) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI21x1_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_650), .B(n_668), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_643), .B(n_649), .Y(n_636) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g1587 ( .A(n_638), .Y(n_1587) );
BUFx2_ASAP7_75t_L g1597 ( .A(n_638), .Y(n_1597) );
INVx1_ASAP7_75t_L g2032 ( .A(n_642), .Y(n_2032) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_643) );
INVx2_ASAP7_75t_L g1224 ( .A(n_644), .Y(n_1224) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx3_ASAP7_75t_L g722 ( .A(n_645), .Y(n_722) );
HB1xp67_ASAP7_75t_L g1592 ( .A(n_653), .Y(n_1592) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g977 ( .A(n_654), .Y(n_977) );
INVx3_ASAP7_75t_L g1644 ( .A(n_654), .Y(n_1644) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_657), .Y(n_1183) );
AOI211xp5_ASAP7_75t_L g2021 ( .A1(n_657), .A2(n_2022), .B(n_2023), .C(n_2026), .Y(n_2021) );
INVx1_ASAP7_75t_L g983 ( .A(n_658), .Y(n_983) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
NAND2x1_ASAP7_75t_SL g701 ( .A(n_662), .B(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_662), .A2(n_707), .B1(n_957), .B2(n_959), .Y(n_988) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
BUFx3_ASAP7_75t_L g1929 ( .A(n_667), .Y(n_1929) );
INVx2_ASAP7_75t_L g868 ( .A(n_668), .Y(n_868) );
OAI31xp33_ASAP7_75t_L g1341 ( .A1(n_668), .A2(n_1342), .A3(n_1347), .B(n_1360), .Y(n_1341) );
AOI22xp5_ASAP7_75t_L g1651 ( .A1(n_668), .A2(n_788), .B1(n_1652), .B2(n_1669), .Y(n_1651) );
AND2x4_ASAP7_75t_L g789 ( .A(n_670), .B(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
XNOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_791), .Y(n_676) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_737), .Y(n_678) );
NOR3xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_698), .C(n_709), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_682), .A2(n_691), .B1(n_1445), .B2(n_1446), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1920 ( .A1(n_682), .A2(n_686), .B1(n_1921), .B2(n_1922), .Y(n_1920) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
AND2x2_ASAP7_75t_L g815 ( .A(n_683), .B(n_684), .Y(n_815) );
INVx2_ASAP7_75t_SL g828 ( .A(n_683), .Y(n_828) );
AND2x2_ASAP7_75t_L g906 ( .A(n_683), .B(n_684), .Y(n_906) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_683), .B(n_684), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_683), .B(n_684), .Y(n_1180) );
AND2x4_ASAP7_75t_L g691 ( .A(n_684), .B(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g696 ( .A(n_684), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_684), .B(n_823), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_684), .A2(n_1017), .B1(n_1071), .B2(n_1076), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_687), .A2(n_809), .B1(n_810), .B2(n_811), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_687), .A2(n_696), .B1(n_901), .B2(n_902), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_687), .A2(n_810), .B1(n_1120), .B2(n_1121), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_687), .A2(n_1174), .B1(n_1175), .B2(n_1176), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_687), .A2(n_695), .B1(n_1401), .B2(n_1402), .Y(n_1400) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_687), .A2(n_1441), .B1(n_1442), .B2(n_1443), .Y(n_1440) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_687), .A2(n_696), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1544 ( .A1(n_687), .A2(n_810), .B1(n_1537), .B2(n_1545), .Y(n_1544) );
AOI22xp33_ASAP7_75t_L g1573 ( .A1(n_687), .A2(n_1175), .B1(n_1574), .B2(n_1575), .Y(n_1573) );
AOI22xp33_ASAP7_75t_L g1626 ( .A1(n_687), .A2(n_695), .B1(n_1627), .B2(n_1628), .Y(n_1626) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_693), .B2(n_694), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g1923 ( .A1(n_690), .A2(n_1924), .B1(n_1925), .B2(n_1926), .Y(n_1923) );
BUFx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_691), .A2(n_813), .B1(n_814), .B2(n_815), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_691), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_691), .A2(n_906), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_691), .A2(n_1178), .B1(n_1179), .B2(n_1180), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_691), .A2(n_1022), .B1(n_1404), .B2(n_1405), .Y(n_1403) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_691), .A2(n_906), .B1(n_1504), .B2(n_1505), .Y(n_1503) );
AOI22xp33_ASAP7_75t_L g1546 ( .A1(n_691), .A2(n_1180), .B1(n_1535), .B2(n_1547), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1576 ( .A1(n_691), .A2(n_1180), .B1(n_1577), .B2(n_1578), .Y(n_1576) );
AOI22xp33_ASAP7_75t_L g1629 ( .A1(n_691), .A2(n_1180), .B1(n_1630), .B2(n_1631), .Y(n_1629) );
BUFx3_ASAP7_75t_L g832 ( .A(n_692), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_692), .A2(n_807), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
INVx1_ASAP7_75t_L g1438 ( .A(n_692), .Y(n_1438) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx2_ASAP7_75t_L g810 ( .A(n_696), .Y(n_810) );
BUFx2_ASAP7_75t_L g1175 ( .A(n_696), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1442 ( .A(n_696), .Y(n_1442) );
BUFx2_ASAP7_75t_L g1926 ( .A(n_696), .Y(n_1926) );
BUFx3_ASAP7_75t_L g725 ( .A(n_697), .Y(n_725) );
INVx1_ASAP7_75t_SL g1009 ( .A(n_697), .Y(n_1009) );
INVx2_ASAP7_75t_L g1072 ( .A(n_697), .Y(n_1072) );
INVx1_ASAP7_75t_L g1292 ( .A(n_697), .Y(n_1292) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g1549 ( .A(n_700), .Y(n_1549) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_701), .Y(n_908) );
NAND2x1p5_ASAP7_75t_L g706 ( .A(n_702), .B(n_707), .Y(n_706) );
AND2x4_ASAP7_75t_L g798 ( .A(n_702), .B(n_799), .Y(n_798) );
AND2x4_ASAP7_75t_L g806 ( .A(n_702), .B(n_807), .Y(n_806) );
INVx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx4f_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
BUFx4f_ASAP7_75t_L g1580 ( .A(n_706), .Y(n_1580) );
BUFx3_ASAP7_75t_L g909 ( .A(n_708), .Y(n_909) );
BUFx2_ASAP7_75t_L g1550 ( .A(n_708), .Y(n_1550) );
BUFx2_ASAP7_75t_L g1581 ( .A(n_708), .Y(n_1581) );
OAI33xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .A3(n_718), .B1(n_726), .B2(n_729), .B3(n_734), .Y(n_709) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI33xp33_ASAP7_75t_L g910 ( .A1(n_711), .A2(n_734), .A3(n_911), .B1(n_917), .B2(n_923), .B3(n_927), .Y(n_910) );
OAI33xp33_ASAP7_75t_L g1407 ( .A1(n_711), .A2(n_734), .A3(n_1408), .B1(n_1412), .B2(n_1416), .B3(n_1417), .Y(n_1407) );
OAI33xp33_ASAP7_75t_L g1507 ( .A1(n_711), .A2(n_736), .A3(n_1508), .B1(n_1511), .B2(n_1515), .B3(n_1517), .Y(n_1507) );
OAI33xp33_ASAP7_75t_L g1551 ( .A1(n_711), .A2(n_734), .A3(n_1552), .B1(n_1556), .B2(n_1561), .B3(n_1562), .Y(n_1551) );
OAI33xp33_ASAP7_75t_L g1582 ( .A1(n_711), .A2(n_734), .A3(n_1583), .B1(n_1589), .B2(n_1594), .B3(n_1599), .Y(n_1582) );
INVx1_ASAP7_75t_L g1635 ( .A(n_711), .Y(n_1635) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_714), .B1(n_716), .B2(n_717), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_714), .A2(n_720), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g981 ( .A(n_715), .Y(n_981) );
INVx1_ASAP7_75t_L g1238 ( .A(n_715), .Y(n_1238) );
OAI22xp33_ASAP7_75t_L g1508 ( .A1(n_717), .A2(n_912), .B1(n_1509), .B2(n_1510), .Y(n_1508) );
OAI22xp33_ASAP7_75t_L g1562 ( .A1(n_717), .A2(n_1524), .B1(n_1528), .B2(n_1563), .Y(n_1562) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_723), .B2(n_724), .Y(n_718) );
BUFx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_721), .A2(n_975), .B1(n_976), .B2(n_978), .Y(n_974) );
INVx2_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g966 ( .A(n_722), .Y(n_966) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_724), .A2(n_730), .B1(n_731), .B2(n_733), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g1645 ( .A1(n_724), .A2(n_1241), .B1(n_1646), .B2(n_1647), .Y(n_1645) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g1418 ( .A(n_725), .Y(n_1418) );
CKINVDCx5p33_ASAP7_75t_R g1931 ( .A(n_725), .Y(n_1931) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_727), .A2(n_730), .B1(n_781), .B2(n_783), .Y(n_780) );
AOI211xp5_ASAP7_75t_L g739 ( .A1(n_728), .A2(n_740), .B(n_744), .C(n_750), .Y(n_739) );
BUFx3_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_732), .A2(n_912), .B1(n_915), .B2(n_916), .Y(n_911) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_732), .A2(n_1413), .B1(n_1414), .B2(n_1415), .Y(n_1412) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_733), .A2(n_759), .B1(n_763), .B2(n_768), .C(n_774), .Y(n_758) );
OAI33xp33_ASAP7_75t_L g1633 ( .A1(n_734), .A2(n_1634), .A3(n_1636), .B1(n_1640), .B2(n_1645), .B3(n_1648), .Y(n_1633) );
INVx1_ASAP7_75t_L g1936 ( .A(n_734), .Y(n_1936) );
CKINVDCx8_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
INVx5_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx6_ASAP7_75t_L g834 ( .A(n_736), .Y(n_834) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_758), .C(n_780), .Y(n_738) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI211xp5_ASAP7_75t_SL g838 ( .A1(n_741), .A2(n_839), .B(n_840), .C(n_844), .Y(n_838) );
AOI211xp5_ASAP7_75t_L g1138 ( .A1(n_741), .A2(n_1139), .B(n_1140), .C(n_1142), .Y(n_1138) );
AOI211xp5_ASAP7_75t_L g1192 ( .A1(n_741), .A2(n_1193), .B(n_1194), .C(n_1195), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1395 ( .A(n_741), .B(n_1396), .Y(n_1395) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_741), .A2(n_1478), .B1(n_1479), .B2(n_1481), .C(n_1483), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_741), .B(n_1540), .Y(n_1539) );
AOI211xp5_ASAP7_75t_L g1605 ( .A1(n_741), .A2(n_1596), .B(n_1606), .C(n_1608), .Y(n_1605) );
AOI22xp33_ASAP7_75t_L g1668 ( .A1(n_741), .A2(n_781), .B1(n_1646), .B2(n_1649), .Y(n_1668) );
AOI211xp5_ASAP7_75t_L g1940 ( .A1(n_741), .A2(n_1941), .B(n_1942), .C(n_1943), .Y(n_1940) );
AND2x4_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
BUFx3_ASAP7_75t_L g1267 ( .A(n_742), .Y(n_1267) );
INVx2_ASAP7_75t_SL g1615 ( .A(n_742), .Y(n_1615) );
AOI222xp33_ASAP7_75t_L g1084 ( .A1(n_743), .A2(n_883), .B1(n_885), .B2(n_1060), .C1(n_1061), .C2(n_1085), .Y(n_1084) );
INVx2_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g841 ( .A(n_746), .Y(n_841) );
INVx2_ASAP7_75t_SL g1361 ( .A(n_746), .Y(n_1361) );
AOI322xp5_ASAP7_75t_L g1380 ( .A1(n_746), .A2(n_885), .A3(n_1381), .B1(n_1382), .B2(n_1383), .C1(n_1384), .C2(n_1385), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_746), .A2(n_843), .B1(n_1531), .B2(n_1532), .Y(n_1530) );
INVx1_ASAP7_75t_L g1607 ( .A(n_746), .Y(n_1607) );
INVx3_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g1465 ( .A(n_753), .Y(n_1465) );
INVx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g1197 ( .A(n_756), .Y(n_1197) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_761), .A2(n_776), .B1(n_854), .B2(n_855), .C(n_859), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g1147 ( .A1(n_761), .A2(n_776), .B1(n_1148), .B2(n_1149), .C(n_1154), .Y(n_1147) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_761), .A2(n_776), .B1(n_1201), .B2(n_1205), .C(n_1208), .Y(n_1200) );
AOI221xp5_ASAP7_75t_L g1612 ( .A1(n_761), .A2(n_776), .B1(n_1598), .B2(n_1613), .C(n_1617), .Y(n_1612) );
AOI221xp5_ASAP7_75t_L g1662 ( .A1(n_761), .A2(n_776), .B1(n_1650), .B2(n_1663), .C(n_1666), .Y(n_1662) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g886 ( .A1(n_762), .A2(n_887), .B1(n_889), .B2(n_890), .C(n_891), .Y(n_886) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_762), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g1386 ( .A1(n_762), .A2(n_891), .B1(n_1387), .B2(n_1388), .C(n_1391), .Y(n_1386) );
HB1xp67_ASAP7_75t_L g1460 ( .A(n_762), .Y(n_1460) );
HB1xp67_ASAP7_75t_L g1486 ( .A(n_762), .Y(n_1486) );
AOI221xp5_ASAP7_75t_L g1523 ( .A1(n_762), .A2(n_891), .B1(n_1524), .B2(n_1525), .C(n_1526), .Y(n_1523) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
BUFx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g1153 ( .A(n_767), .Y(n_1153) );
BUFx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g992 ( .A(n_770), .B(n_993), .Y(n_992) );
A2O1A1Ixp33_ASAP7_75t_L g1047 ( .A1(n_770), .A2(n_1048), .B(n_1049), .C(n_1054), .Y(n_1047) );
INVx2_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g1155 ( .A(n_771), .Y(n_1155) );
INVx1_ASAP7_75t_L g1354 ( .A(n_771), .Y(n_1354) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g1947 ( .A1(n_776), .A2(n_1486), .B1(n_1948), .B2(n_1949), .C(n_1952), .Y(n_1947) );
AND2x4_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g949 ( .A(n_779), .Y(n_949) );
BUFx6f_ASAP7_75t_L g1664 ( .A(n_779), .Y(n_1664) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_781), .A2(n_783), .B1(n_866), .B2(n_867), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_781), .A2(n_783), .B1(n_894), .B2(n_895), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_781), .A2(n_783), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_781), .A2(n_783), .B1(n_1210), .B2(n_1211), .Y(n_1209) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_781), .A2(n_783), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_781), .A2(n_783), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
AOI22xp33_ASAP7_75t_L g1494 ( .A1(n_781), .A2(n_783), .B1(n_1495), .B2(n_1496), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_781), .A2(n_783), .B1(n_1528), .B2(n_1529), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g1619 ( .A1(n_781), .A2(n_783), .B1(n_1600), .B2(n_1601), .Y(n_1619) );
AOI22xp33_ASAP7_75t_L g1955 ( .A1(n_781), .A2(n_783), .B1(n_1956), .B2(n_1957), .Y(n_1955) );
INVx6_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI211xp5_ASAP7_75t_L g1653 ( .A1(n_783), .A2(n_1647), .B(n_1654), .C(n_1655), .Y(n_1653) );
INVx4_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_788), .A2(n_836), .B(n_837), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g1135 ( .A1(n_788), .A2(n_1136), .B(n_1137), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_788), .A2(n_1448), .B1(n_1522), .B2(n_1541), .Y(n_1521) );
AOI21xp33_ASAP7_75t_SL g1602 ( .A1(n_788), .A2(n_1603), .B(n_1604), .Y(n_1602) );
INVx5_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_SL g897 ( .A(n_789), .Y(n_897) );
INVx1_ASAP7_75t_L g1189 ( .A(n_789), .Y(n_1189) );
INVx2_ASAP7_75t_L g1470 ( .A(n_789), .Y(n_1470) );
INVx2_ASAP7_75t_L g1069 ( .A(n_790), .Y(n_1069) );
AO22x2_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_869), .B1(n_932), .B2(n_933), .Y(n_791) );
INVx1_ASAP7_75t_L g933 ( .A(n_792), .Y(n_933) );
XNOR2x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
AND2x4_ASAP7_75t_L g794 ( .A(n_795), .B(n_835), .Y(n_794) );
AND4x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_808), .C(n_812), .D(n_816), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_801), .B1(n_802), .B2(n_805), .C(n_806), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g1116 ( .A1(n_797), .A2(n_802), .B1(n_806), .B2(n_1117), .C(n_1118), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_798), .A2(n_804), .B1(n_806), .B2(n_1060), .C(n_1061), .Y(n_1059) );
INVx1_ASAP7_75t_L g1169 ( .A(n_798), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1364 ( .A1(n_798), .A2(n_804), .B1(n_806), .B2(n_1365), .C(n_1366), .Y(n_1364) );
AOI221xp5_ASAP7_75t_L g1422 ( .A1(n_798), .A2(n_804), .B1(n_806), .B2(n_1423), .C(n_1424), .Y(n_1422) );
AOI221xp5_ASAP7_75t_L g1917 ( .A1(n_798), .A2(n_804), .B1(n_806), .B2(n_1918), .C(n_1919), .Y(n_1917) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g1167 ( .A1(n_804), .A2(n_1168), .B1(n_1170), .B2(n_1171), .C(n_1172), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_806), .Y(n_1172) );
HB1xp67_ASAP7_75t_L g1933 ( .A(n_807), .Y(n_1933) );
INVx1_ASAP7_75t_L g2013 ( .A(n_807), .Y(n_2013) );
OAI221xp5_ASAP7_75t_L g848 ( .A1(n_811), .A2(n_813), .B1(n_849), .B2(n_850), .C(n_852), .Y(n_848) );
AOI33xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_819), .A3(n_824), .B1(n_829), .B2(n_831), .B3(n_834), .Y(n_816) );
BUFx3_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g1127 ( .A(n_818), .Y(n_1127) );
INVx2_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g833 ( .A(n_822), .Y(n_833) );
INVx2_ASAP7_75t_SL g822 ( .A(n_823), .Y(n_822) );
BUFx6f_ASAP7_75t_L g1187 ( .A(n_823), .Y(n_1187) );
INVx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AOI33xp33_ASAP7_75t_L g1125 ( .A1(n_834), .A2(n_1126), .A3(n_1128), .B1(n_1129), .B2(n_1133), .B3(n_1134), .Y(n_1125) );
AOI33xp33_ASAP7_75t_L g1181 ( .A1(n_834), .A2(n_1126), .A3(n_1182), .B1(n_1184), .B2(n_1185), .B3(n_1186), .Y(n_1181) );
INVx1_ASAP7_75t_L g1335 ( .A(n_834), .Y(n_1335) );
AOI33xp33_ASAP7_75t_L g1425 ( .A1(n_834), .A2(n_1426), .A3(n_1427), .B1(n_1428), .B2(n_1432), .B3(n_1436), .Y(n_1425) );
AOI33xp33_ASAP7_75t_L g2005 ( .A1(n_834), .A2(n_1126), .A3(n_2006), .B1(n_2007), .B2(n_2009), .B3(n_2011), .Y(n_2005) );
AOI31xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_853), .A3(n_865), .B(n_868), .Y(n_837) );
INVx2_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
BUFx3_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_847), .Y(n_878) );
INVx1_ASAP7_75t_L g1269 ( .A(n_847), .Y(n_1269) );
OAI211xp5_ASAP7_75t_L g1042 ( .A1(n_849), .A2(n_1043), .B(n_1044), .C(n_1045), .Y(n_1042) );
OAI211xp5_ASAP7_75t_L g1455 ( .A1(n_849), .A2(n_1443), .B(n_1456), .C(n_1457), .Y(n_1455) );
OAI221xp5_ASAP7_75t_L g1611 ( .A1(n_849), .A2(n_852), .B1(n_1146), .B2(n_1575), .C(n_1577), .Y(n_1611) );
OAI221xp5_ASAP7_75t_L g1660 ( .A1(n_849), .A2(n_1146), .B1(n_1628), .B2(n_1630), .C(n_1661), .Y(n_1660) );
OAI22xp5_ASAP7_75t_L g1038 ( .A1(n_850), .A2(n_1010), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
OAI221xp5_ASAP7_75t_L g1196 ( .A1(n_850), .A2(n_1176), .B1(n_1178), .B2(n_1197), .C(n_1198), .Y(n_1196) );
OAI221xp5_ASAP7_75t_L g1306 ( .A1(n_850), .A2(n_1303), .B1(n_1307), .B2(n_1308), .C(n_1309), .Y(n_1306) );
INVx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
BUFx6f_ASAP7_75t_L g1099 ( .A(n_862), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g1536 ( .A(n_864), .Y(n_1536) );
AOI31xp33_ASAP7_75t_L g1137 ( .A1(n_868), .A2(n_1138), .A3(n_1147), .B(n_1156), .Y(n_1137) );
INVx1_ASAP7_75t_L g1448 ( .A(n_868), .Y(n_1448) );
AOI31xp33_ASAP7_75t_L g1604 ( .A1(n_868), .A2(n_1605), .A3(n_1612), .B(n_1619), .Y(n_1604) );
INVx3_ASAP7_75t_L g932 ( .A(n_869), .Y(n_932) );
INVx1_ASAP7_75t_L g930 ( .A(n_870), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_898), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g872 ( .A(n_873), .B(n_886), .C(n_893), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_877), .B1(n_879), .B2(n_880), .C(n_881), .Y(n_873) );
INVx1_ASAP7_75t_L g1951 ( .A(n_875), .Y(n_1951) );
INVx1_ASAP7_75t_L g1946 ( .A(n_876), .Y(n_1946) );
INVx1_ASAP7_75t_L g1030 ( .A(n_879), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_880), .A2(n_895), .B1(n_918), .B2(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx4_ASAP7_75t_L g1454 ( .A(n_883), .Y(n_1454) );
INVx2_ASAP7_75t_SL g884 ( .A(n_885), .Y(n_884) );
INVx2_ASAP7_75t_L g1484 ( .A(n_885), .Y(n_1484) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_890), .A2(n_894), .B1(n_912), .B2(n_928), .Y(n_927) );
AOI21xp5_ASAP7_75t_L g1091 ( .A1(n_891), .A2(n_1092), .B(n_1098), .Y(n_1091) );
INVx1_ASAP7_75t_L g1346 ( .A(n_891), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g1459 ( .A1(n_891), .A2(n_1460), .B1(n_1461), .B2(n_1462), .C(n_1463), .Y(n_1459) );
AOI221xp5_ASAP7_75t_L g1485 ( .A1(n_891), .A2(n_1486), .B1(n_1487), .B2(n_1488), .C(n_1493), .Y(n_1485) );
BUFx3_ASAP7_75t_L g1054 ( .A(n_892), .Y(n_1054) );
AOI22xp5_ASAP7_75t_L g1378 ( .A1(n_897), .A2(n_1213), .B1(n_1379), .B2(n_1397), .Y(n_1378) );
NOR3xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_907), .C(n_910), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_903), .Y(n_899) );
OAI22xp33_ASAP7_75t_L g1416 ( .A1(n_912), .A2(n_1229), .B1(n_1387), .B2(n_1393), .Y(n_1416) );
OAI22xp33_ASAP7_75t_L g1552 ( .A1(n_912), .A2(n_1553), .B1(n_1554), .B2(n_1555), .Y(n_1552) );
INVx2_ASAP7_75t_SL g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g972 ( .A(n_913), .Y(n_972) );
INVx1_ASAP7_75t_L g1413 ( .A(n_913), .Y(n_1413) );
INVx2_ASAP7_75t_SL g913 ( .A(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_918), .A2(n_1409), .B1(n_1410), .B2(n_1411), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1417 ( .A1(n_918), .A2(n_1394), .B1(n_1396), .B2(n_1418), .Y(n_1417) );
BUFx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
BUFx2_ASAP7_75t_L g1333 ( .A(n_919), .Y(n_1333) );
INVx2_ASAP7_75t_SL g1559 ( .A(n_921), .Y(n_1559) );
OAI22xp5_ASAP7_75t_L g1561 ( .A1(n_921), .A2(n_1516), .B1(n_1529), .B2(n_1540), .Y(n_1561) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
XNOR2x2_ASAP7_75t_L g935 ( .A(n_936), .B(n_1161), .Y(n_935) );
AO22x2_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_1113), .B1(n_1159), .B2(n_1160), .Y(n_936) );
INVx1_ASAP7_75t_L g1159 ( .A(n_937), .Y(n_1159) );
XNOR2xp5_ASAP7_75t_L g937 ( .A(n_938), .B(n_999), .Y(n_937) );
NAND4xp75_ASAP7_75t_L g939 ( .A(n_940), .B(n_960), .C(n_991), .D(n_995), .Y(n_939) );
AND2x2_ASAP7_75t_SL g940 ( .A(n_941), .B(n_956), .Y(n_940) );
AOI33xp33_ASAP7_75t_L g941 ( .A1(n_942), .A2(n_943), .A3(n_947), .B1(n_950), .B2(n_951), .B3(n_955), .Y(n_941) );
AOI33xp33_ASAP7_75t_L g2014 ( .A1(n_942), .A2(n_1270), .A3(n_2015), .B1(n_2017), .B2(n_2018), .B3(n_2019), .Y(n_2014) );
BUFx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
BUFx3_ASAP7_75t_L g952 ( .A(n_945), .Y(n_952) );
INVx1_ASAP7_75t_L g1144 ( .A(n_945), .Y(n_1144) );
INVx2_ASAP7_75t_L g1657 ( .A(n_945), .Y(n_1657) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_969), .B1(n_974), .B2(n_979), .C(n_984), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_965), .A2(n_966), .B1(n_967), .B2(n_968), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_968), .A2(n_1332), .B1(n_1333), .B2(n_1334), .Y(n_1331) );
INVx1_ASAP7_75t_L g2008 ( .A(n_968), .Y(n_2008) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_975), .A2(n_980), .B1(n_996), .B2(n_998), .Y(n_995) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OAI221xp5_ASAP7_75t_L g1235 ( .A1(n_983), .A2(n_1236), .B1(n_1237), .B2(n_1238), .C(n_1239), .Y(n_1235) );
AOI21xp5_ASAP7_75t_L g984 ( .A1(n_985), .A2(n_986), .B(n_987), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_992), .A2(n_996), .B1(n_1239), .B2(n_1243), .Y(n_1254) );
AOI221xp5_ASAP7_75t_L g1310 ( .A1(n_992), .A2(n_996), .B1(n_1311), .B2(n_1312), .C(n_1313), .Y(n_1310) );
AND2x2_ASAP7_75t_L g996 ( .A(n_993), .B(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_994), .A2(n_998), .B1(n_1237), .B2(n_1244), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_997), .A2(n_1330), .B1(n_1332), .B2(n_1345), .Y(n_1344) );
XNOR2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1056), .Y(n_999) );
NAND3xp33_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1019), .C(n_1028), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1018), .Y(n_1002) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1009), .B2(n_1010), .C(n_1011), .Y(n_1006) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1007), .Y(n_1242) );
BUFx2_ASAP7_75t_L g1439 ( .A(n_1012), .Y(n_1439) );
NAND3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1016), .C(n_1017), .Y(n_1013) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1015), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g1431 ( .A(n_1015), .Y(n_1431) );
NOR2xp33_ASAP7_75t_SL g1019 ( .A(n_1020), .B(n_1025), .Y(n_1019) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1022), .Y(n_1338) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVxp67_ASAP7_75t_L g1339 ( .A(n_1024), .Y(n_1339) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
OAI31xp33_ASAP7_75t_SL g1028 ( .A1(n_1029), .A2(n_1031), .A3(n_1033), .B(n_1055), .Y(n_1028) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1030), .Y(n_1451) );
OAI211xp5_ASAP7_75t_SL g1033 ( .A1(n_1034), .A2(n_1038), .B(n_1042), .C(n_1047), .Y(n_1033) );
INVx2_ASAP7_75t_L g1610 ( .A(n_1037), .Y(n_1610) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
NAND2xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1051), .Y(n_1049) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1050), .Y(n_1351) );
NAND2xp5_ASAP7_75t_SL g1056 ( .A(n_1057), .B(n_1109), .Y(n_1056) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1058), .Y(n_1111) );
NAND3xp33_ASAP7_75t_SL g1058 ( .A(n_1059), .B(n_1062), .C(n_1070), .Y(n_1058) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1068), .B2(n_1069), .Y(n_1062) );
BUFx2_ASAP7_75t_L g1426 ( .A(n_1063), .Y(n_1426) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_1068), .A2(n_1102), .B1(n_1105), .B2(n_1106), .Y(n_1101) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1072), .Y(n_1435) );
BUFx3_ASAP7_75t_L g1130 ( .A(n_1077), .Y(n_1130) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1083), .Y(n_1110) );
AOI31xp33_ASAP7_75t_SL g1083 ( .A1(n_1084), .A2(n_1091), .A3(n_1101), .B(n_1108), .Y(n_1083) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1088), .Y(n_1100) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1095), .Y(n_1263) );
INVxp67_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx3_ASAP7_75t_L g1492 ( .A(n_1097), .Y(n_1492) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1097), .Y(n_1665) );
HB1xp67_ASAP7_75t_L g1262 ( .A(n_1103), .Y(n_1262) );
BUFx3_ASAP7_75t_L g1618 ( .A(n_1103), .Y(n_1618) );
HB1xp67_ASAP7_75t_L g1616 ( .A(n_1104), .Y(n_1616) );
HB1xp67_ASAP7_75t_L g1990 ( .A(n_1104), .Y(n_1990) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
NAND3xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .C(n_1112), .Y(n_1109) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1113), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1135), .Y(n_1114) );
AND4x1_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1119), .C(n_1122), .D(n_1125), .Y(n_1115) );
AOI33xp33_ASAP7_75t_L g1927 ( .A1(n_1126), .A2(n_1928), .A3(n_1932), .B1(n_1934), .B2(n_1935), .B3(n_1936), .Y(n_1927) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g1240 ( .A1(n_1132), .A2(n_1241), .B1(n_1243), .B2(n_1244), .Y(n_1240) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_1146), .A2(n_1295), .B1(n_1296), .B2(n_1303), .C(n_1305), .Y(n_1302) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g1161 ( .A1(n_1162), .A2(n_1275), .B1(n_1369), .B2(n_1370), .Y(n_1161) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1162), .Y(n_1369) );
XNOR2xp5_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1216), .Y(n_1162) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1188), .Y(n_1165) );
AND4x1_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1173), .C(n_1177), .D(n_1181), .Y(n_1166) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
AOI21xp33_ASAP7_75t_SL g1188 ( .A1(n_1189), .A2(n_1190), .B(n_1191), .Y(n_1188) );
AOI31xp33_ASAP7_75t_L g1191 ( .A1(n_1192), .A2(n_1200), .A3(n_1209), .B(n_1212), .Y(n_1191) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
CKINVDCx8_ASAP7_75t_R g1213 ( .A(n_1214), .Y(n_1213) );
OAI31xp33_ASAP7_75t_L g1219 ( .A1(n_1214), .A2(n_1220), .A3(n_1221), .B(n_1234), .Y(n_1219) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
NAND3xp33_ASAP7_75t_SL g1218 ( .A(n_1219), .B(n_1249), .C(n_1251), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1225), .B1(n_1226), .B2(n_1227), .Y(n_1222) );
OAI22xp5_ASAP7_75t_L g1589 ( .A1(n_1223), .A2(n_1590), .B1(n_1591), .B2(n_1593), .Y(n_1589) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx2_ASAP7_75t_L g1512 ( .A(n_1224), .Y(n_1512) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1224), .Y(n_1516) );
INVx2_ASAP7_75t_L g1595 ( .A(n_1224), .Y(n_1595) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1230), .Y(n_1236) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1230), .Y(n_1554) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
NOR2xp33_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1255), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1254), .Y(n_1252) );
NAND3xp33_ASAP7_75t_SL g1255 ( .A(n_1256), .B(n_1258), .C(n_1271), .Y(n_1255) );
AOI33xp33_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1260), .A3(n_1261), .B1(n_1264), .B2(n_1266), .B3(n_1270), .Y(n_1258) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
HB1xp67_ASAP7_75t_L g1370 ( .A(n_1276), .Y(n_1370) );
XNOR2x1_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1316), .Y(n_1276) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1278), .Y(n_1314) );
NAND4xp25_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1297), .C(n_1299), .D(n_1310), .Y(n_1278) );
AOI21xp5_ASAP7_75t_L g1284 ( .A1(n_1285), .A2(n_1286), .B(n_1287), .Y(n_1284) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1291), .B1(n_1292), .B2(n_1293), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_1290), .A2(n_1320), .B1(n_1321), .B2(n_1322), .Y(n_1319) );
INVx2_ASAP7_75t_SL g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1304), .Y(n_1357) );
INVx1_ASAP7_75t_SL g1368 ( .A(n_1317), .Y(n_1368) );
NAND4xp75_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1336), .C(n_1341), .D(n_1364), .Y(n_1317) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
OAI211xp5_ASAP7_75t_L g1356 ( .A1(n_1326), .A2(n_1357), .B(n_1358), .C(n_1359), .Y(n_1356) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1328), .Y(n_1564) );
BUFx2_ASAP7_75t_L g1584 ( .A(n_1328), .Y(n_1584) );
NOR2x1_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1340), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1356), .Y(n_1347) );
OAI211xp5_ASAP7_75t_L g1348 ( .A1(n_1349), .A2(n_1350), .B(n_1352), .C(n_1353), .Y(n_1348) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1355), .Y(n_1661) );
OAI22xp5_ASAP7_75t_L g1726 ( .A1(n_1367), .A2(n_1681), .B1(n_1690), .B2(n_1727), .Y(n_1726) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1566), .B1(n_1567), .B2(n_1671), .Y(n_1372) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1373), .Y(n_1671) );
XNOR2x2_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1472), .Y(n_1373) );
XNOR2xp5_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1419), .Y(n_1374) );
XNOR2xp5_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1377), .Y(n_1375) );
OAI22xp33_ASAP7_75t_L g1763 ( .A1(n_1376), .A2(n_1764), .B1(n_1765), .B2(n_1766), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1378), .B(n_1398), .Y(n_1377) );
NAND4xp25_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1386), .C(n_1392), .D(n_1395), .Y(n_1379) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
NOR3xp33_ASAP7_75t_SL g1398 ( .A(n_1399), .B(n_1406), .C(n_1407), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1403), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1511 ( .A1(n_1410), .A2(n_1512), .B1(n_1513), .B2(n_1514), .Y(n_1511) );
OAI22xp5_ASAP7_75t_L g1515 ( .A1(n_1418), .A2(n_1478), .B1(n_1496), .B2(n_1516), .Y(n_1515) );
XNOR2x1_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1471), .Y(n_1419) );
NAND2x1_ASAP7_75t_L g1420 ( .A(n_1421), .B(n_1447), .Y(n_1420) );
AND4x1_ASAP7_75t_L g1421 ( .A(n_1422), .B(n_1425), .C(n_1440), .D(n_1444), .Y(n_1421) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
INVx2_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
AOI22xp5_ASAP7_75t_L g1447 ( .A1(n_1448), .A2(n_1449), .B1(n_1469), .B2(n_1470), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g1475 ( .A1(n_1448), .A2(n_1470), .B1(n_1476), .B2(n_1497), .Y(n_1475) );
NAND3xp33_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1459), .C(n_1466), .Y(n_1449) );
AOI21xp5_ASAP7_75t_SL g1450 ( .A1(n_1451), .A2(n_1452), .B(n_1453), .Y(n_1450) );
HB1xp67_ASAP7_75t_L g1953 ( .A(n_1464), .Y(n_1953) );
AOI21xp5_ASAP7_75t_L g1937 ( .A1(n_1470), .A2(n_1938), .B(n_1939), .Y(n_1937) );
XNOR2xp5_ASAP7_75t_L g1472 ( .A(n_1473), .B(n_1519), .Y(n_1472) );
XOR2x2_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1518), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_1475), .B(n_1498), .Y(n_1474) );
NAND3xp33_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1485), .C(n_1494), .Y(n_1476) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1482), .Y(n_1534) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
NOR3xp33_ASAP7_75t_L g1498 ( .A(n_1499), .B(n_1506), .C(n_1507), .Y(n_1498) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1500), .B(n_1503), .Y(n_1499) );
OAI22xp5_ASAP7_75t_L g1556 ( .A1(n_1512), .A2(n_1557), .B1(n_1558), .B2(n_1560), .Y(n_1556) );
XNOR2x1_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1565), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1542), .Y(n_1520) );
NAND5xp2_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1527), .C(n_1530), .D(n_1533), .E(n_1539), .Y(n_1522) );
OAI221xp5_ASAP7_75t_SL g1533 ( .A1(n_1534), .A2(n_1535), .B1(n_1536), .B2(n_1537), .C(n_1538), .Y(n_1533) );
NOR3xp33_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1548), .C(n_1551), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1546), .Y(n_1543) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
OAI22xp5_ASAP7_75t_L g1567 ( .A1(n_1568), .A2(n_1569), .B1(n_1621), .B2(n_1670), .Y(n_1567) );
INVx2_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
XNOR2x1_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1620), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1602), .Y(n_1570) );
NOR3xp33_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1579), .C(n_1582), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1572 ( .A(n_1573), .B(n_1576), .Y(n_1572) );
OAI22xp33_ASAP7_75t_L g1583 ( .A1(n_1584), .A2(n_1585), .B1(n_1586), .B2(n_1588), .Y(n_1583) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
OAI22xp5_ASAP7_75t_L g1594 ( .A1(n_1595), .A2(n_1596), .B1(n_1597), .B2(n_1598), .Y(n_1594) );
OAI22xp5_ASAP7_75t_L g1640 ( .A1(n_1595), .A2(n_1641), .B1(n_1642), .B2(n_1643), .Y(n_1640) );
INVx2_ASAP7_75t_SL g1609 ( .A(n_1610), .Y(n_1609) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1621), .Y(n_1670) );
XNOR2x1_ASAP7_75t_SL g1621 ( .A(n_1622), .B(n_1623), .Y(n_1621) );
AND2x2_ASAP7_75t_L g1623 ( .A(n_1624), .B(n_1651), .Y(n_1623) );
NOR3xp33_ASAP7_75t_SL g1624 ( .A(n_1625), .B(n_1632), .C(n_1633), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1629), .Y(n_1625) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
NAND3xp33_ASAP7_75t_L g1652 ( .A(n_1653), .B(n_1662), .C(n_1668), .Y(n_1652) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
INVx1_ASAP7_75t_L g1944 ( .A(n_1659), .Y(n_1944) );
INVx1_ASAP7_75t_L g1954 ( .A(n_1659), .Y(n_1954) );
OAI221xp5_ASAP7_75t_L g1672 ( .A1(n_1673), .A2(n_1908), .B1(n_1911), .B2(n_1958), .C(n_1962), .Y(n_1672) );
AOI311xp33_ASAP7_75t_L g1673 ( .A1(n_1674), .A2(n_1767), .A3(n_1795), .B(n_1802), .C(n_1874), .Y(n_1673) );
OAI211xp5_ASAP7_75t_L g1674 ( .A1(n_1675), .A2(n_1703), .B(n_1728), .C(n_1754), .Y(n_1674) );
A2O1A1Ixp33_ASAP7_75t_L g1728 ( .A1(n_1675), .A2(n_1729), .B(n_1733), .C(n_1739), .Y(n_1728) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
NAND2xp5_ASAP7_75t_L g1819 ( .A(n_1676), .B(n_1820), .Y(n_1819) );
AND2x2_ASAP7_75t_L g1901 ( .A(n_1676), .B(n_1796), .Y(n_1901) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
INVx2_ASAP7_75t_SL g1744 ( .A(n_1677), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1778 ( .A(n_1677), .B(n_1736), .Y(n_1778) );
AND2x4_ASAP7_75t_L g1792 ( .A(n_1677), .B(n_1735), .Y(n_1792) );
NAND2xp5_ASAP7_75t_L g1817 ( .A(n_1677), .B(n_1796), .Y(n_1817) );
AND2x2_ASAP7_75t_L g1823 ( .A(n_1677), .B(n_1824), .Y(n_1823) );
NOR2xp33_ASAP7_75t_L g1865 ( .A(n_1677), .B(n_1824), .Y(n_1865) );
HB1xp67_ASAP7_75t_L g1892 ( .A(n_1677), .Y(n_1892) );
CKINVDCx5p33_ASAP7_75t_R g1677 ( .A(n_1678), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1678), .B(n_1736), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1830 ( .A(n_1678), .B(n_1735), .Y(n_1830) );
OR2x2_ASAP7_75t_L g1678 ( .A(n_1679), .B(n_1693), .Y(n_1678) );
OAI22xp5_ASAP7_75t_L g1679 ( .A1(n_1680), .A2(n_1687), .B1(n_1688), .B2(n_1692), .Y(n_1679) );
BUFx3_ASAP7_75t_L g1764 ( .A(n_1680), .Y(n_1764) );
BUFx6f_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
OR2x2_ASAP7_75t_L g1681 ( .A(n_1682), .B(n_1683), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1690 ( .A(n_1682), .B(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1682), .Y(n_1710) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1683), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1686), .Y(n_1683) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1686), .Y(n_1697) );
HB1xp67_ASAP7_75t_L g1766 ( .A(n_1688), .Y(n_1766) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1691), .Y(n_1712) );
OAI22xp5_ASAP7_75t_L g1693 ( .A1(n_1694), .A2(n_1699), .B1(n_1700), .B2(n_1702), .Y(n_1693) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
BUFx3_ASAP7_75t_L g1762 ( .A(n_1695), .Y(n_1762) );
AND2x4_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1698), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1696), .B(n_1698), .Y(n_1719) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
AND2x4_ASAP7_75t_L g1701 ( .A(n_1697), .B(n_1698), .Y(n_1701) );
INVx2_ASAP7_75t_L g1761 ( .A(n_1700), .Y(n_1761) );
INVx2_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
OR2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1714), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1730 ( .A(n_1704), .B(n_1731), .Y(n_1730) );
OAI321xp33_ASAP7_75t_SL g1815 ( .A1(n_1704), .A2(n_1816), .A3(n_1817), .B1(n_1818), .B2(n_1819), .C(n_1821), .Y(n_1815) );
NAND2xp5_ASAP7_75t_L g1827 ( .A(n_1704), .B(n_1746), .Y(n_1827) );
INVx2_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1814 ( .A(n_1705), .B(n_1720), .Y(n_1814) );
NAND2xp5_ASAP7_75t_SL g1849 ( .A(n_1705), .B(n_1850), .Y(n_1849) );
AND2x2_ASAP7_75t_L g1880 ( .A(n_1705), .B(n_1778), .Y(n_1880) );
BUFx2_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1706), .B(n_1743), .Y(n_1742) );
INVx2_ASAP7_75t_L g1750 ( .A(n_1706), .Y(n_1750) );
NAND2xp5_ASAP7_75t_L g1770 ( .A(n_1706), .B(n_1771), .Y(n_1770) );
OR2x2_ASAP7_75t_L g1788 ( .A(n_1706), .B(n_1776), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1807 ( .A(n_1706), .B(n_1732), .Y(n_1807) );
INVx2_ASAP7_75t_L g1824 ( .A(n_1706), .Y(n_1824) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1713), .Y(n_1706) );
AND2x4_ASAP7_75t_L g1708 ( .A(n_1709), .B(n_1710), .Y(n_1708) );
AND2x4_ASAP7_75t_L g1711 ( .A(n_1710), .B(n_1712), .Y(n_1711) );
BUFx2_ASAP7_75t_L g1800 ( .A(n_1711), .Y(n_1800) );
HB1xp67_ASAP7_75t_L g2047 ( .A(n_1712), .Y(n_2047) );
INVx2_ASAP7_75t_L g1755 ( .A(n_1714), .Y(n_1755) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1715), .B(n_1720), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1715), .B(n_1742), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1715), .B(n_1752), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1715), .B(n_1747), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1715), .B(n_1757), .Y(n_1777) );
INVxp67_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
BUFx2_ASAP7_75t_L g1732 ( .A(n_1716), .Y(n_1732) );
BUFx3_ASAP7_75t_L g1776 ( .A(n_1716), .Y(n_1776) );
OR2x2_ASAP7_75t_L g1860 ( .A(n_1716), .B(n_1725), .Y(n_1860) );
AND2x2_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1718), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1775 ( .A(n_1720), .B(n_1776), .Y(n_1775) );
NOR2xp33_ASAP7_75t_L g1858 ( .A(n_1720), .B(n_1859), .Y(n_1858) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1720), .Y(n_1869) );
NAND3xp33_ASAP7_75t_SL g1887 ( .A(n_1720), .B(n_1749), .C(n_1811), .Y(n_1887) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1724), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1721), .B(n_1725), .Y(n_1743) );
INVx2_ASAP7_75t_L g1748 ( .A(n_1721), .Y(n_1748) );
OR2x2_ASAP7_75t_L g1753 ( .A(n_1721), .B(n_1725), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1822 ( .A(n_1721), .B(n_1776), .Y(n_1822) );
NOR2xp33_ASAP7_75t_L g1850 ( .A(n_1721), .B(n_1776), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1722), .B(n_1723), .Y(n_1721) );
NOR2x1_ASAP7_75t_L g1731 ( .A(n_1724), .B(n_1732), .Y(n_1731) );
AND2x2_ASAP7_75t_L g1873 ( .A(n_1724), .B(n_1776), .Y(n_1873) );
INVx2_ASAP7_75t_SL g1724 ( .A(n_1725), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1725), .B(n_1748), .Y(n_1747) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
NOR2xp33_ASAP7_75t_L g1885 ( .A(n_1730), .B(n_1832), .Y(n_1885) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1731), .Y(n_1871) );
AND2x2_ASAP7_75t_L g1746 ( .A(n_1732), .B(n_1747), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_1732), .B(n_1743), .Y(n_1794) );
A2O1A1Ixp33_ASAP7_75t_L g1739 ( .A1(n_1733), .A2(n_1740), .B(n_1744), .C(n_1745), .Y(n_1739) );
OAI221xp5_ASAP7_75t_L g1779 ( .A1(n_1733), .A2(n_1734), .B1(n_1780), .B2(n_1782), .C(n_1784), .Y(n_1779) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
AOI22xp33_ASAP7_75t_L g1889 ( .A1(n_1734), .A2(n_1768), .B1(n_1830), .B2(n_1890), .Y(n_1889) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1820 ( .A(n_1735), .B(n_1798), .Y(n_1820) );
OR2x2_ASAP7_75t_L g1832 ( .A(n_1735), .B(n_1833), .Y(n_1832) );
INVx3_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
OR2x2_ASAP7_75t_L g1856 ( .A(n_1736), .B(n_1798), .Y(n_1856) );
AND2x2_ASAP7_75t_L g1897 ( .A(n_1736), .B(n_1797), .Y(n_1897) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1737), .B(n_1738), .Y(n_1736) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1818 ( .A(n_1742), .Y(n_1818) );
O2A1O1Ixp33_ASAP7_75t_L g1875 ( .A1(n_1742), .A2(n_1876), .B(n_1877), .C(n_1878), .Y(n_1875) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1743), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1783 ( .A(n_1743), .B(n_1750), .Y(n_1783) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1744), .B(n_1750), .Y(n_1749) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1744), .Y(n_1769) );
NOR2xp33_ASAP7_75t_L g1786 ( .A(n_1744), .B(n_1787), .Y(n_1786) );
NOR2xp33_ASAP7_75t_L g1846 ( .A(n_1744), .B(n_1832), .Y(n_1846) );
INVx2_ASAP7_75t_L g1854 ( .A(n_1744), .Y(n_1854) );
AOI21xp33_ASAP7_75t_SL g1745 ( .A1(n_1746), .A2(n_1749), .B(n_1751), .Y(n_1745) );
OAI211xp5_ASAP7_75t_L g1843 ( .A1(n_1746), .A2(n_1824), .B(n_1830), .C(n_1844), .Y(n_1843) );
A2O1A1Ixp33_ASAP7_75t_SL g1888 ( .A1(n_1746), .A2(n_1862), .B(n_1889), .C(n_1894), .Y(n_1888) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1747), .B(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1747), .Y(n_1838) );
NAND2xp5_ASAP7_75t_L g1816 ( .A(n_1748), .B(n_1776), .Y(n_1816) );
OAI321xp33_ASAP7_75t_L g1878 ( .A1(n_1748), .A2(n_1867), .A3(n_1879), .B1(n_1881), .B2(n_1882), .C(n_1884), .Y(n_1878) );
NOR2xp33_ASAP7_75t_L g1752 ( .A(n_1750), .B(n_1753), .Y(n_1752) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1750), .B(n_1757), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1883 ( .A(n_1750), .B(n_1822), .Y(n_1883) );
INVx1_ASAP7_75t_L g1893 ( .A(n_1751), .Y(n_1893) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1753), .Y(n_1757) );
OR2x2_ASAP7_75t_L g1787 ( .A(n_1753), .B(n_1788), .Y(n_1787) );
NOR2xp33_ASAP7_75t_L g1828 ( .A(n_1753), .B(n_1829), .Y(n_1828) );
O2A1O1Ixp33_ASAP7_75t_L g1754 ( .A1(n_1755), .A2(n_1756), .B(n_1758), .C(n_1759), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1876 ( .A(n_1756), .B(n_1776), .Y(n_1876) );
AND2x2_ASAP7_75t_L g1855 ( .A(n_1757), .B(n_1807), .Y(n_1855) );
CKINVDCx5p33_ASAP7_75t_R g1812 ( .A(n_1758), .Y(n_1812) );
AOI211xp5_ASAP7_75t_SL g1825 ( .A1(n_1758), .A2(n_1826), .B(n_1828), .C(n_1831), .Y(n_1825) );
NAND4xp25_ASAP7_75t_L g1905 ( .A(n_1758), .B(n_1807), .C(n_1844), .D(n_1906), .Y(n_1905) );
INVx3_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
INVx3_ASAP7_75t_L g1784 ( .A(n_1760), .Y(n_1784) );
A2O1A1Ixp33_ASAP7_75t_SL g1802 ( .A1(n_1760), .A2(n_1803), .B(n_1825), .C(n_1841), .Y(n_1802) );
AND2x2_ASAP7_75t_L g1862 ( .A(n_1760), .B(n_1863), .Y(n_1862) );
BUFx2_ASAP7_75t_SL g1910 ( .A(n_1766), .Y(n_1910) );
NAND4xp25_ASAP7_75t_L g1767 ( .A(n_1768), .B(n_1772), .C(n_1785), .D(n_1789), .Y(n_1767) );
OR2x2_ASAP7_75t_L g1768 ( .A(n_1769), .B(n_1770), .Y(n_1768) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1770), .Y(n_1896) );
AOI21xp33_ASAP7_75t_L g1772 ( .A1(n_1773), .A2(n_1778), .B(n_1779), .Y(n_1772) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
NOR2xp33_ASAP7_75t_L g1774 ( .A(n_1775), .B(n_1777), .Y(n_1774) );
OR2x2_ASAP7_75t_L g1780 ( .A(n_1776), .B(n_1781), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1835 ( .A(n_1776), .B(n_1783), .Y(n_1835) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1777), .Y(n_1866) );
AOI221xp5_ASAP7_75t_L g1803 ( .A1(n_1778), .A2(n_1804), .B1(n_1808), .B2(n_1813), .C(n_1815), .Y(n_1803) );
AOI21xp5_ASAP7_75t_L g1894 ( .A1(n_1778), .A2(n_1792), .B(n_1834), .Y(n_1894) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1780), .Y(n_1851) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
NAND2xp5_ASAP7_75t_L g1795 ( .A(n_1784), .B(n_1796), .Y(n_1795) );
O2A1O1Ixp33_ASAP7_75t_L g1852 ( .A1(n_1784), .A2(n_1814), .B(n_1853), .C(n_1856), .Y(n_1852) );
OAI211xp5_ASAP7_75t_L g1874 ( .A1(n_1784), .A2(n_1875), .B(n_1888), .C(n_1895), .Y(n_1874) );
INVxp67_ASAP7_75t_SL g1785 ( .A(n_1786), .Y(n_1785) );
O2A1O1Ixp33_ASAP7_75t_L g1895 ( .A1(n_1786), .A2(n_1896), .B(n_1897), .C(n_1898), .Y(n_1895) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1787), .B(n_1805), .Y(n_1804) );
NOR2xp33_ASAP7_75t_L g1904 ( .A(n_1787), .B(n_1892), .Y(n_1904) );
OR2x2_ASAP7_75t_L g1868 ( .A(n_1788), .B(n_1869), .Y(n_1868) );
INVxp67_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
NOR2xp33_ASAP7_75t_L g1790 ( .A(n_1791), .B(n_1793), .Y(n_1790) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
AND2x2_ASAP7_75t_L g1840 ( .A(n_1792), .B(n_1796), .Y(n_1840) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
OAI332xp33_ASAP7_75t_L g1857 ( .A1(n_1795), .A2(n_1854), .A3(n_1858), .B1(n_1861), .B2(n_1864), .B3(n_1866), .C1(n_1867), .C2(n_1868), .Y(n_1857) );
INVx2_ASAP7_75t_L g1844 ( .A(n_1796), .Y(n_1844) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1797), .Y(n_1796) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1797), .Y(n_1811) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1798), .Y(n_1833) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1798), .Y(n_1881) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1799), .B(n_1801), .Y(n_1798) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1806), .Y(n_1805) );
NAND2xp5_ASAP7_75t_L g1845 ( .A(n_1806), .B(n_1846), .Y(n_1845) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
OR2x2_ASAP7_75t_L g1809 ( .A(n_1810), .B(n_1812), .Y(n_1809) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1811), .Y(n_1810) );
INVx1_ASAP7_75t_L g1863 ( .A(n_1811), .Y(n_1863) );
AOI211xp5_ASAP7_75t_L g1870 ( .A1(n_1811), .A2(n_1829), .B(n_1871), .C(n_1872), .Y(n_1870) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
INVx1_ASAP7_75t_L g1877 ( .A(n_1817), .Y(n_1877) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1820), .Y(n_1867) );
NAND2xp5_ASAP7_75t_L g1821 ( .A(n_1822), .B(n_1823), .Y(n_1821) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1824), .B(n_1830), .Y(n_1829) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
OAI21xp33_ASAP7_75t_L g1831 ( .A1(n_1832), .A2(n_1834), .B(n_1836), .Y(n_1831) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
INVxp33_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
NOR2xp33_ASAP7_75t_L g1837 ( .A(n_1838), .B(n_1839), .Y(n_1837) );
NAND2xp5_ASAP7_75t_L g1907 ( .A(n_1838), .B(n_1869), .Y(n_1907) );
INVx1_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
OAI21xp5_ASAP7_75t_L g1847 ( .A1(n_1840), .A2(n_1848), .B(n_1851), .Y(n_1847) );
NOR4xp25_ASAP7_75t_L g1841 ( .A(n_1842), .B(n_1852), .C(n_1857), .D(n_1870), .Y(n_1841) );
NAND3xp33_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1845), .C(n_1847), .Y(n_1842) );
A2O1A1Ixp33_ASAP7_75t_L g1898 ( .A1(n_1844), .A2(n_1899), .B(n_1903), .C(n_1905), .Y(n_1898) );
INVx1_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
NAND2xp5_ASAP7_75t_L g1853 ( .A(n_1854), .B(n_1855), .Y(n_1853) );
INVx1_ASAP7_75t_L g1859 ( .A(n_1860), .Y(n_1859) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1862), .Y(n_1861) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
INVxp67_ASAP7_75t_L g1902 ( .A(n_1868), .Y(n_1902) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1883), .Y(n_1882) );
NOR2xp33_ASAP7_75t_L g1884 ( .A(n_1885), .B(n_1886), .Y(n_1884) );
INVx1_ASAP7_75t_L g1886 ( .A(n_1887), .Y(n_1886) );
INVxp33_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
NOR2xp33_ASAP7_75t_L g1891 ( .A(n_1892), .B(n_1893), .Y(n_1891) );
NAND2xp5_ASAP7_75t_L g1899 ( .A(n_1900), .B(n_1902), .Y(n_1899) );
INVx1_ASAP7_75t_L g1900 ( .A(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g1903 ( .A(n_1904), .Y(n_1903) );
INVx1_ASAP7_75t_L g1906 ( .A(n_1907), .Y(n_1906) );
CKINVDCx5p33_ASAP7_75t_R g1908 ( .A(n_1909), .Y(n_1908) );
INVx1_ASAP7_75t_SL g1909 ( .A(n_1910), .Y(n_1909) );
INVx1_ASAP7_75t_L g1913 ( .A(n_1914), .Y(n_1913) );
BUFx2_ASAP7_75t_L g1914 ( .A(n_1915), .Y(n_1914) );
NAND2xp5_ASAP7_75t_L g1915 ( .A(n_1916), .B(n_1937), .Y(n_1915) );
AND4x1_ASAP7_75t_L g1916 ( .A(n_1917), .B(n_1920), .C(n_1923), .D(n_1927), .Y(n_1916) );
INVx1_ASAP7_75t_L g1930 ( .A(n_1931), .Y(n_1930) );
INVx1_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
CKINVDCx5p33_ASAP7_75t_R g1958 ( .A(n_1959), .Y(n_1958) );
BUFx2_ASAP7_75t_L g1959 ( .A(n_1960), .Y(n_1959) );
OAI21xp5_ASAP7_75t_L g2046 ( .A1(n_1961), .A2(n_2047), .B(n_2048), .Y(n_2046) );
INVx1_ASAP7_75t_L g1963 ( .A(n_1964), .Y(n_1963) );
INVx1_ASAP7_75t_L g1964 ( .A(n_1965), .Y(n_1964) );
INVx1_ASAP7_75t_L g1965 ( .A(n_1966), .Y(n_1965) );
INVx1_ASAP7_75t_L g1966 ( .A(n_1967), .Y(n_1966) );
INVx1_ASAP7_75t_L g2044 ( .A(n_1969), .Y(n_2044) );
AOI211x1_ASAP7_75t_SL g1969 ( .A1(n_1970), .A2(n_2001), .B(n_2004), .C(n_2020), .Y(n_1969) );
NAND4xp25_ASAP7_75t_SL g1970 ( .A(n_1971), .B(n_1981), .C(n_1988), .D(n_1998), .Y(n_1970) );
AOI22xp33_ASAP7_75t_L g1971 ( .A1(n_1972), .A2(n_1973), .B1(n_1977), .B2(n_1978), .Y(n_1971) );
AND2x4_ASAP7_75t_L g1973 ( .A(n_1974), .B(n_1976), .Y(n_1973) );
INVx1_ASAP7_75t_SL g1974 ( .A(n_1975), .Y(n_1974) );
INVx1_ASAP7_75t_L g2000 ( .A(n_1979), .Y(n_2000) );
INVx1_ASAP7_75t_L g1979 ( .A(n_1980), .Y(n_1979) );
AOI22xp33_ASAP7_75t_L g1981 ( .A1(n_1982), .A2(n_1983), .B1(n_1986), .B2(n_1987), .Y(n_1981) );
AOI22xp33_ASAP7_75t_L g2038 ( .A1(n_1982), .A2(n_2039), .B1(n_2040), .B2(n_2041), .Y(n_2038) );
AND2x4_ASAP7_75t_L g1993 ( .A(n_1984), .B(n_1994), .Y(n_1993) );
INVx1_ASAP7_75t_L g1984 ( .A(n_1985), .Y(n_1984) );
AOI222xp33_ASAP7_75t_L g1988 ( .A1(n_1989), .A2(n_1990), .B1(n_1991), .B2(n_1992), .C1(n_1996), .C2(n_1997), .Y(n_1988) );
BUFx4f_ASAP7_75t_L g1992 ( .A(n_1993), .Y(n_1992) );
INVx1_ASAP7_75t_L g1994 ( .A(n_1995), .Y(n_1994) );
INVx5_ASAP7_75t_L g1998 ( .A(n_1999), .Y(n_1998) );
BUFx6f_ASAP7_75t_L g2001 ( .A(n_2002), .Y(n_2001) );
NAND2xp5_ASAP7_75t_L g2004 ( .A(n_2005), .B(n_2014), .Y(n_2004) );
INVx1_ASAP7_75t_L g2012 ( .A(n_2013), .Y(n_2012) );
AOI31xp33_ASAP7_75t_L g2020 ( .A1(n_2021), .A2(n_2030), .A3(n_2038), .B(n_2043), .Y(n_2020) );
INVx1_ASAP7_75t_L g2024 ( .A(n_2025), .Y(n_2024) );
INVx2_ASAP7_75t_L g2027 ( .A(n_2028), .Y(n_2027) );
AOI22xp33_ASAP7_75t_L g2030 ( .A1(n_2031), .A2(n_2033), .B1(n_2034), .B2(n_2037), .Y(n_2030) );
AND2x4_ASAP7_75t_L g2034 ( .A(n_2032), .B(n_2035), .Y(n_2034) );
INVx1_ASAP7_75t_L g2035 ( .A(n_2036), .Y(n_2035) );
INVx5_ASAP7_75t_L g2041 ( .A(n_2042), .Y(n_2041) );
BUFx2_ASAP7_75t_L g2045 ( .A(n_2046), .Y(n_2045) );
endmodule