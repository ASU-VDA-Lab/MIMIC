module real_jpeg_11733_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_37),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_37),
.B1(n_62),
.B2(n_63),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_3),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_4),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_145),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_145),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_145),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_5),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_59),
.B(n_62),
.C(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_5),
.B(n_101),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_5),
.B(n_32),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_SL g246 ( 
.A1(n_5),
.A2(n_32),
.B(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_5),
.B(n_46),
.C(n_51),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_180),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_5),
.A2(n_85),
.B1(n_86),
.B2(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_41),
.Y(n_281)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_66),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_66),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_183),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_183),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_183),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_13),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_172),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_172),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_172),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_40),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_15),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_120),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_102),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_19),
.B(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_83),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_20),
.B(n_73),
.CI(n_83),
.CON(n_147),
.SN(n_147)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_57),
.B2(n_72),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_56),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_23),
.B(n_56),
.C(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_35),
.B(n_38),
.Y(n_24)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_25),
.A2(n_38),
.B(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_25),
.A2(n_26),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_25),
.A2(n_26),
.B1(n_186),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_25),
.A2(n_111),
.B(n_187),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_25),
.A2(n_26),
.B1(n_206),
.B2(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_26),
.A2(n_81),
.B(n_114),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_27),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_27),
.A2(n_29),
.B(n_231),
.C(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_27),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_SL g233 ( 
.A(n_28),
.B(n_30),
.C(n_33),
.Y(n_233)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_32),
.A2(n_60),
.B(n_180),
.Y(n_199)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_36),
.A2(n_41),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_39),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_41),
.B(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_42),
.A2(n_56),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_49),
.B(n_53),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_43),
.A2(n_53),
.B(n_95),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_43),
.A2(n_75),
.B(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_44),
.A2(n_76),
.B1(n_93),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_44),
.A2(n_76),
.B1(n_227),
.B2(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_44),
.A2(n_76),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_44),
.A2(n_76),
.B1(n_248),
.B2(n_258),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_49),
.A2(n_77),
.B(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_49),
.B(n_180),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_50),
.B(n_267),
.Y(n_266)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_72),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B(n_67),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_61),
.B1(n_69),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_58),
.A2(n_69),
.B1(n_144),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_58),
.A2(n_69),
.B1(n_171),
.B2(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_70)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_68),
.A2(n_101),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_98),
.B(n_100),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_73),
.A2(n_74),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B(n_96),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_96),
.B1(n_97),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_84),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_84),
.A2(n_91),
.B1(n_92),
.B2(n_126),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_85),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_85),
.A2(n_86),
.B1(n_261),
.B2(n_269),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_85),
.A2(n_135),
.B(n_263),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_86),
.B(n_180),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_89),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_87),
.A2(n_163),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_87),
.A2(n_136),
.B(n_196),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_87),
.A2(n_195),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_89),
.A2(n_165),
.B(n_195),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_125),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_101),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_115),
.B2(n_116),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_148),
.B(n_310),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_147),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_123),
.B(n_147),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_128),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_127),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_129),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_142),
.C(n_143),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_131),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_132),
.A2(n_133),
.B1(n_138),
.B2(n_139),
.Y(n_298)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_143),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g313 ( 
.A(n_147),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_173),
.B(n_309),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_150),
.B(n_153),
.Y(n_309)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.C(n_159),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_158),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_159),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.C(n_169),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_160),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_166),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_300)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_303),
.B(n_308),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_216),
.B(n_294),
.C(n_302),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_207),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_176),
.B(n_207),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_191),
.C(n_200),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_188),
.C(n_190),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_192),
.B1(n_200),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_205),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_208),
.B(n_214),
.C(n_215),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_292),
.B(n_293),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_236),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_219),
.B(n_222),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_228),
.B1(n_229),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_234),
.B1(n_235),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_249),
.B(n_291),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_241),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_247),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_285),
.B(n_290),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_275),
.B(n_284),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_264),
.B(n_274),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_256),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_270),
.B(n_273),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_277),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_280),
.C(n_283),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_289),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_301),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_301),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);


endmodule