module fake_netlist_1_8809_n_1381 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1381);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1381;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_298;
wire n_411;
wire n_1341;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g292 ( .A(n_126), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_233), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_215), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_136), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_178), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_236), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_148), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_96), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_138), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_208), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_165), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_255), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_90), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_50), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_214), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_252), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_114), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_111), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_231), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_153), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_282), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_86), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_219), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_160), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_128), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_173), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_15), .Y(n_319) );
INVxp33_ASAP7_75t_L g320 ( .A(n_60), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_270), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_184), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_281), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_15), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_217), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_38), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_197), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_146), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_66), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_85), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_5), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_46), .Y(n_332) );
INVxp67_ASAP7_75t_SL g333 ( .A(n_285), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_266), .Y(n_334) );
INVxp67_ASAP7_75t_SL g335 ( .A(n_30), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_260), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_55), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_177), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_92), .B(n_141), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_287), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_5), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_47), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_121), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_89), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_198), .Y(n_345) );
INVx2_ASAP7_75t_SL g346 ( .A(n_11), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_249), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_3), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_51), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_53), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_118), .Y(n_351) );
INVx2_ASAP7_75t_SL g352 ( .A(n_137), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_75), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_207), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_191), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_180), .Y(n_356) );
INVxp33_ASAP7_75t_SL g357 ( .A(n_77), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_284), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_76), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_68), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_83), .Y(n_361) );
CKINVDCx16_ASAP7_75t_R g362 ( .A(n_35), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_174), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_39), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_27), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_21), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_228), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_97), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_31), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_17), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_182), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_104), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_216), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_48), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_263), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_254), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_13), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_268), .Y(n_378) );
BUFx5_ASAP7_75t_L g379 ( .A(n_25), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_279), .Y(n_380) );
CKINVDCx16_ASAP7_75t_R g381 ( .A(n_98), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_27), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_22), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_45), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_94), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_91), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_212), .Y(n_387) );
INVxp33_ASAP7_75t_L g388 ( .A(n_53), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_139), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_156), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_21), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_206), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_131), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_258), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_168), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_81), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_251), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_103), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_26), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_218), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_65), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_66), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_64), .Y(n_403) );
INVxp67_ASAP7_75t_SL g404 ( .A(n_199), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_162), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_119), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_1), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_196), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_275), .Y(n_409) );
INVxp33_ASAP7_75t_L g410 ( .A(n_68), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_152), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_3), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_129), .Y(n_413) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_259), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_43), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_147), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_230), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_122), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_262), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_9), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_123), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_245), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_239), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_172), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_221), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_19), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_242), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_192), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_176), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_38), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_246), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_14), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_117), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_203), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_79), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_320), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_379), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_320), .B(n_0), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_379), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_292), .B(n_0), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_388), .B(n_1), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_379), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_295), .B(n_2), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_379), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_362), .Y(n_446) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_392), .B(n_291), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_379), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_295), .B(n_2), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_346), .B(n_4), .Y(n_451) );
AND3x2_ASAP7_75t_L g452 ( .A(n_332), .B(n_4), .C(n_6), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_379), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_314), .B(n_6), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_314), .B(n_7), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_379), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_313), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_319), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_319), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_297), .Y(n_460) );
CKINVDCx5p33_ASAP7_75t_R g461 ( .A(n_381), .Y(n_461) );
XOR2x2_ASAP7_75t_L g462 ( .A(n_426), .B(n_7), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_350), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_328), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_366), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_409), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_346), .B(n_8), .Y(n_467) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_293), .B(n_8), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_352), .B(n_9), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_449), .A2(n_324), .B1(n_331), .B2(n_306), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_447), .B(n_294), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_445), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_464), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_445), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_449), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_436), .B(n_388), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_449), .B(n_329), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_445), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_436), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_438), .B(n_410), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_457), .B(n_352), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_438), .B(n_410), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_457), .B(n_367), .Y(n_485) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_439), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_449), .B(n_329), .Y(n_491) );
INVx5_ASAP7_75t_L g492 ( .A(n_439), .Y(n_492) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_451), .A2(n_403), .B1(n_337), .B2(n_377), .Y(n_493) );
BUFx10_ASAP7_75t_L g494 ( .A(n_449), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_447), .B(n_294), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
AND2x2_ASAP7_75t_SL g497 ( .A(n_447), .B(n_339), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_457), .Y(n_498) );
NAND2xp33_ASAP7_75t_L g499 ( .A(n_460), .B(n_304), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_439), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_439), .Y(n_501) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_450), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_454), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_438), .B(n_348), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_442), .B(n_348), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_457), .B(n_367), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_454), .A2(n_342), .B1(n_349), .B2(n_341), .Y(n_507) );
INVx4_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
INVx4_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_440), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_443), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_443), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_448), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_461), .B(n_340), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_454), .B(n_360), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_448), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_475), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_497), .A2(n_442), .B1(n_469), .B2(n_455), .Y(n_518) );
BUFx4f_ASAP7_75t_L g519 ( .A(n_497), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_475), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_477), .Y(n_521) );
INVx4_ASAP7_75t_L g522 ( .A(n_475), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_477), .Y(n_523) );
AND2x6_ASAP7_75t_L g524 ( .A(n_503), .B(n_469), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_477), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_475), .Y(n_526) );
NOR2xp33_ASAP7_75t_R g527 ( .A(n_473), .B(n_446), .Y(n_527) );
AOI22xp5_ASAP7_75t_SL g528 ( .A1(n_479), .A2(n_403), .B1(n_337), .B2(n_465), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_504), .B(n_469), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_497), .A2(n_442), .B1(n_469), .B2(n_444), .Y(n_532) );
NOR2xp67_ASAP7_75t_L g533 ( .A(n_471), .B(n_469), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_508), .B(n_453), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_479), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_482), .B(n_451), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_476), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_482), .B(n_467), .Y(n_538) );
INVx4_ASAP7_75t_L g539 ( .A(n_508), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_476), .B(n_462), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_476), .B(n_462), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_477), .Y(n_542) );
INVx4_ASAP7_75t_L g543 ( .A(n_508), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_482), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_491), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_508), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_491), .A2(n_453), .B1(n_456), .B2(n_467), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_484), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_484), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_484), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_508), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g552 ( .A1(n_495), .A2(n_456), .B(n_459), .C(n_458), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_509), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_509), .B(n_296), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_509), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_491), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_509), .B(n_298), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_491), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_491), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_515), .A2(n_468), .B1(n_441), .B2(n_459), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_504), .B(n_452), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_504), .Y(n_562) );
INVx4_ASAP7_75t_L g563 ( .A(n_509), .Y(n_563) );
INVx4_ASAP7_75t_L g564 ( .A(n_494), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_515), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_505), .B(n_304), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_515), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_505), .Y(n_569) );
OR2x6_ASAP7_75t_L g570 ( .A(n_505), .B(n_441), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_515), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_515), .B(n_311), .Y(n_572) );
INVx5_ASAP7_75t_L g573 ( .A(n_494), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_470), .B(n_462), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_470), .B(n_311), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_507), .B(n_452), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_507), .B(n_353), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_503), .B(n_468), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_494), .B(n_299), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_503), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_494), .Y(n_581) );
AND2x4_ASAP7_75t_SL g582 ( .A(n_503), .B(n_328), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_480), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_483), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_483), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_514), .B(n_357), .Y(n_586) );
AND2x6_ASAP7_75t_SL g587 ( .A(n_493), .B(n_364), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_SL g588 ( .A1(n_485), .A2(n_305), .B(n_316), .C(n_300), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_506), .B(n_353), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_480), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_485), .B(n_357), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_506), .B(n_359), .Y(n_592) );
BUFx12f_ASAP7_75t_L g593 ( .A(n_493), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_487), .A2(n_458), .B1(n_365), .B2(n_370), .Y(n_594) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_502), .Y(n_595) );
NOR2x2_ASAP7_75t_L g596 ( .A(n_499), .B(n_374), .Y(n_596) );
INVx4_ASAP7_75t_L g597 ( .A(n_480), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_487), .A2(n_369), .B1(n_383), .B2(n_382), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_472), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_488), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_472), .Y(n_601) );
NOR2xp33_ASAP7_75t_R g602 ( .A(n_474), .B(n_374), .Y(n_602) );
AND2x6_ASAP7_75t_SL g603 ( .A(n_488), .B(n_391), .Y(n_603) );
INVx5_ASAP7_75t_L g604 ( .A(n_498), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_474), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_478), .B(n_359), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_489), .A2(n_377), .B1(n_399), .B2(n_384), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_478), .B(n_301), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_580), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_534), .A2(n_498), .B(n_489), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_521), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_534), .A2(n_498), .B(n_510), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_537), .B(n_384), .Y(n_613) );
BUFx8_ASAP7_75t_L g614 ( .A(n_535), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_523), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_602), .Y(n_616) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_573), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_537), .B(n_399), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_562), .A2(n_510), .B(n_512), .C(n_511), .Y(n_619) );
INVx6_ASAP7_75t_SL g620 ( .A(n_561), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_582), .Y(n_621) );
OR2x6_ASAP7_75t_L g622 ( .A(n_593), .B(n_414), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_530), .A2(n_512), .B(n_513), .C(n_511), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_528), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_519), .A2(n_516), .B1(n_513), .B2(n_407), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_525), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_576), .A2(n_401), .B1(n_432), .B2(n_407), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g628 ( .A1(n_530), .A2(n_516), .B(n_402), .C(n_415), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_529), .Y(n_629) );
INVx4_ASAP7_75t_L g630 ( .A(n_573), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_573), .B(n_363), .Y(n_631) );
O2A1O1Ixp5_ASAP7_75t_SL g632 ( .A1(n_608), .A2(n_463), .B(n_302), .C(n_307), .Y(n_632) );
NAND3xp33_ASAP7_75t_SL g633 ( .A(n_527), .B(n_432), .C(n_401), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_562), .A2(n_335), .B(n_420), .C(n_412), .Y(n_634) );
OR2x6_ASAP7_75t_SL g635 ( .A(n_596), .B(n_363), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_600), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_517), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_517), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_574), .A2(n_430), .B1(n_326), .B2(n_350), .C1(n_397), .C2(n_394), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_536), .B(n_373), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_564), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_540), .A2(n_350), .B1(n_380), .B2(n_389), .C(n_373), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_579), .A2(n_321), .B(n_312), .Y(n_643) );
BUFx3_ASAP7_75t_L g644 ( .A(n_582), .Y(n_644) );
INVx5_ASAP7_75t_L g645 ( .A(n_573), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_526), .Y(n_646) );
INVx3_ASAP7_75t_SL g647 ( .A(n_576), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_519), .A2(n_395), .B1(n_405), .B2(n_389), .Y(n_648) );
AOI222xp33_ASAP7_75t_L g649 ( .A1(n_541), .A2(n_350), .B1(n_333), .B2(n_330), .C1(n_368), .C2(n_404), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_602), .Y(n_650) );
OR2x6_ASAP7_75t_L g651 ( .A(n_561), .B(n_303), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_527), .Y(n_652) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_518), .A2(n_310), .B(n_315), .C(n_309), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_550), .A2(n_544), .B1(n_532), .B2(n_548), .Y(n_654) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_584), .A2(n_318), .B(n_322), .C(n_317), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_569), .B(n_434), .Y(n_656) );
NOR2xp33_ASAP7_75t_SL g657 ( .A(n_564), .B(n_395), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_526), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_607), .B(n_538), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_585), .B(n_567), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_601), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_548), .Y(n_662) );
INVx5_ASAP7_75t_L g663 ( .A(n_597), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_542), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_549), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_549), .A2(n_323), .B1(n_334), .B2(n_325), .Y(n_666) );
OR2x6_ASAP7_75t_L g667 ( .A(n_570), .B(n_336), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_587), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_603), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_551), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_545), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_572), .Y(n_672) );
INVx3_ASAP7_75t_L g673 ( .A(n_520), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_556), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_524), .A2(n_338), .B1(n_344), .B2(n_343), .Y(n_675) );
BUFx3_ASAP7_75t_L g676 ( .A(n_578), .Y(n_676) );
XOR2xp5_ASAP7_75t_L g677 ( .A(n_575), .B(n_405), .Y(n_677) );
INVx4_ASAP7_75t_L g678 ( .A(n_520), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_578), .A2(n_351), .B(n_354), .C(n_345), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_558), .Y(n_680) );
BUFx12f_ASAP7_75t_L g681 ( .A(n_570), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_570), .Y(n_682) );
INVx2_ASAP7_75t_SL g683 ( .A(n_577), .Y(n_683) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_522), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_598), .A2(n_425), .B1(n_408), .B2(n_424), .C(n_433), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_547), .B(n_408), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_559), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_606), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_524), .A2(n_355), .B1(n_361), .B2(n_356), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_551), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_589), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_586), .B(n_424), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_565), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_568), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_547), .B(n_425), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_571), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_586), .A2(n_435), .B1(n_433), .B2(n_372), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g698 ( .A1(n_552), .A2(n_375), .B(n_376), .C(n_371), .Y(n_698) );
INVx3_ASAP7_75t_L g699 ( .A(n_522), .Y(n_699) );
OR2x2_ASAP7_75t_L g700 ( .A(n_560), .B(n_435), .Y(n_700) );
INVx4_ASAP7_75t_L g701 ( .A(n_539), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_591), .B(n_308), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_553), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_553), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_591), .A2(n_385), .B1(n_390), .B2(n_386), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_533), .A2(n_393), .B1(n_400), .B2(n_396), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_539), .B(n_406), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_592), .A2(n_411), .B1(n_416), .B2(n_413), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_560), .B(n_327), .Y(n_709) );
OR2x6_ASAP7_75t_L g710 ( .A(n_543), .B(n_417), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_555), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_598), .B(n_421), .C(n_419), .Y(n_712) );
OA22x2_ASAP7_75t_L g713 ( .A1(n_554), .A2(n_423), .B1(n_427), .B2(n_422), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_594), .B(n_10), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_597), .A2(n_429), .B1(n_431), .B2(n_428), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_555), .A2(n_305), .B(n_316), .C(n_300), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_546), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_583), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_543), .B(n_313), .Y(n_719) );
INVx1_ASAP7_75t_SL g720 ( .A(n_608), .Y(n_720) );
NAND2x1p5_ASAP7_75t_L g721 ( .A(n_563), .B(n_387), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_594), .A2(n_418), .B1(n_387), .B2(n_378), .C1(n_347), .C2(n_358), .Y(n_722) );
BUFx2_ASAP7_75t_L g723 ( .A(n_563), .Y(n_723) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_524), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_531), .Y(n_725) );
BUFx5_ASAP7_75t_L g726 ( .A(n_524), .Y(n_726) );
INVx5_ASAP7_75t_L g727 ( .A(n_524), .Y(n_727) );
BUFx2_ASAP7_75t_L g728 ( .A(n_531), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_566), .B(n_418), .Y(n_729) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_566), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_583), .Y(n_731) );
AND2x4_ASAP7_75t_SL g732 ( .A(n_581), .B(n_347), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_579), .A2(n_490), .B(n_481), .Y(n_733) );
INVx6_ASAP7_75t_L g734 ( .A(n_604), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_590), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_605), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_599), .B(n_358), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_554), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_557), .B(n_378), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_557), .Y(n_740) );
BUFx3_ASAP7_75t_L g741 ( .A(n_604), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_604), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_588), .A2(n_490), .B(n_481), .Y(n_743) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_617), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_665), .B(n_588), .Y(n_745) );
AO31x2_ASAP7_75t_L g746 ( .A1(n_716), .A2(n_466), .A3(n_450), .B(n_398), .Y(n_746) );
O2A1O1Ixp33_ASAP7_75t_L g747 ( .A1(n_628), .A2(n_463), .B(n_398), .C(n_450), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_662), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_660), .B(n_604), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_659), .B(n_10), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_654), .B(n_11), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_714), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g753 ( .A(n_645), .B(n_595), .Y(n_753) );
OAI21x1_ASAP7_75t_L g754 ( .A1(n_743), .A2(n_490), .B(n_481), .Y(n_754) );
OAI21x1_ASAP7_75t_L g755 ( .A1(n_733), .A2(n_500), .B(n_496), .Y(n_755) );
AO21x2_ASAP7_75t_L g756 ( .A1(n_623), .A2(n_466), .B(n_496), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_672), .B(n_12), .Y(n_757) );
INVx3_ASAP7_75t_L g758 ( .A(n_630), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_661), .B(n_595), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_647), .B(n_636), .Y(n_760) );
OAI21x1_ASAP7_75t_L g761 ( .A1(n_632), .A2(n_500), .B(n_496), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_737), .A2(n_595), .B(n_501), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_613), .B(n_618), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_637), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_661), .Y(n_765) );
BUFx2_ASAP7_75t_SL g766 ( .A(n_645), .Y(n_766) );
OAI21x1_ASAP7_75t_L g767 ( .A1(n_721), .A2(n_729), .B(n_612), .Y(n_767) );
INVx4_ASAP7_75t_SL g768 ( .A(n_617), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_610), .A2(n_595), .B(n_501), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_619), .A2(n_463), .B(n_466), .C(n_409), .Y(n_770) );
INVxp33_ASAP7_75t_SL g771 ( .A(n_657), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_683), .A2(n_463), .B1(n_502), .B2(n_500), .Y(n_772) );
NAND2x1p5_ASAP7_75t_L g773 ( .A(n_645), .B(n_492), .Y(n_773) );
AO21x2_ASAP7_75t_L g774 ( .A1(n_655), .A2(n_501), .B(n_486), .Y(n_774) );
AO21x2_ASAP7_75t_L g775 ( .A1(n_653), .A2(n_486), .B(n_502), .Y(n_775) );
BUFx2_ASAP7_75t_L g776 ( .A(n_614), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_638), .Y(n_777) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_667), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_SL g779 ( .A1(n_679), .A2(n_142), .B(n_290), .C(n_289), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_630), .B(n_16), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_688), .B(n_16), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_707), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_710), .A2(n_502), .B1(n_486), .B2(n_19), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g784 ( .A1(n_634), .A2(n_502), .B1(n_486), .B2(n_20), .C(n_22), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_663), .Y(n_785) );
OAI21x1_ASAP7_75t_SL g786 ( .A1(n_625), .A2(n_17), .B(n_18), .Y(n_786) );
BUFx3_ASAP7_75t_L g787 ( .A(n_614), .Y(n_787) );
AO21x2_ASAP7_75t_L g788 ( .A1(n_739), .A2(n_486), .B(n_502), .Y(n_788) );
OAI21x1_ASAP7_75t_L g789 ( .A1(n_609), .A2(n_486), .B(n_71), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_663), .B(n_492), .Y(n_790) );
INVx4_ASAP7_75t_L g791 ( .A(n_663), .Y(n_791) );
OA21x2_ASAP7_75t_L g792 ( .A1(n_609), .A2(n_486), .B(n_502), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_707), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_646), .Y(n_794) );
A2O1A1Ixp33_ASAP7_75t_L g795 ( .A1(n_698), .A2(n_492), .B(n_20), .C(n_23), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_676), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_682), .B(n_18), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_727), .B(n_23), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_624), .B(n_24), .Y(n_799) );
OAI21x1_ASAP7_75t_L g800 ( .A1(n_718), .A2(n_72), .B(n_70), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_713), .A2(n_492), .B1(n_25), .B2(n_26), .Y(n_801) );
OAI21x1_ASAP7_75t_L g802 ( .A1(n_731), .A2(n_74), .B(n_73), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_617), .Y(n_803) );
BUFx2_ASAP7_75t_L g804 ( .A(n_620), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_621), .Y(n_805) );
OAI21x1_ASAP7_75t_L g806 ( .A1(n_735), .A2(n_80), .B(n_78), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g807 ( .A1(n_705), .A2(n_24), .B1(n_28), .B2(n_29), .C(n_30), .Y(n_807) );
INVx2_ASAP7_75t_SL g808 ( .A(n_644), .Y(n_808) );
INVx4_ASAP7_75t_L g809 ( .A(n_727), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_693), .Y(n_810) );
BUFx6f_ASAP7_75t_L g811 ( .A(n_684), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_611), .A2(n_84), .B(n_82), .Y(n_812) );
INVx4_ASAP7_75t_L g813 ( .A(n_727), .Y(n_813) );
NOR2xp33_ASAP7_75t_SL g814 ( .A(n_652), .B(n_28), .Y(n_814) );
AO21x2_ASAP7_75t_L g815 ( .A1(n_706), .A2(n_88), .B(n_87), .Y(n_815) );
OAI21x1_ASAP7_75t_L g816 ( .A1(n_615), .A2(n_95), .B(n_93), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_658), .Y(n_817) );
NOR2xp33_ASAP7_75t_SL g818 ( .A(n_669), .B(n_29), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_712), .A2(n_492), .B1(n_32), .B2(n_33), .Y(n_819) );
INVx3_ASAP7_75t_L g820 ( .A(n_641), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_616), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_821) );
NOR2xp67_ASAP7_75t_L g822 ( .A(n_633), .B(n_34), .Y(n_822) );
OAI22xp5_ASAP7_75t_SL g823 ( .A1(n_668), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_694), .Y(n_824) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_667), .A2(n_36), .B1(n_37), .B2(n_39), .Y(n_825) );
AO21x2_ASAP7_75t_L g826 ( .A1(n_643), .A2(n_100), .B(n_99), .Y(n_826) );
OA21x2_ASAP7_75t_L g827 ( .A1(n_675), .A2(n_492), .B(n_102), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_627), .B(n_37), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_696), .B(n_40), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_626), .B(n_40), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_629), .Y(n_831) );
AOI21xp5_ASAP7_75t_L g832 ( .A1(n_738), .A2(n_492), .B(n_169), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_691), .A2(n_492), .B1(n_42), .B2(n_43), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_656), .A2(n_41), .B1(n_42), .B2(n_44), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_670), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_664), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_671), .B(n_41), .Y(n_837) );
OAI21x1_ASAP7_75t_L g838 ( .A1(n_674), .A2(n_171), .B(n_286), .Y(n_838) );
INVx1_ASAP7_75t_SL g839 ( .A(n_620), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_690), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_651), .B(n_44), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g842 ( .A(n_635), .Y(n_842) );
OAI21x1_ASAP7_75t_L g843 ( .A1(n_680), .A2(n_170), .B(n_283), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_687), .B(n_45), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_649), .B(n_46), .Y(n_845) );
INVx1_ASAP7_75t_SL g846 ( .A(n_650), .Y(n_846) );
OAI21x1_ASAP7_75t_L g847 ( .A1(n_641), .A2(n_175), .B(n_280), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_651), .B(n_47), .Y(n_848) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_730), .Y(n_849) );
OA21x2_ASAP7_75t_L g850 ( .A1(n_689), .A2(n_179), .B(n_278), .Y(n_850) );
OAI21x1_ASAP7_75t_L g851 ( .A1(n_673), .A2(n_699), .B(n_736), .Y(n_851) );
OA21x2_ASAP7_75t_L g852 ( .A1(n_709), .A2(n_167), .B(n_277), .Y(n_852) );
BUFx3_ASAP7_75t_L g853 ( .A(n_741), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_710), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_656), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_673), .A2(n_166), .B(n_276), .Y(n_856) );
O2A1O1Ixp33_ASAP7_75t_L g857 ( .A1(n_708), .A2(n_48), .B(n_49), .C(n_50), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_640), .B(n_49), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_711), .B(n_51), .Y(n_859) );
NAND2xp33_ASAP7_75t_SL g860 ( .A(n_724), .B(n_52), .Y(n_860) );
OAI21x1_ASAP7_75t_L g861 ( .A1(n_699), .A2(n_183), .B(n_274), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_703), .A2(n_181), .B(n_273), .Y(n_862) );
INVx3_ASAP7_75t_L g863 ( .A(n_684), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_639), .B(n_52), .Y(n_864) );
OR2x6_ASAP7_75t_L g865 ( .A(n_622), .B(n_54), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_677), .B(n_54), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_704), .Y(n_867) );
AND2x4_ASAP7_75t_L g868 ( .A(n_678), .B(n_55), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_692), .B(n_56), .Y(n_869) );
OR2x6_ASAP7_75t_L g870 ( .A(n_622), .B(n_56), .Y(n_870) );
AND2x4_ASAP7_75t_L g871 ( .A(n_678), .B(n_57), .Y(n_871) );
OA21x2_ASAP7_75t_L g872 ( .A1(n_666), .A2(n_719), .B(n_715), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_717), .Y(n_873) );
OA21x2_ASAP7_75t_L g874 ( .A1(n_719), .A2(n_186), .B(n_272), .Y(n_874) );
AO31x2_ASAP7_75t_L g875 ( .A1(n_702), .A2(n_57), .A3(n_58), .B(n_59), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_725), .Y(n_876) );
OAI21x1_ASAP7_75t_L g877 ( .A1(n_631), .A2(n_185), .B(n_269), .Y(n_877) );
OAI21x1_ASAP7_75t_L g878 ( .A1(n_742), .A2(n_164), .B(n_267), .Y(n_878) );
NAND2xp33_ASAP7_75t_R g879 ( .A(n_740), .B(n_58), .Y(n_879) );
INVx2_ASAP7_75t_SL g880 ( .A(n_732), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_686), .A2(n_187), .B(n_265), .Y(n_881) );
BUFx2_ASAP7_75t_L g882 ( .A(n_684), .Y(n_882) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_730), .Y(n_883) );
AO21x1_ASAP7_75t_L g884 ( .A1(n_695), .A2(n_163), .B(n_264), .Y(n_884) );
OR2x2_ASAP7_75t_L g885 ( .A(n_648), .B(n_59), .Y(n_885) );
OAI21x1_ASAP7_75t_L g886 ( .A1(n_700), .A2(n_161), .B(n_261), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_685), .B(n_60), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_722), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_728), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_864), .B(n_642), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_751), .A2(n_681), .B1(n_720), .B2(n_726), .Y(n_891) );
OAI21x1_ASAP7_75t_SL g892 ( .A1(n_749), .A2(n_701), .B(n_726), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_829), .Y(n_893) );
OR2x2_ASAP7_75t_L g894 ( .A(n_748), .B(n_854), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_763), .A2(n_697), .B1(n_723), .B2(n_701), .C(n_730), .Y(n_895) );
INVx3_ASAP7_75t_L g896 ( .A(n_791), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_829), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_751), .A2(n_726), .B1(n_734), .B2(n_63), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_830), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_765), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_805), .B(n_61), .Y(n_901) );
OAI211xp5_ASAP7_75t_L g902 ( .A1(n_833), .A2(n_726), .B(n_64), .C(n_65), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_787), .Y(n_903) );
OAI21x1_ASAP7_75t_L g904 ( .A1(n_754), .A2(n_726), .B(n_734), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_750), .A2(n_62), .B1(n_67), .B2(n_69), .Y(n_905) );
OAI21xp5_ASAP7_75t_L g906 ( .A1(n_750), .A2(n_67), .B(n_69), .Y(n_906) );
OR2x2_ASAP7_75t_L g907 ( .A(n_776), .B(n_101), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_830), .Y(n_908) );
OAI211xp5_ASAP7_75t_SL g909 ( .A1(n_807), .A2(n_105), .B(n_106), .C(n_107), .Y(n_909) );
OR2x2_ASAP7_75t_L g910 ( .A(n_760), .B(n_108), .Y(n_910) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_865), .A2(n_109), .B1(n_110), .B2(n_112), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_866), .B(n_113), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_752), .A2(n_115), .B1(n_116), .B2(n_120), .Y(n_913) );
AOI222xp33_ASAP7_75t_L g914 ( .A1(n_845), .A2(n_823), .B1(n_807), .B2(n_841), .C1(n_848), .C2(n_828), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_749), .A2(n_124), .B(n_125), .Y(n_915) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_771), .A2(n_127), .B1(n_130), .B2(n_132), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_837), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_837), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_865), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_762), .A2(n_140), .B(n_143), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_865), .A2(n_144), .B1(n_145), .B2(n_149), .Y(n_921) );
A2O1A1Ixp33_ASAP7_75t_L g922 ( .A1(n_747), .A2(n_150), .B(n_151), .C(n_154), .Y(n_922) );
A2O1A1Ixp33_ASAP7_75t_L g923 ( .A1(n_747), .A2(n_155), .B(n_157), .C(n_158), .Y(n_923) );
OAI222xp33_ASAP7_75t_L g924 ( .A1(n_870), .A2(n_159), .B1(n_188), .B2(n_189), .C1(n_190), .C2(n_193), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_844), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g926 ( .A1(n_762), .A2(n_194), .B(n_195), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_781), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_888), .A2(n_204), .B1(n_205), .B2(n_209), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_870), .A2(n_210), .B1(n_211), .B2(n_213), .Y(n_929) );
AOI22xp33_ASAP7_75t_SL g930 ( .A1(n_870), .A2(n_220), .B1(n_222), .B2(n_223), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_888), .A2(n_872), .B1(n_869), .B2(n_885), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_855), .B(n_288), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_845), .A2(n_887), .B1(n_784), .B2(n_872), .Y(n_933) );
OAI21xp5_ASAP7_75t_SL g934 ( .A1(n_778), .A2(n_224), .B(n_225), .Y(n_934) );
AOI21xp33_ASAP7_75t_L g935 ( .A1(n_869), .A2(n_226), .B(n_227), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_810), .B(n_229), .Y(n_936) );
AOI21xp5_ASAP7_75t_L g937 ( .A1(n_769), .A2(n_232), .B(n_234), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_784), .A2(n_235), .B1(n_237), .B2(n_238), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_769), .A2(n_240), .B(n_241), .Y(n_939) );
BUFx2_ASAP7_75t_L g940 ( .A(n_785), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_781), .A2(n_243), .B1(n_244), .B2(n_247), .C(n_248), .Y(n_941) );
AO21x1_ASAP7_75t_L g942 ( .A1(n_783), .A2(n_250), .B(n_253), .Y(n_942) );
AOI21xp5_ASAP7_75t_L g943 ( .A1(n_759), .A2(n_256), .B(n_257), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_844), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_873), .Y(n_945) );
NAND4xp25_ASAP7_75t_L g946 ( .A(n_818), .B(n_799), .C(n_879), .D(n_797), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_824), .B(n_831), .Y(n_947) );
INVx2_ASAP7_75t_L g948 ( .A(n_836), .Y(n_948) );
AOI21x1_ASAP7_75t_L g949 ( .A1(n_827), .A2(n_852), .B(n_884), .Y(n_949) );
OAI21x1_ASAP7_75t_L g950 ( .A1(n_755), .A2(n_789), .B(n_761), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_764), .Y(n_951) );
OA21x2_ASAP7_75t_L g952 ( .A1(n_881), .A2(n_886), .B(n_832), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_778), .A2(n_825), .B1(n_757), .B2(n_858), .Y(n_953) );
AND2x4_ASAP7_75t_L g954 ( .A(n_768), .B(n_791), .Y(n_954) );
OAI21xp5_ASAP7_75t_L g955 ( .A1(n_745), .A2(n_858), .B(n_770), .Y(n_955) );
A2O1A1Ixp33_ASAP7_75t_L g956 ( .A1(n_857), .A2(n_795), .B(n_757), .C(n_860), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_825), .A2(n_834), .B1(n_871), .B2(n_868), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_879), .A2(n_868), .B1(n_871), .B2(n_797), .Y(n_958) );
AND2x4_ASAP7_75t_L g959 ( .A(n_768), .B(n_758), .Y(n_959) );
OAI22xp5_ASAP7_75t_SL g960 ( .A1(n_842), .A2(n_821), .B1(n_880), .B2(n_834), .Y(n_960) );
AO21x2_ASAP7_75t_L g961 ( .A1(n_756), .A2(n_770), .B(n_775), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_859), .Y(n_962) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_832), .A2(n_812), .B(n_816), .Y(n_963) );
OAI22xp33_ASAP7_75t_SL g964 ( .A1(n_814), .A2(n_783), .B1(n_780), .B2(n_798), .Y(n_964) );
AOI22xp33_ASAP7_75t_SL g965 ( .A1(n_780), .A2(n_786), .B1(n_798), .B2(n_766), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_801), .A2(n_782), .B1(n_793), .B2(n_821), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_801), .A2(n_822), .B1(n_859), .B2(n_889), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_785), .Y(n_968) );
OR2x2_ASAP7_75t_L g969 ( .A(n_846), .B(n_853), .Y(n_969) );
AOI222xp33_ASAP7_75t_L g970 ( .A1(n_839), .A2(n_804), .B1(n_796), .B2(n_808), .C1(n_795), .C2(n_819), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_875), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_882), .B(n_817), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_777), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_819), .A2(n_775), .B1(n_756), .B2(n_774), .Y(n_974) );
OAI21x1_ASAP7_75t_L g975 ( .A1(n_851), .A2(n_767), .B(n_792), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_803), .B(n_863), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_774), .A2(n_758), .B1(n_815), .B2(n_876), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_875), .Y(n_978) );
OA21x2_ASAP7_75t_L g979 ( .A1(n_838), .A2(n_843), .B(n_802), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_820), .B(n_809), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_794), .B(n_840), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_875), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_759), .A2(n_835), .B1(n_867), .B2(n_857), .Y(n_983) );
NAND2xp33_ASAP7_75t_L g984 ( .A(n_744), .B(n_811), .Y(n_984) );
AOI222xp33_ASAP7_75t_L g985 ( .A1(n_820), .A2(n_813), .B1(n_809), .B2(n_803), .C1(n_768), .C2(n_863), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_744), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_811), .B(n_744), .Y(n_987) );
BUFx4f_ASAP7_75t_SL g988 ( .A(n_811), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_875), .Y(n_989) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_744), .Y(n_990) );
NOR2x1_ASAP7_75t_SL g991 ( .A(n_813), .B(n_883), .Y(n_991) );
INVx3_ASAP7_75t_L g992 ( .A(n_773), .Y(n_992) );
OAI21x1_ASAP7_75t_L g993 ( .A1(n_792), .A2(n_800), .B(n_806), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_815), .A2(n_826), .B1(n_850), .B2(n_827), .Y(n_994) );
CKINVDCx11_ASAP7_75t_R g995 ( .A(n_849), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_826), .A2(n_850), .B1(n_874), .B2(n_772), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_790), .B(n_773), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_790), .B(n_772), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g999 ( .A1(n_874), .A2(n_852), .B1(n_878), .B2(n_847), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_753), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_753), .B(n_746), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_746), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_746), .B(n_883), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_746), .Y(n_1004) );
AOI21xp5_ASAP7_75t_L g1005 ( .A1(n_788), .A2(n_779), .B(n_862), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_849), .B(n_883), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_788), .Y(n_1007) );
OA21x2_ASAP7_75t_L g1008 ( .A1(n_856), .A2(n_861), .B(n_862), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_849), .A2(n_883), .B1(n_877), .B2(n_779), .Y(n_1009) );
O2A1O1Ixp33_ASAP7_75t_SL g1010 ( .A1(n_849), .A2(n_749), .B(n_795), .C(n_770), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_864), .B(n_535), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_829), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_785), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1014 ( .A1(n_763), .A2(n_624), .B1(n_535), .B2(n_479), .C(n_528), .Y(n_1014) );
INVx2_ASAP7_75t_L g1015 ( .A(n_765), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1016 ( .A(n_768), .B(n_645), .Y(n_1016) );
OR2x6_ASAP7_75t_L g1017 ( .A(n_766), .B(n_776), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_864), .B(n_535), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_829), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_971), .Y(n_1020) );
NAND2xp33_ASAP7_75t_SL g1021 ( .A(n_957), .B(n_960), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_890), .B(n_1011), .Y(n_1022) );
INVx4_ASAP7_75t_L g1023 ( .A(n_988), .Y(n_1023) );
OAI211xp5_ASAP7_75t_L g1024 ( .A1(n_958), .A2(n_914), .B(n_946), .C(n_957), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_978), .Y(n_1025) );
AND2x4_ASAP7_75t_SL g1026 ( .A(n_1017), .B(n_997), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_1013), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_1013), .B(n_940), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_982), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_951), .B(n_973), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_989), .Y(n_1031) );
OAI221xp5_ASAP7_75t_SL g1032 ( .A1(n_1014), .A2(n_953), .B1(n_966), .B2(n_898), .C(n_891), .Y(n_1032) );
BUFx2_ASAP7_75t_L g1033 ( .A(n_1001), .Y(n_1033) );
INVx3_ASAP7_75t_L g1034 ( .A(n_1016), .Y(n_1034) );
BUFx3_ASAP7_75t_L g1035 ( .A(n_988), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_900), .B(n_1015), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_1006), .B(n_1003), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_962), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_945), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_893), .B(n_1019), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_897), .B(n_899), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_908), .Y(n_1042) );
INVx2_ASAP7_75t_L g1043 ( .A(n_975), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_953), .A2(n_1018), .B1(n_966), .B2(n_898), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_917), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_947), .B(n_948), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1047 ( .A(n_970), .B(n_905), .C(n_967), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_1002), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_918), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_925), .Y(n_1050) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_931), .A2(n_933), .B1(n_944), .B2(n_1012), .C(n_967), .Y(n_1051) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1004), .Y(n_1052) );
BUFx3_ASAP7_75t_L g1053 ( .A(n_995), .Y(n_1053) );
INVxp67_ASAP7_75t_L g1054 ( .A(n_1017), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_891), .B(n_933), .Y(n_1055) );
AOI21xp5_ASAP7_75t_L g1056 ( .A1(n_1005), .A2(n_999), .B(n_994), .Y(n_1056) );
AND2x4_ASAP7_75t_L g1057 ( .A(n_986), .B(n_1000), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_968), .B(n_894), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_981), .B(n_976), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_964), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1061 ( .A(n_972), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_896), .B(n_992), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_990), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_990), .Y(n_1064) );
INVx2_ASAP7_75t_SL g1065 ( .A(n_1017), .Y(n_1065) );
NOR2x1_ASAP7_75t_L g1066 ( .A(n_911), .B(n_934), .Y(n_1066) );
INVx2_ASAP7_75t_L g1067 ( .A(n_993), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_906), .B(n_992), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_950), .Y(n_1069) );
INVx2_ASAP7_75t_L g1070 ( .A(n_961), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_896), .B(n_905), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_969), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_987), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_959), .B(n_954), .Y(n_1074) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_998), .Y(n_1075) );
INVx3_ASAP7_75t_L g1076 ( .A(n_1016), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_910), .B(n_956), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1078 ( .A1(n_895), .A2(n_983), .B1(n_902), .B2(n_911), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_959), .B(n_954), .Y(n_1079) );
AOI222xp33_ASAP7_75t_L g1080 ( .A1(n_912), .A2(n_924), .B1(n_929), .B2(n_919), .C1(n_921), .C2(n_909), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g1081 ( .A(n_901), .Y(n_1081) );
OR2x2_ASAP7_75t_L g1082 ( .A(n_955), .B(n_961), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_936), .Y(n_1083) );
NOR2xp33_ASAP7_75t_L g1084 ( .A(n_903), .B(n_907), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1085 ( .A(n_974), .B(n_980), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_965), .B(n_930), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1087 ( .A(n_965), .B(n_930), .Y(n_1087) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_991), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_985), .B(n_929), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_904), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_919), .B(n_921), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1092 ( .A(n_920), .B(n_926), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_916), .B(n_938), .Y(n_1093) );
AND2x4_ASAP7_75t_SL g1094 ( .A(n_913), .B(n_927), .Y(n_1094) );
BUFx3_ASAP7_75t_L g1095 ( .A(n_892), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_916), .B(n_938), .Y(n_1096) );
INVxp67_ASAP7_75t_L g1097 ( .A(n_932), .Y(n_1097) );
INVx3_ASAP7_75t_L g1098 ( .A(n_1008), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_913), .B(n_974), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g1100 ( .A(n_924), .Y(n_1100) );
INVx3_ASAP7_75t_L g1101 ( .A(n_1008), .Y(n_1101) );
OAI31xp33_ASAP7_75t_L g1102 ( .A1(n_909), .A2(n_928), .A3(n_941), .B(n_1010), .Y(n_1102) );
OAI21x1_ASAP7_75t_L g1103 ( .A1(n_949), .A2(n_1009), .B(n_994), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g1104 ( .A(n_984), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_977), .B(n_942), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_979), .Y(n_1106) );
BUFx2_ASAP7_75t_L g1107 ( .A(n_979), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_943), .Y(n_1108) );
AND2x4_ASAP7_75t_L g1109 ( .A(n_1009), .B(n_939), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_977), .B(n_996), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_996), .B(n_922), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_915), .B(n_999), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_923), .B(n_952), .Y(n_1113) );
INVx2_ASAP7_75t_SL g1114 ( .A(n_952), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_935), .B(n_937), .Y(n_1115) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_963), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_963), .B(n_951), .Y(n_1117) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1007), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_971), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_1013), .Y(n_1120) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_1014), .A2(n_493), .B1(n_634), .B2(n_890), .C(n_1011), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_1028), .Y(n_1122) );
INVx3_ASAP7_75t_L g1123 ( .A(n_1095), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1033), .B(n_1037), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g1125 ( .A1(n_1024), .A2(n_1087), .B1(n_1086), .B2(n_1100), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1126 ( .A(n_1028), .Y(n_1126) );
INVxp67_ASAP7_75t_SL g1127 ( .A(n_1033), .Y(n_1127) );
AO221x2_ASAP7_75t_L g1128 ( .A1(n_1047), .A2(n_1021), .B1(n_1055), .B2(n_1045), .C(n_1042), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1020), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_1027), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1020), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1037), .B(n_1059), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1040), .B(n_1041), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1025), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1106), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1025), .Y(n_1136) );
INVx3_ASAP7_75t_L g1137 ( .A(n_1095), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1029), .Y(n_1138) );
AOI221xp5_ASAP7_75t_L g1139 ( .A1(n_1121), .A2(n_1044), .B1(n_1032), .B2(n_1022), .C(n_1051), .Y(n_1139) );
INVx2_ASAP7_75t_SL g1140 ( .A(n_1026), .Y(n_1140) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1106), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1142 ( .A(n_1120), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1037), .B(n_1059), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1037), .B(n_1029), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1031), .B(n_1119), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1085), .B(n_1075), .Y(n_1146) );
NAND2x1p5_ASAP7_75t_L g1147 ( .A(n_1034), .B(n_1076), .Y(n_1147) );
BUFx3_ASAP7_75t_L g1148 ( .A(n_1026), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1031), .B(n_1119), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1040), .B(n_1041), .Y(n_1150) );
BUFx6f_ASAP7_75t_L g1151 ( .A(n_1098), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1085), .B(n_1075), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1036), .B(n_1110), .Y(n_1153) );
OAI211xp5_ASAP7_75t_SL g1154 ( .A1(n_1054), .A2(n_1058), .B(n_1081), .C(n_1039), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1036), .B(n_1110), .Y(n_1155) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_1086), .A2(n_1087), .B1(n_1066), .B2(n_1089), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1039), .B(n_1073), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1117), .Y(n_1158) );
INVx2_ASAP7_75t_SL g1159 ( .A(n_1065), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1073), .B(n_1030), .Y(n_1160) );
AOI21xp33_ASAP7_75t_L g1161 ( .A1(n_1080), .A2(n_1089), .B(n_1066), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1162 ( .A(n_1117), .B(n_1052), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1030), .B(n_1063), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1063), .B(n_1064), .Y(n_1164) );
BUFx3_ASAP7_75t_L g1165 ( .A(n_1034), .Y(n_1165) );
INVx1_ASAP7_75t_SL g1166 ( .A(n_1053), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1064), .B(n_1050), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1038), .B(n_1050), .Y(n_1168) );
HB1xp67_ASAP7_75t_L g1169 ( .A(n_1072), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1038), .B(n_1049), .Y(n_1170) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_1118), .Y(n_1171) );
BUFx2_ASAP7_75t_L g1172 ( .A(n_1088), .Y(n_1172) );
NAND4xp25_ASAP7_75t_L g1173 ( .A(n_1077), .B(n_1078), .C(n_1049), .D(n_1045), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1042), .B(n_1052), .Y(n_1174) );
INVxp67_ASAP7_75t_L g1175 ( .A(n_1084), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1048), .B(n_1105), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_1061), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1105), .B(n_1099), .Y(n_1178) );
AOI221xp5_ASAP7_75t_L g1179 ( .A1(n_1060), .A2(n_1046), .B1(n_1077), .B2(n_1071), .C(n_1097), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1068), .B(n_1071), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1082), .B(n_1065), .Y(n_1181) );
OAI21xp33_ASAP7_75t_L g1182 ( .A1(n_1078), .A2(n_1093), .B(n_1096), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1068), .B(n_1074), .Y(n_1183) );
AND2x4_ASAP7_75t_L g1184 ( .A(n_1114), .B(n_1116), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1099), .B(n_1082), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1057), .B(n_1079), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1057), .B(n_1079), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1057), .B(n_1074), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1114), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1107), .Y(n_1190) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_1062), .Y(n_1191) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1098), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1057), .B(n_1111), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1062), .B(n_1034), .Y(n_1194) );
AND2x4_ASAP7_75t_L g1195 ( .A(n_1116), .B(n_1101), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1107), .Y(n_1196) );
INVxp33_ASAP7_75t_L g1197 ( .A(n_1035), .Y(n_1197) );
A2O1A1Ixp33_ASAP7_75t_L g1198 ( .A1(n_1093), .A2(n_1096), .B(n_1102), .C(n_1094), .Y(n_1198) );
BUFx2_ASAP7_75t_L g1199 ( .A(n_1104), .Y(n_1199) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_1083), .A2(n_1091), .B1(n_1056), .B2(n_1070), .C(n_1112), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1160), .B(n_1091), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1153), .B(n_1070), .Y(n_1202) );
INVx1_ASAP7_75t_SL g1203 ( .A(n_1166), .Y(n_1203) );
INVxp67_ASAP7_75t_SL g1204 ( .A(n_1177), .Y(n_1204) );
OAI31xp33_ASAP7_75t_L g1205 ( .A1(n_1198), .A2(n_1094), .A3(n_1035), .B(n_1053), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1146), .B(n_1101), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1146), .B(n_1103), .Y(n_1207) );
HB1xp67_ASAP7_75t_L g1208 ( .A(n_1172), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1153), .B(n_1111), .Y(n_1209) );
HB1xp67_ASAP7_75t_L g1210 ( .A(n_1172), .Y(n_1210) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1135), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_1156), .A2(n_1076), .B1(n_1023), .B2(n_1083), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1155), .B(n_1113), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1129), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1160), .B(n_1076), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1155), .B(n_1113), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1133), .B(n_1023), .Y(n_1217) );
BUFx3_ASAP7_75t_L g1218 ( .A(n_1148), .Y(n_1218) );
NOR3x1_ASAP7_75t_L g1219 ( .A(n_1140), .B(n_1115), .C(n_1023), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1185), .B(n_1043), .Y(n_1220) );
AND2x4_ASAP7_75t_L g1221 ( .A(n_1158), .B(n_1067), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1150), .B(n_1108), .Y(n_1222) );
NAND4xp25_ASAP7_75t_L g1223 ( .A(n_1161), .B(n_1139), .C(n_1125), .D(n_1156), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1131), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1185), .B(n_1043), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1152), .B(n_1069), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1178), .B(n_1069), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1178), .B(n_1067), .Y(n_1228) );
INVx1_ASAP7_75t_SL g1229 ( .A(n_1169), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1152), .B(n_1090), .Y(n_1230) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_1127), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1144), .B(n_1090), .Y(n_1232) );
NOR2xp33_ASAP7_75t_L g1233 ( .A(n_1175), .B(n_1092), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1144), .B(n_1176), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1176), .B(n_1109), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1131), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1158), .B(n_1109), .Y(n_1237) );
BUFx2_ASAP7_75t_L g1238 ( .A(n_1123), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1134), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1193), .B(n_1109), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1134), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1193), .B(n_1109), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1136), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1180), .B(n_1092), .Y(n_1244) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_1182), .A2(n_1092), .B1(n_1128), .B2(n_1179), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1136), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1163), .B(n_1092), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1132), .B(n_1143), .Y(n_1248) );
NAND2xp33_ASAP7_75t_SL g1249 ( .A(n_1140), .B(n_1124), .Y(n_1249) );
OAI33xp33_ASAP7_75t_L g1250 ( .A1(n_1182), .A2(n_1154), .A3(n_1173), .B1(n_1183), .B2(n_1138), .B3(n_1164), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1122), .B(n_1126), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1132), .B(n_1143), .Y(n_1252) );
BUFx2_ASAP7_75t_L g1253 ( .A(n_1123), .Y(n_1253) );
CKINVDCx16_ASAP7_75t_R g1254 ( .A(n_1148), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1163), .B(n_1157), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1138), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1162), .B(n_1149), .Y(n_1257) );
INVx4_ASAP7_75t_L g1258 ( .A(n_1148), .Y(n_1258) );
NAND3xp33_ASAP7_75t_SL g1259 ( .A(n_1197), .B(n_1142), .C(n_1130), .Y(n_1259) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1141), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1157), .B(n_1170), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1181), .B(n_1164), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1251), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1204), .Y(n_1264) );
NOR2xp33_ASAP7_75t_L g1265 ( .A(n_1223), .B(n_1250), .Y(n_1265) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1211), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1209), .B(n_1128), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1257), .B(n_1162), .Y(n_1268) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_1208), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1255), .B(n_1124), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1271 ( .A(n_1210), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1262), .B(n_1181), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1209), .B(n_1128), .Y(n_1273) );
AND2x4_ASAP7_75t_L g1274 ( .A(n_1257), .B(n_1123), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1262), .B(n_1171), .Y(n_1275) );
NOR2xp33_ASAP7_75t_R g1276 ( .A(n_1249), .B(n_1123), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1248), .B(n_1187), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1214), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1201), .B(n_1128), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g1280 ( .A(n_1231), .Y(n_1280) );
INVx2_ASAP7_75t_L g1281 ( .A(n_1211), .Y(n_1281) );
AOI22xp5_ASAP7_75t_L g1282 ( .A1(n_1223), .A2(n_1173), .B1(n_1187), .B2(n_1186), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1224), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1229), .B(n_1167), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1234), .B(n_1162), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1261), .B(n_1167), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1234), .B(n_1168), .Y(n_1287) );
INVx2_ASAP7_75t_SL g1288 ( .A(n_1254), .Y(n_1288) );
HB1xp67_ASAP7_75t_L g1289 ( .A(n_1231), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1248), .B(n_1168), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1236), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1239), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1252), .B(n_1170), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1239), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1252), .B(n_1188), .Y(n_1295) );
INVxp67_ASAP7_75t_L g1296 ( .A(n_1259), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1228), .B(n_1149), .Y(n_1297) );
NOR2x1_ASAP7_75t_L g1298 ( .A(n_1258), .B(n_1137), .Y(n_1298) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_1237), .B(n_1137), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g1300 ( .A(n_1219), .Y(n_1300) );
AND2x4_ASAP7_75t_L g1301 ( .A(n_1237), .B(n_1137), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1264), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1287), .B(n_1290), .Y(n_1303) );
AOI22xp5_ASAP7_75t_L g1304 ( .A1(n_1265), .A2(n_1233), .B1(n_1212), .B2(n_1245), .Y(n_1304) );
AOI211xp5_ASAP7_75t_L g1305 ( .A1(n_1265), .A2(n_1205), .B(n_1203), .C(n_1244), .Y(n_1305) );
NAND4xp25_ASAP7_75t_L g1306 ( .A(n_1282), .B(n_1205), .C(n_1219), .D(n_1217), .Y(n_1306) );
INVx2_ASAP7_75t_SL g1307 ( .A(n_1276), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1263), .B(n_1213), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1279), .B(n_1213), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1267), .B(n_1216), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_1273), .A2(n_1244), .B1(n_1188), .B2(n_1186), .Y(n_1311) );
OAI221xp5_ASAP7_75t_SL g1312 ( .A1(n_1296), .A2(n_1247), .B1(n_1215), .B2(n_1218), .C(n_1207), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1272), .Y(n_1313) );
OAI332xp33_ASAP7_75t_L g1314 ( .A1(n_1300), .A2(n_1254), .A3(n_1222), .B1(n_1207), .B2(n_1206), .B3(n_1256), .C1(n_1241), .C2(n_1246), .Y(n_1314) );
AOI322xp5_ASAP7_75t_L g1315 ( .A1(n_1288), .A2(n_1216), .A3(n_1235), .B1(n_1240), .B2(n_1242), .C1(n_1227), .C2(n_1228), .Y(n_1315) );
INVx4_ASAP7_75t_L g1316 ( .A(n_1288), .Y(n_1316) );
AOI322xp5_ASAP7_75t_L g1317 ( .A1(n_1293), .A2(n_1235), .A3(n_1240), .B1(n_1242), .B2(n_1227), .C1(n_1202), .C2(n_1200), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1275), .Y(n_1318) );
INVx1_ASAP7_75t_SL g1319 ( .A(n_1276), .Y(n_1319) );
INVxp67_ASAP7_75t_SL g1320 ( .A(n_1280), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1297), .B(n_1202), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1285), .B(n_1220), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1285), .B(n_1220), .Y(n_1323) );
AOI222xp33_ASAP7_75t_L g1324 ( .A1(n_1284), .A2(n_1225), .B1(n_1246), .B2(n_1256), .C1(n_1241), .C2(n_1243), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1325 ( .A(n_1270), .B(n_1206), .Y(n_1325) );
O2A1O1Ixp33_ASAP7_75t_L g1326 ( .A1(n_1280), .A2(n_1159), .B(n_1191), .C(n_1199), .Y(n_1326) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_1289), .A2(n_1243), .B1(n_1225), .B2(n_1145), .C(n_1238), .Y(n_1327) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1286), .B(n_1145), .Y(n_1328) );
OAI21xp33_ASAP7_75t_L g1329 ( .A1(n_1289), .A2(n_1232), .B(n_1226), .Y(n_1329) );
XNOR2xp5_ASAP7_75t_L g1330 ( .A(n_1305), .B(n_1277), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_1306), .A2(n_1274), .B1(n_1299), .B2(n_1301), .Y(n_1331) );
OAI221xp5_ASAP7_75t_L g1332 ( .A1(n_1304), .A2(n_1269), .B1(n_1271), .B2(n_1298), .C(n_1253), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1324), .B(n_1269), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1302), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1325), .Y(n_1335) );
XOR2x2_ASAP7_75t_L g1336 ( .A(n_1316), .B(n_1258), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g1337 ( .A1(n_1307), .A2(n_1258), .B1(n_1274), .B2(n_1218), .Y(n_1337) );
AOI21xp33_ASAP7_75t_L g1338 ( .A1(n_1326), .A2(n_1271), .B(n_1159), .Y(n_1338) );
NAND2xp5_ASAP7_75t_SL g1339 ( .A(n_1307), .B(n_1258), .Y(n_1339) );
NAND2xp5_ASAP7_75t_SL g1340 ( .A(n_1319), .B(n_1218), .Y(n_1340) );
CKINVDCx20_ASAP7_75t_R g1341 ( .A(n_1316), .Y(n_1341) );
OAI21xp33_ASAP7_75t_L g1342 ( .A1(n_1315), .A2(n_1274), .B(n_1268), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1318), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1322), .B(n_1295), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1323), .B(n_1268), .Y(n_1345) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1320), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1313), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1348 ( .A(n_1333), .B(n_1314), .Y(n_1348) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_1341), .A2(n_1316), .B1(n_1312), .B2(n_1311), .Y(n_1349) );
INVx1_ASAP7_75t_SL g1350 ( .A(n_1341), .Y(n_1350) );
XNOR2x1_ASAP7_75t_L g1351 ( .A(n_1330), .B(n_1303), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_1342), .A2(n_1311), .B1(n_1309), .B2(n_1327), .Y(n_1352) );
OA21x2_ASAP7_75t_L g1353 ( .A1(n_1346), .A2(n_1320), .B(n_1329), .Y(n_1353) );
O2A1O1Ixp33_ASAP7_75t_L g1354 ( .A1(n_1332), .A2(n_1312), .B(n_1310), .C(n_1308), .Y(n_1354) );
OAI222xp33_ASAP7_75t_L g1355 ( .A1(n_1331), .A2(n_1339), .B1(n_1340), .B2(n_1337), .C1(n_1335), .C2(n_1347), .Y(n_1355) );
AOI221xp5_ASAP7_75t_SL g1356 ( .A1(n_1340), .A2(n_1321), .B1(n_1328), .B2(n_1317), .C(n_1294), .Y(n_1356) );
OAI221xp5_ASAP7_75t_L g1357 ( .A1(n_1339), .A2(n_1253), .B1(n_1238), .B2(n_1278), .C(n_1291), .Y(n_1357) );
OR2x2_ASAP7_75t_L g1358 ( .A(n_1343), .B(n_1226), .Y(n_1358) );
AOI211xp5_ASAP7_75t_L g1359 ( .A1(n_1355), .A2(n_1338), .B(n_1334), .C(n_1336), .Y(n_1359) );
OAI22xp33_ASAP7_75t_L g1360 ( .A1(n_1349), .A2(n_1336), .B1(n_1137), .B2(n_1345), .Y(n_1360) );
AOI321xp33_ASAP7_75t_L g1361 ( .A1(n_1348), .A2(n_1299), .A3(n_1301), .B1(n_1345), .B2(n_1344), .C(n_1283), .Y(n_1361) );
NOR3xp33_ASAP7_75t_L g1362 ( .A(n_1356), .B(n_1199), .C(n_1292), .Y(n_1362) );
AOI211xp5_ASAP7_75t_SL g1363 ( .A1(n_1357), .A2(n_1301), .B(n_1299), .C(n_1194), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1358), .Y(n_1364) );
OR2x2_ASAP7_75t_L g1365 ( .A(n_1364), .B(n_1352), .Y(n_1365) );
BUFx6f_ASAP7_75t_L g1366 ( .A(n_1359), .Y(n_1366) );
AOI22xp5_ASAP7_75t_SL g1367 ( .A1(n_1361), .A2(n_1350), .B1(n_1353), .B2(n_1351), .Y(n_1367) );
AOI21xp33_ASAP7_75t_L g1368 ( .A1(n_1360), .A2(n_1354), .B(n_1353), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_1367), .A2(n_1353), .B1(n_1362), .B2(n_1363), .Y(n_1369) );
NOR4xp75_ASAP7_75t_L g1370 ( .A(n_1366), .B(n_1232), .C(n_1174), .D(n_1147), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1365), .B(n_1281), .Y(n_1371) );
OAI21xp5_ASAP7_75t_L g1372 ( .A1(n_1369), .A2(n_1368), .B(n_1366), .Y(n_1372) );
OAI21xp5_ASAP7_75t_L g1373 ( .A1(n_1371), .A2(n_1147), .B(n_1194), .Y(n_1373) );
AOI322xp5_ASAP7_75t_L g1374 ( .A1(n_1370), .A2(n_1281), .A3(n_1266), .B1(n_1221), .B2(n_1190), .C1(n_1196), .C2(n_1174), .Y(n_1374) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_1372), .A2(n_1230), .B1(n_1165), .B2(n_1266), .Y(n_1375) );
BUFx2_ASAP7_75t_L g1376 ( .A(n_1373), .Y(n_1376) );
XNOR2xp5_ASAP7_75t_L g1377 ( .A(n_1376), .B(n_1374), .Y(n_1377) );
AOI22xp5_ASAP7_75t_SL g1378 ( .A1(n_1375), .A2(n_1165), .B1(n_1190), .B2(n_1196), .Y(n_1378) );
AOI211xp5_ASAP7_75t_L g1379 ( .A1(n_1377), .A2(n_1195), .B(n_1184), .C(n_1221), .Y(n_1379) );
AOI22x1_ASAP7_75t_L g1380 ( .A1(n_1379), .A2(n_1378), .B1(n_1192), .B2(n_1189), .Y(n_1380) );
AOI222xp33_ASAP7_75t_L g1381 ( .A1(n_1380), .A2(n_1195), .B1(n_1221), .B2(n_1184), .C1(n_1151), .C2(n_1260), .Y(n_1381) );
endmodule