module fake_jpeg_6422_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_20),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_30),
.B1(n_24),
.B2(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_30),
.B1(n_19),
.B2(n_28),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_30),
.B1(n_23),
.B2(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_56),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_35),
.C(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_61),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_33),
.B1(n_25),
.B2(n_17),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_15),
.B1(n_16),
.B2(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_0),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_26),
.C(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_32),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_22),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_68),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_67),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_32),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_53),
.B1(n_48),
.B2(n_57),
.Y(n_86)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_41),
.B1(n_40),
.B2(n_32),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_57),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_27),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_56),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_101),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_40),
.B1(n_41),
.B2(n_59),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_75),
.B1(n_51),
.B2(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_96),
.B1(n_27),
.B2(n_29),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_70),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_98),
.B(n_63),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_73),
.B1(n_74),
.B2(n_71),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_46),
.C(n_59),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_75),
.C(n_77),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_59),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_64),
.B(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_112),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_74),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_113),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_85),
.B1(n_110),
.B2(n_120),
.Y(n_144)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_78),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_121),
.C(n_98),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_104),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_120),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_69),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_99),
.B(n_85),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_77),
.B1(n_51),
.B2(n_29),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_63),
.C(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_127),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_133),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_136),
.C(n_101),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_85),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_144),
.B1(n_67),
.B2(n_63),
.Y(n_163)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_103),
.C(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

AOI322xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_117),
.A3(n_113),
.B1(n_109),
.B2(n_95),
.C1(n_111),
.C2(n_107),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_116),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_85),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_114),
.B1(n_84),
.B2(n_121),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_139),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_87),
.C(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_84),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_91),
.B1(n_100),
.B2(n_83),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_163),
.B1(n_146),
.B2(n_140),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_100),
.B1(n_89),
.B2(n_83),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_141),
.B1(n_127),
.B2(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_134),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_170),
.Y(n_189)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_137),
.C(n_130),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_171),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_177),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_151),
.B1(n_154),
.B2(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_63),
.C(n_89),
.Y(n_190)
);

OAI321xp33_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_136),
.A3(n_138),
.B1(n_135),
.B2(n_67),
.C(n_89),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_155),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_183),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_173),
.Y(n_183)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_158),
.B1(n_153),
.B2(n_149),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_192),
.C(n_31),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_20),
.Y(n_191)
);

NAND4xp25_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_31),
.C(n_29),
.D(n_3),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_82),
.C(n_20),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_176),
.B1(n_170),
.B2(n_167),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_194),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_175),
.B1(n_165),
.B2(n_172),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_172),
.B1(n_82),
.B2(n_31),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_5),
.B(n_7),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_197),
.B(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_192),
.C(n_7),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_202),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_190),
.B(n_196),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_207),
.B(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_194),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_189),
.B(n_180),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_183),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_209),
.C(n_201),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_204),
.B1(n_203),
.B2(n_10),
.Y(n_216)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g220 ( 
.A1(n_211),
.A2(n_8),
.B(n_9),
.C(n_10),
.D(n_11),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_213),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_7),
.C(n_8),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_8),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_13),
.Y(n_223)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_9),
.B(n_10),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_222),
.B(n_223),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_9),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_217),
.B(n_12),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_224),
.Y(n_227)
);


endmodule