module fake_jpeg_13588_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_29),
.B(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_16),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_17),
.B(n_13),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_78),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_60),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_1),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_55),
.B1(n_51),
.B2(n_52),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_90),
.B1(n_62),
.B2(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_87),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_65),
.C(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_66),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_61),
.B1(n_67),
.B2(n_57),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_5),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_102),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_73),
.B1(n_71),
.B2(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_111),
.B1(n_113),
.B2(n_4),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_58),
.B(n_63),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_6),
.B(n_7),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_63),
.B1(n_73),
.B2(n_64),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_112),
.B1(n_8),
.B2(n_9),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_59),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_108),
.Y(n_129)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_60),
.B1(n_54),
.B2(n_41),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_85),
.B1(n_40),
.B2(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_2),
.B(n_3),
.Y(n_117)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_134),
.B(n_14),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_126),
.B1(n_28),
.B2(n_30),
.Y(n_146)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_38),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_14),
.Y(n_139)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_10),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_95),
.C(n_13),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_10),
.B(n_11),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_138),
.C(n_139),
.Y(n_150)
);

NAND2x1_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_12),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_146),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_31),
.C(n_24),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_15),
.B1(n_26),
.B2(n_27),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_114),
.A2(n_116),
.B1(n_134),
.B2(n_119),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_114),
.B1(n_118),
.B2(n_131),
.Y(n_152)
);

OAI322xp33_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_151),
.A3(n_153),
.B1(n_147),
.B2(n_130),
.C1(n_136),
.C2(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_143),
.B1(n_145),
.B2(n_121),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_149),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_155),
.A3(n_152),
.B1(n_138),
.B2(n_140),
.C1(n_142),
.C2(n_154),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_158),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_159),
.C(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_118),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule