module real_jpeg_27113_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_320, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_320;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_0),
.B(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_0),
.B(n_95),
.Y(n_94)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_0),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_0),
.B(n_194),
.Y(n_199)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_4),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_21),
.B1(n_48),
.B2(n_50),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_21),
.B1(n_42),
.B2(n_46),
.Y(n_98)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_6),
.B1(n_20),
.B2(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_5),
.B1(n_20),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_5),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_104),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_5),
.A2(n_42),
.B1(n_46),
.B2(n_104),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_104),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_6),
.A2(n_42),
.B1(n_46),
.B2(n_72),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_274)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_10),
.B(n_48),
.Y(n_184)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_9),
.A2(n_10),
.B(n_42),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_10),
.A2(n_20),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_20),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_42),
.B1(n_46),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_10),
.B(n_33),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_10),
.B(n_58),
.Y(n_188)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_11),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_16),
.C(n_281),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_81),
.B(n_316),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_34),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_16),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_29),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_17),
.A2(n_25),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_18),
.B(n_102),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_22),
.B(n_31),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_22),
.A2(n_25),
.B(n_31),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_24),
.Y(n_125)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_25),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_26),
.B(n_28),
.Y(n_123)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_27),
.A2(n_58),
.B(n_66),
.C(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_27),
.B(n_66),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_27),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_27),
.A2(n_54),
.B(n_59),
.C(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_29),
.B(n_115),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_32),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_35),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_73),
.C(n_75),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_36),
.A2(n_37),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_55),
.C(n_69),
.Y(n_37)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_38),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_38),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_38),
.B(n_55),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_51),
.B(n_52),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_39),
.A2(n_97),
.B(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_40),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_40),
.B(n_98),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_40),
.B(n_164),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_47),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_46),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_42),
.A2(n_44),
.B(n_54),
.C(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_47),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_47),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_47),
.B(n_53),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_50),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_51),
.B(n_54),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_51),
.A2(n_165),
.B(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_54),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_61),
.B(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_57),
.A2(n_64),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_58),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_68),
.Y(n_141)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_62),
.B(n_65),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_110),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_65),
.A2(n_258),
.B(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_69),
.A2(n_70),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_73),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_73),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_73),
.A2(n_75),
.B1(n_242),
.B2(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_75),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_76),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_79),
.B(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_309),
.B(n_315),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_286),
.A3(n_304),
.B1(n_307),
.B2(n_308),
.C(n_320),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_266),
.B(n_285),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_246),
.B(n_265),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_147),
.B(n_228),
.C(n_245),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_133),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_87),
.B(n_133),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_111),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_100),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_89),
.B(n_100),
.C(n_111),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_90),
.B(n_96),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_93),
.B(n_94),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_92),
.B(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_92),
.A2(n_128),
.B(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_92),
.B(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_127),
.B(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_94),
.B(n_193),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_175),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_99),
.B(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_107),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_105),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_106),
.B(n_290),
.C(n_294),
.Y(n_303)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_109),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_121),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_113),
.B(n_118),
.C(n_121),
.Y(n_243)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_126),
.Y(n_138)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_128),
.B(n_146),
.Y(n_192)
);

INVx5_ASAP7_75t_SL g210 ( 
.A(n_128),
.Y(n_210)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_130),
.B(n_192),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_139),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_134),
.A2(n_135),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_141),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_199),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_227),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_220),
.B(n_226),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_177),
.B(n_219),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_166),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_151),
.B(n_166),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.C(n_161),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_152),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_156),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_155),
.A2(n_156),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_155),
.B(n_262),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_155),
.A2(n_156),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_156),
.A2(n_277),
.B(n_282),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_160),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_165),
.B(n_174),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_173),
.C(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_214),
.B(n_218),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_195),
.B(n_213),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_185),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_190),
.C(n_191),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_202),
.B(n_212),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_197),
.B(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_206),
.B(n_211),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_230),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_243),
.B2(n_244),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_237),
.C(n_244),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_248),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_264),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_260),
.B2(n_261),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_261),
.C(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_254),
.C(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_268),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_283),
.B2(n_284),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_276),
.C(n_284),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_273),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_274),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_288),
.C(n_296),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_275),
.B(n_288),
.CI(n_296),
.CON(n_306),
.SN(n_306)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_297),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_290),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_299),
.C(n_303),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_303),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_305),
.B(n_306),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_312),
.Y(n_314)
);


endmodule