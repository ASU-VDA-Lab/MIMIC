module fake_jpeg_23382_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_20),
.B1(n_19),
.B2(n_22),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_23),
.B1(n_15),
.B2(n_22),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_15),
.C(n_22),
.Y(n_64)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_64),
.B(n_35),
.CI(n_37),
.CON(n_107),
.SN(n_107)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_83),
.B1(n_86),
.B2(n_45),
.Y(n_101)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_29),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_24),
.B1(n_28),
.B2(n_36),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_84),
.B1(n_87),
.B2(n_25),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_54),
.Y(n_109)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OA22x2_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_22),
.B1(n_40),
.B2(n_38),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_28),
.B1(n_21),
.B2(n_22),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_26),
.B1(n_17),
.B2(n_18),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_49),
.B1(n_58),
.B2(n_45),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_112),
.B1(n_74),
.B2(n_81),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_101),
.B1(n_82),
.B2(n_79),
.Y(n_113)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_17),
.Y(n_119)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_42),
.B1(n_62),
.B2(n_53),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_131)
);

INVx2_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_105),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_66),
.B(n_64),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_72),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_42),
.B1(n_52),
.B2(n_26),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_130),
.B1(n_108),
.B2(n_98),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_118),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_120),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_79),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_132),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_110),
.B1(n_90),
.B2(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_95),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_81),
.B1(n_25),
.B2(n_60),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_0),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_138),
.B(n_97),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_38),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_137),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_69),
.B1(n_25),
.B2(n_13),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_154),
.B1(n_124),
.B2(n_120),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_107),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_92),
.B1(n_101),
.B2(n_111),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_153),
.B1(n_126),
.B2(n_133),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_93),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_136),
.B(n_129),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_91),
.C(n_94),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_151),
.C(n_160),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_91),
.C(n_94),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_112),
.B1(n_108),
.B2(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_155),
.B(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_157),
.B(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_122),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_40),
.C(n_41),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_37),
.B1(n_60),
.B2(n_72),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_129),
.C(n_138),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_169),
.C(n_184),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_129),
.C(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_171),
.B(n_182),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_146),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_148),
.B(n_152),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_158),
.A2(n_133),
.B1(n_127),
.B2(n_136),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_181),
.B1(n_29),
.B2(n_16),
.Y(n_210)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_179),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_163),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_127),
.B(n_119),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_178),
.B(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_121),
.C(n_41),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_190),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_40),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_37),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_156),
.C(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_204),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g193 ( 
.A1(n_175),
.A2(n_161),
.B(n_158),
.C(n_162),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_193),
.A2(n_195),
.B(n_196),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_200),
.C(n_166),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_161),
.B(n_159),
.C(n_157),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_205),
.B(n_14),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_152),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_121),
.C(n_144),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_190),
.B1(n_173),
.B2(n_179),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_14),
.B(n_13),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_211),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_16),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_214),
.B1(n_115),
.B2(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_16),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_183),
.B(n_29),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_186),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_115),
.B1(n_99),
.B2(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_221),
.B(n_226),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_220),
.C(n_192),
.Y(n_237)
);

NAND2x1_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_176),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_219),
.A2(n_29),
.B(n_2),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_167),
.C(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_199),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_222),
.A2(n_225),
.B1(n_29),
.B2(n_30),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_227),
.B1(n_195),
.B2(n_193),
.Y(n_248)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_172),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_0),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_0),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_0),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_236),
.B(n_1),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_238),
.C(n_251),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_220),
.C(n_192),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_193),
.B1(n_196),
.B2(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_207),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_242),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_207),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_212),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_246),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_194),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_209),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_248),
.A2(n_225),
.B1(n_255),
.B2(n_249),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_195),
.B1(n_201),
.B2(n_205),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_16),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_232),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_222),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_236),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_255),
.A2(n_231),
.B(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

AOI221xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_271),
.B1(n_219),
.B2(n_233),
.C(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_267),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_270),
.B1(n_1),
.B2(n_3),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_221),
.B1(n_234),
.B2(n_217),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_219),
.B1(n_239),
.B2(n_230),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_241),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_242),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_247),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_224),
.Y(n_269)
);

FAx1_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_230),
.CI(n_251),
.CON(n_277),
.SN(n_277)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_252),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_273),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_279),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_238),
.C(n_237),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_277),
.B1(n_272),
.B2(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_260),
.C(n_257),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_250),
.C(n_3),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_1),
.C(n_3),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_286),
.C(n_4),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_259),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_266),
.A2(n_29),
.B1(n_5),
.B2(n_6),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_258),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_4),
.C(n_5),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_292),
.B(n_277),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_297),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_264),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_265),
.C(n_262),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_7),
.C(n_8),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_4),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_4),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_274),
.B1(n_6),
.B2(n_7),
.Y(n_300)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_300),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_5),
.CI(n_7),
.CON(n_303),
.SN(n_303)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_287),
.B1(n_294),
.B2(n_10),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_288),
.C(n_306),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_8),
.B(n_9),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_309),
.B(n_312),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_316),
.B(n_307),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_303),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_315),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_308),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_307),
.B(n_301),
.C(n_11),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_9),
.B(n_11),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_9),
.C(n_30),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_30),
.B(n_295),
.C(n_305),
.Y(n_323)
);


endmodule