module fake_jpeg_584_n_184 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_11),
.B(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_37),
.B(n_40),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_2),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_55),
.Y(n_87)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_32),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_34),
.A2(n_27),
.B1(n_24),
.B2(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_34),
.A2(n_21),
.B1(n_25),
.B2(n_7),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_48),
.B(n_25),
.C(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_81),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_4),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_84),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_39),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_8),
.B(n_52),
.C(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_67),
.Y(n_96)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_88),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_103),
.Y(n_123)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_87),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_62),
.B(n_74),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_64),
.B(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_111),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_60),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_65),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_61),
.B(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_85),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_83),
.A3(n_61),
.B1(n_76),
.B2(n_72),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_126),
.B(n_101),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_56),
.B1(n_64),
.B2(n_79),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_122),
.A2(n_125),
.B1(n_92),
.B2(n_103),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_97),
.A2(n_90),
.B1(n_102),
.B2(n_95),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_56),
.B1(n_69),
.B2(n_83),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_93),
.B1(n_94),
.B2(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_109),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_79),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_103),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_90),
.B1(n_95),
.B2(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_135),
.B1(n_137),
.B2(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_127),
.B(n_111),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_140),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_96),
.B(n_106),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_141),
.A2(n_123),
.B(n_119),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_129),
.C(n_119),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_91),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_126),
.C(n_142),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_152),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_142),
.C(n_131),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_135),
.B1(n_134),
.B2(n_133),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_153),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_94),
.C(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_160),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_148),
.B1(n_130),
.B2(n_117),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_130),
.B(n_120),
.C(n_115),
.D(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_154),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_169),
.B1(n_159),
.B2(n_155),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_161),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_172),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_157),
.C(n_163),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_158),
.C(n_164),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_113),
.Y(n_178)
);

OAI221xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_167),
.B1(n_166),
.B2(n_169),
.C(n_173),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_113),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_105),
.C(n_108),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_181),
.B1(n_79),
.B2(n_100),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_91),
.Y(n_184)
);


endmodule