module fake_jpeg_14204_n_95 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_7),
.B(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_2),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_55),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_68),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_37),
.B1(n_53),
.B2(n_38),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_70),
.B(n_72),
.C(n_3),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_60),
.A2(n_32),
.B(n_33),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_71),
.Y(n_78)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_43),
.A3(n_42),
.B1(n_45),
.B2(n_35),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_55),
.B(n_54),
.C(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_44),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_40),
.B1(n_34),
.B2(n_45),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_17),
.B(n_28),
.C(n_5),
.D(n_11),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_80),
.B(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_4),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_86),
.B(n_85),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_90),
.A2(n_88),
.B1(n_83),
.B2(n_80),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_13),
.B(n_14),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_15),
.A3(n_22),
.B1(n_23),
.B2(n_24),
.C1(n_25),
.C2(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_81),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_94),
.Y(n_95)
);


endmodule