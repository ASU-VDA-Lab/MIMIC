module fake_jpeg_31045_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_4),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_16),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_10),
.B1(n_16),
.B2(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_22),
.B1(n_10),
.B2(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_20),
.C(n_21),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_23),
.C(n_21),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_36),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_22),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_37),
.B1(n_28),
.B2(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_22),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_41),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_18),
.C(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_34),
.B1(n_30),
.B2(n_26),
.Y(n_46)
);

OAI322xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_31),
.A3(n_15),
.B1(n_38),
.B2(n_9),
.C1(n_13),
.C2(n_18),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.C(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_9),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_50),
.B(n_48),
.Y(n_53)
);

FAx1_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_13),
.CI(n_1),
.CON(n_54),
.SN(n_54)
);

AOI31xp67_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_54),
.A3(n_6),
.B(n_0),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_2),
.B(n_5),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B(n_6),
.Y(n_57)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_0),
.A3(n_6),
.B1(n_11),
.B2(n_14),
.C1(n_24),
.C2(n_56),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_11),
.Y(n_59)
);


endmodule