module fake_jpeg_6528_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_41),
.B1(n_27),
.B2(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_51),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_47),
.B1(n_57),
.B2(n_50),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_41),
.B1(n_29),
.B2(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_39),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_77),
.B1(n_20),
.B2(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_29),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_89),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_40),
.B1(n_26),
.B2(n_17),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_81),
.B1(n_20),
.B2(n_28),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_25),
.B(n_32),
.C(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_80),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_52),
.B1(n_51),
.B2(n_41),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_32),
.CI(n_33),
.CON(n_78),
.SN(n_78)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_78),
.B(n_14),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_23),
.B1(n_30),
.B2(n_33),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_23),
.B1(n_25),
.B2(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_90),
.B1(n_56),
.B2(n_62),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_59),
.A2(n_37),
.B1(n_36),
.B2(n_40),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_71),
.A3(n_37),
.B1(n_36),
.B2(n_75),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_91),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_32),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_32),
.B1(n_20),
.B2(n_17),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_60),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_99),
.B1(n_108),
.B2(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_0),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_115),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_36),
.B1(n_37),
.B2(n_56),
.Y(n_99)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_108),
.B1(n_99),
.B2(n_111),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_69),
.B1(n_110),
.B2(n_118),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_64),
.B1(n_84),
.B2(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_112),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_37),
.B1(n_20),
.B2(n_28),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_31),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_89),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_0),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_12),
.B(n_1),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_67),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_69),
.B1(n_76),
.B2(n_67),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_122),
.B1(n_137),
.B2(n_144),
.Y(n_159)
);

NAND2x1p5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_76),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_142),
.B(n_150),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_72),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_149),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_126),
.A2(n_128),
.B1(n_129),
.B2(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_89),
.B1(n_65),
.B2(n_75),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_68),
.B1(n_66),
.B2(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_92),
.C(n_83),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_107),
.C(n_105),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_95),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_98),
.A2(n_62),
.B1(n_91),
.B2(n_31),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_62),
.B1(n_31),
.B2(n_21),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_143),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_31),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_62),
.B1(n_21),
.B2(n_60),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_146),
.Y(n_164)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_95),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_21),
.B(n_1),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_172),
.C(n_173),
.Y(n_192)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_153),
.B(n_158),
.Y(n_193)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_177),
.B(n_181),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_123),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_171),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_165),
.B(n_167),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_94),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g186 ( 
.A(n_170),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_95),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_95),
.C(n_112),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_86),
.C(n_93),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_109),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_175),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_136),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_21),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_86),
.B1(n_88),
.B2(n_74),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_148),
.B1(n_143),
.B2(n_141),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_86),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_184),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_122),
.A2(n_0),
.B(n_1),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_134),
.A2(n_113),
.B(n_106),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_134),
.A2(n_106),
.B(n_2),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_126),
.B(n_149),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_148),
.B1(n_138),
.B2(n_142),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_177),
.B1(n_179),
.B2(n_168),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_137),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_168),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_172),
.C(n_160),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.C(n_208),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_142),
.C(n_135),
.Y(n_200)
);

NOR4xp25_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_10),
.C(n_3),
.D(n_4),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_161),
.C(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_139),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_206),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_164),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_150),
.C(n_144),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_106),
.B1(n_88),
.B2(n_74),
.Y(n_209)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_182),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_213),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_214),
.A2(n_219),
.B1(n_221),
.B2(n_232),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_212),
.A2(n_170),
.B1(n_158),
.B2(n_173),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_220),
.A2(n_236),
.B1(n_197),
.B2(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_177),
.B1(n_181),
.B2(n_159),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_162),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_224),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_228),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_151),
.C(n_157),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_233),
.C(n_192),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_230),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_165),
.B1(n_183),
.B2(n_163),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_152),
.C(n_156),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_0),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_236),
.A2(n_191),
.B(n_195),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_186),
.C(n_202),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_241),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_202),
.CI(n_189),
.CON(n_239),
.SN(n_239)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_239),
.B(n_254),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_232),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_192),
.C(n_189),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_199),
.C(n_190),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_251),
.B1(n_226),
.B2(n_215),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_211),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_199),
.C(n_193),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_252),
.C(n_256),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_210),
.C(n_187),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_2),
.C(n_3),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_220),
.Y(n_265)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_262),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_249),
.C(n_240),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_221),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_269),
.Y(n_274)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_268),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_265),
.A2(n_257),
.B(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_273),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_218),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_214),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_217),
.B1(n_226),
.B2(n_216),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_248),
.B1(n_244),
.B2(n_239),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_264),
.C(n_267),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_6),
.B(n_7),
.Y(n_296)
);

INVx11_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_284),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_260),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_249),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_274),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_239),
.B1(n_241),
.B2(n_5),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_269),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_287),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_258),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_291),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_264),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_283),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_267),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_295),
.C(n_277),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_298),
.B(n_278),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_276),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_278),
.A2(n_7),
.B(n_8),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_290),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_306),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_285),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_275),
.B(n_286),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_305),
.B(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_284),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_289),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_308),
.B(n_310),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_282),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_314),
.B(n_295),
.Y(n_315)
);

OAI21x1_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_299),
.B(n_304),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_292),
.A3(n_294),
.B1(n_313),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_316)
);

OAI321xp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_179),
.C(n_121),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_8),
.Y(n_318)
);


endmodule