module fake_jpeg_18411_n_230 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_33),
.Y(n_44)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_38),
.Y(n_47)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_30),
.B1(n_23),
.B2(n_22),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_49),
.B1(n_26),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_30),
.B1(n_23),
.B2(n_21),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_53),
.B1(n_33),
.B2(n_37),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_22),
.B1(n_21),
.B2(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_29),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_33),
.B1(n_32),
.B2(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_74),
.B1(n_77),
.B2(n_41),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_75),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_29),
.B1(n_17),
.B2(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_20),
.B1(n_24),
.B2(n_27),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_54),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_70),
.C(n_36),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_93),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_43),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_91),
.B(n_36),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_43),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_63),
.B1(n_64),
.B2(n_60),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_41),
.B1(n_66),
.B2(n_78),
.Y(n_115)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_99),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_72),
.B(n_54),
.C(n_75),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_69),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_53),
.Y(n_101)
);

AO21x1_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_90),
.B(n_102),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_59),
.B(n_73),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_103),
.A2(n_122),
.B1(n_80),
.B2(n_91),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_20),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_66),
.B1(n_41),
.B2(n_58),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_76),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_120),
.C(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_87),
.B1(n_91),
.B2(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_69),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_24),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_115),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_24),
.Y(n_125)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_138),
.B1(n_34),
.B2(n_20),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_131),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_104),
.A2(n_122),
.B1(n_103),
.B2(n_107),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_142),
.B1(n_131),
.B2(n_139),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_123),
.B(n_94),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_94),
.B1(n_87),
.B2(n_86),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_97),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_144),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_100),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_113),
.A2(n_86),
.B1(n_100),
.B2(n_93),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_106),
.B1(n_119),
.B2(n_116),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_27),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_109),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_151),
.B(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_125),
.C(n_118),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_161),
.C(n_164),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

AOI22x1_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_124),
.B1(n_108),
.B2(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_147),
.B1(n_140),
.B2(n_130),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_139),
.B1(n_144),
.B2(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_36),
.C(n_34),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_27),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_34),
.C(n_20),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_167),
.B(n_11),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_8),
.Y(n_168)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_136),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_151),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_158),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_143),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_147),
.C(n_137),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_150),
.C(n_157),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_176),
.B1(n_183),
.B2(n_174),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_177),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_192),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_160),
.B1(n_152),
.B2(n_164),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_196),
.B1(n_8),
.B2(n_1),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_170),
.C(n_184),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_173),
.B(n_1),
.Y(n_204)
);

AO221x1_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_165),
.B1(n_152),
.B2(n_2),
.C(n_3),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_178),
.C(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_201),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_202),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_187),
.C(n_185),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_205),
.B(n_11),
.Y(n_209)
);

XOR2x1_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_8),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_206),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_194),
.B1(n_186),
.B2(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_212),
.Y(n_217)
);

OAI321xp33_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_213),
.A3(n_14),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_203),
.C(n_199),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_192),
.C(n_1),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_198),
.B(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_212),
.C(n_210),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_218),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_4),
.B(n_5),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_10),
.C(n_12),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_210),
.C(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_221),
.B(n_10),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_0),
.A3(n_5),
.B1(n_10),
.B2(n_12),
.C1(n_13),
.C2(n_219),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_224),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_227),
.B(n_13),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_0),
.Y(n_230)
);


endmodule