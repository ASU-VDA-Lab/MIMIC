module fake_jpeg_3968_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_23),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_4),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_24),
.B1(n_31),
.B2(n_17),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_54),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_24),
.B1(n_31),
.B2(n_19),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_31),
.B1(n_16),
.B2(n_19),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_23),
.B1(n_27),
.B2(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_27),
.B1(n_21),
.B2(n_30),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_73),
.B1(n_64),
.B2(n_70),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_32),
.A2(n_21),
.B1(n_15),
.B2(n_29),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_66),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_60),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_29),
.B(n_26),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_59),
.A2(n_64),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_70),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

AOI222xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_29),
.B1(n_26),
.B2(n_20),
.C1(n_11),
.C2(n_15),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_20),
.B(n_26),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_20),
.B1(n_6),
.B2(n_7),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_4),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_34),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_34),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_9),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_99),
.B1(n_97),
.B2(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_56),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_71),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_101),
.A2(n_77),
.B(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_68),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_57),
.B1(n_62),
.B2(n_72),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_106),
.B1(n_114),
.B2(n_115),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_72),
.B1(n_75),
.B2(n_77),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_110),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_119),
.B(n_123),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_65),
.C(n_76),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_76),
.Y(n_111)
);

XOR2x2_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_108),
.Y(n_135)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_100),
.B1(n_85),
.B2(n_91),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_87),
.B1(n_91),
.B2(n_80),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_96),
.B1(n_80),
.B2(n_89),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_118),
.B1(n_114),
.B2(n_115),
.Y(n_131)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_104),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_92),
.B(n_86),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_101),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_122),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_88),
.B1(n_83),
.B2(n_95),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_129),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_81),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_112),
.B1(n_117),
.B2(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_136),
.C(n_130),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_103),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_138),
.Y(n_147)
);

AOI211xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_111),
.B(n_106),
.C(n_124),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_143),
.B(n_140),
.C(n_125),
.D(n_129),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_139),
.A2(n_121),
.B(n_110),
.C(n_116),
.D(n_117),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_148),
.B(n_151),
.CI(n_125),
.CON(n_158),
.SN(n_158)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_140),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_112),
.C(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_146),
.B(n_142),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_153),
.B(n_154),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_136),
.B(n_127),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_128),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_157),
.B(n_158),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_160),
.C(n_145),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_151),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_165),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_141),
.B1(n_146),
.B2(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_158),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_147),
.C(n_128),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_158),
.C(n_147),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_169),
.B(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_162),
.B(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_163),
.Y(n_175)
);

OAI211xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_176),
.B(n_164),
.C(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_126),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_173),
.Y(n_180)
);


endmodule