module fake_netlist_6_883_n_331 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_92, n_42, n_8, n_90, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_331);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_92;
input n_42;
input n_8;
input n_90;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_331;

wire n_326;
wire n_256;
wire n_209;
wire n_223;
wire n_278;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_125;
wire n_168;
wire n_297;
wire n_106;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_142;
wire n_143;
wire n_180;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_280;
wire n_287;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_111;
wire n_314;
wire n_183;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_97;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_107;
wire n_103;
wire n_272;
wire n_185;
wire n_293;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_166;
wire n_184;
wire n_216;
wire n_323;
wire n_152;
wire n_321;
wire n_105;
wire n_227;
wire n_132;
wire n_102;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_231;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_317;
wire n_149;
wire n_328;
wire n_195;
wire n_285;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_267;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_170;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVxp67_ASAP7_75t_SL g114 ( 
.A(n_13),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_44),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_41),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_52),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_3),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_15),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVxp33_ASAP7_75t_SL g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_43),
.Y(n_124)
);

INVxp33_ASAP7_75t_SL g125 ( 
.A(n_36),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_79),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_20),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_53),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_48),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_39),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_0),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_100),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_1),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_127),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

BUFx8_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_97),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_6),
.Y(n_164)
);

AO22x2_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_124),
.B1(n_136),
.B2(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_114),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

AO22x2_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_164),
.B1(n_146),
.B2(n_159),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_97),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_111),
.Y(n_177)
);

OAI221xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_130),
.B1(n_122),
.B2(n_133),
.C(n_132),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

OR2x6_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_113),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_125),
.Y(n_185)
);

OR2x2_ASAP7_75t_SL g186 ( 
.A(n_140),
.B(n_137),
.Y(n_186)
);

AO22x2_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_128),
.B1(n_126),
.B2(n_115),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_120),
.B1(n_121),
.B2(n_134),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_117),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

AO22x2_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_7),
.B1(n_8),
.B2(n_125),
.Y(n_196)
);

AO22x2_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_8),
.B1(n_123),
.B2(n_106),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_106),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_116),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_100),
.B1(n_14),
.B2(n_16),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_11),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_168),
.B(n_17),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_175),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_172),
.B1(n_194),
.B2(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_18),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_19),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_21),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_32),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_189),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_34),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_38),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_40),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_42),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_172),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_165),
.B(n_49),
.Y(n_226)
);

AND3x1_ASAP7_75t_SL g227 ( 
.A(n_178),
.B(n_51),
.C(n_55),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_56),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_59),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_60),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_62),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_165),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_235),
.A2(n_73),
.B(n_76),
.C(n_77),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_80),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_82),
.B(n_84),
.C(n_85),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_87),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_88),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_89),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_90),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_204),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_91),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_234),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_201),
.B(n_222),
.C(n_223),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_211),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_199),
.A2(n_200),
.B1(n_225),
.B2(n_228),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_209),
.A2(n_231),
.B1(n_233),
.B2(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_229),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

BUFx4_ASAP7_75t_R g257 ( 
.A(n_229),
.Y(n_257)
);

NOR2x2_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_224),
.B(n_218),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_212),
.A2(n_215),
.B(n_227),
.C(n_213),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_213),
.B(n_244),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_213),
.B1(n_244),
.B2(n_252),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_213),
.B1(n_255),
.B2(n_240),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_261),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_254),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_246),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_236),
.A2(n_247),
.B(n_238),
.C(n_239),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_245),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_256),
.Y(n_276)
);

AOI221xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_260),
.B1(n_257),
.B2(n_259),
.C(n_258),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_258),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_246),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_R g282 ( 
.A(n_242),
.B(n_198),
.Y(n_282)
);

AO21x2_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_262),
.B(n_263),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_265),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_280),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_278),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_291),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_267),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

OR2x6_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_272),
.Y(n_299)
);

NAND2x1_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_272),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_275),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_292),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_292),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_264),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_294),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_298),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_310),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_300),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_283),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_299),
.B1(n_268),
.B2(n_277),
.Y(n_319)
);

NAND2x1_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_312),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_307),
.B(n_308),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_318),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_316),
.Y(n_326)
);

AOI222xp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_323),
.B1(n_322),
.B2(n_316),
.C1(n_314),
.C2(n_325),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_326),
.B1(n_320),
.B2(n_315),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_329),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_328),
.B1(n_282),
.B2(n_268),
.Y(n_331)
);


endmodule