module fake_netlist_1_2354_n_26 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_4), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_3), .B(n_2), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_6), .B(n_7), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_9), .B(n_0), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_14), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
OAI21xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_14), .B(n_17), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_14), .B1(n_16), .B2(n_15), .Y(n_20) );
AOI322xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_15), .A3(n_16), .B1(n_14), .B2(n_8), .C1(n_11), .C2(n_10), .Y(n_21) );
AOI221xp5_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_16), .B1(n_14), .B2(n_13), .C(n_12), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_22), .Y(n_23) );
CKINVDCx6p67_ASAP7_75t_R g24 ( .A(n_21), .Y(n_24) );
NAND3xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_16), .C(n_3), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_24), .B1(n_16), .B2(n_1), .Y(n_26) );
endmodule