module fake_aes_10431_n_591 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_591);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_591;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g71 ( .A(n_54), .Y(n_71) );
CKINVDCx5p33_ASAP7_75t_R g72 ( .A(n_0), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_10), .Y(n_73) );
INVxp67_ASAP7_75t_SL g74 ( .A(n_57), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_63), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_58), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_13), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_49), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_65), .Y(n_79) );
INVx1_ASAP7_75t_SL g80 ( .A(n_36), .Y(n_80) );
NOR2xp67_ASAP7_75t_L g81 ( .A(n_10), .B(n_34), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_62), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_18), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_70), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_44), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_37), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_40), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_7), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_7), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_6), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_43), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_31), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_28), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_15), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_24), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_61), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_20), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_33), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_1), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_8), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_48), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_5), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_26), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_35), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_39), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_45), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_4), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_53), .Y(n_113) );
BUFx6f_ASAP7_75t_SL g114 ( .A(n_75), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_85), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_85), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_83), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_79), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_89), .B(n_0), .Y(n_119) );
BUFx10_ASAP7_75t_L g120 ( .A(n_113), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_97), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_73), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_72), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_103), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_103), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_91), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_103), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_112), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_109), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_73), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_77), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_88), .Y(n_134) );
AOI21x1_ASAP7_75t_L g135 ( .A1(n_75), .A2(n_25), .B(n_68), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_78), .Y(n_137) );
NOR2xp33_ASAP7_75t_R g138 ( .A(n_76), .B(n_69), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_87), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_109), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_93), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_90), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_111), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_100), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_95), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_95), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_78), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
BUFx8_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
NAND2x1p5_ASAP7_75t_L g152 ( .A(n_137), .B(n_111), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_131), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
OAI221xp5_ASAP7_75t_L g155 ( .A1(n_137), .A2(n_98), .B1(n_110), .B2(n_101), .C(n_106), .Y(n_155) );
AO22x2_ASAP7_75t_L g156 ( .A1(n_119), .A2(n_98), .B1(n_96), .B2(n_107), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_115), .B(n_71), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_115), .B(n_116), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_116), .B(n_71), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_120), .B(n_104), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
AO22x2_ASAP7_75t_L g165 ( .A1(n_119), .A2(n_74), .B1(n_96), .B2(n_107), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_149), .B(n_94), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_122), .A2(n_110), .B1(n_101), .B2(n_106), .Y(n_168) );
OR2x2_ASAP7_75t_SL g169 ( .A(n_134), .B(n_108), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_143), .B(n_108), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_143), .B(n_120), .Y(n_173) );
OR2x2_ASAP7_75t_SL g174 ( .A(n_142), .B(n_105), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_120), .B(n_105), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_149), .A2(n_74), .B1(n_104), .B2(n_99), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_125), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_127), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_139), .B(n_86), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_125), .A2(n_86), .B1(n_99), .B2(n_94), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_124), .B(n_80), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_126), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_139), .B(n_92), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_141), .B(n_92), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_128), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_114), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_114), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_124), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_129), .B(n_80), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_195), .B(n_129), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_195), .B(n_118), .Y(n_198) );
O2A1O1Ixp5_ASAP7_75t_L g199 ( .A1(n_194), .A2(n_135), .B(n_102), .C(n_84), .Y(n_199) );
BUFx4f_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
OAI21xp33_ASAP7_75t_SL g201 ( .A1(n_173), .A2(n_84), .B(n_81), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_170), .A2(n_82), .B(n_81), .C(n_145), .Y(n_203) );
NOR2x1_ASAP7_75t_L g204 ( .A(n_159), .B(n_130), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_152), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_172), .A2(n_145), .B(n_141), .C(n_140), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_157), .B(n_118), .Y(n_208) );
NOR2xp33_ASAP7_75t_R g209 ( .A(n_151), .B(n_121), .Y(n_209) );
AO22x1_ASAP7_75t_L g210 ( .A1(n_151), .A2(n_117), .B1(n_138), .B2(n_4), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g211 ( .A1(n_194), .A2(n_67), .B(n_66), .C(n_64), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_153), .A2(n_60), .B(n_59), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_167), .B(n_56), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_158), .A2(n_55), .B(n_52), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_SL g215 ( .A1(n_162), .A2(n_51), .B(n_50), .C(n_46), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
INVx3_ASAP7_75t_SL g217 ( .A(n_184), .Y(n_217) );
NOR3xp33_ASAP7_75t_SL g218 ( .A(n_184), .B(n_1), .C(n_3), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_160), .A2(n_42), .B(n_41), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_176), .A2(n_5), .B(n_6), .C(n_8), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_183), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_187), .B(n_9), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_179), .A2(n_9), .B(n_11), .C(n_12), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_187), .B(n_11), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_167), .B(n_38), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_171), .A2(n_32), .B(n_30), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_165), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_165), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_188), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_155), .A2(n_16), .B(n_17), .C(n_18), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_165), .A2(n_17), .B1(n_19), .B2(n_20), .Y(n_232) );
AOI221xp5_ASAP7_75t_L g233 ( .A1(n_156), .A2(n_19), .B1(n_21), .B2(n_22), .C(n_23), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_165), .A2(n_21), .B1(n_23), .B2(n_27), .Y(n_234) );
BUFx4f_ASAP7_75t_L g235 ( .A(n_196), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_180), .A2(n_29), .B(n_182), .C(n_185), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_177), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_177), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_156), .A2(n_161), .B1(n_181), .B2(n_168), .Y(n_239) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_189), .A2(n_190), .B(n_175), .Y(n_240) );
NOR2xp33_ASAP7_75t_R g241 ( .A(n_151), .B(n_193), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_191), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_178), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_186), .B(n_181), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_196), .B(n_192), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
OAI22xp33_ASAP7_75t_SL g248 ( .A1(n_234), .A2(n_181), .B1(n_186), .B2(n_156), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_209), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_202), .B(n_156), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_205), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_221), .Y(n_252) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_199), .A2(n_154), .B(n_150), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_226), .Y(n_254) );
AO31x2_ASAP7_75t_L g255 ( .A1(n_245), .A2(n_150), .A3(n_166), .B(n_163), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_213), .A2(n_154), .B(n_163), .Y(n_256) );
INVx4_ASAP7_75t_SL g257 ( .A(n_205), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_213), .A2(n_164), .B(n_166), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_235), .B(n_181), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_203), .A2(n_164), .B(n_186), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_242), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_198), .B(n_174), .Y(n_262) );
INVxp67_ASAP7_75t_L g263 ( .A(n_205), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_245), .A2(n_186), .B(n_169), .Y(n_265) );
NAND2x1p5_ASAP7_75t_L g266 ( .A(n_216), .B(n_169), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_243), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_227), .A2(n_174), .B(n_219), .Y(n_268) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_219), .B(n_214), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_235), .B(n_197), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_200), .A2(n_240), .B(n_244), .Y(n_271) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_214), .A2(n_236), .B(n_212), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_225), .A2(n_222), .B(n_238), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_240), .B(n_216), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_216), .B(n_224), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_217), .Y(n_276) );
AO21x2_ASAP7_75t_L g277 ( .A1(n_215), .A2(n_211), .B(n_223), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_246), .B(n_200), .Y(n_278) );
OR2x6_ASAP7_75t_L g279 ( .A(n_222), .B(n_234), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_226), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_226), .B(n_230), .Y(n_281) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_220), .A2(n_229), .B(n_232), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_238), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_239), .A2(n_228), .B(n_232), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_228), .A2(n_231), .B(n_233), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_230), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_279), .A2(n_233), .B1(n_204), .B2(n_208), .Y(n_287) );
OAI222xp33_ASAP7_75t_L g288 ( .A1(n_279), .A2(n_218), .B1(n_210), .B2(n_201), .C1(n_207), .C2(n_241), .Y(n_288) );
NOR2xp33_ASAP7_75t_R g289 ( .A(n_276), .B(n_230), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_257), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_250), .B(n_261), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_257), .B(n_261), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_250), .B(n_270), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
XNOR2xp5_ASAP7_75t_L g295 ( .A(n_250), .B(n_279), .Y(n_295) );
BUFx10_ASAP7_75t_L g296 ( .A(n_250), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_270), .B(n_279), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_251), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g299 ( .A(n_249), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_262), .B(n_278), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_279), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_251), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_257), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_262), .B(n_278), .Y(n_305) );
BUFx4f_ASAP7_75t_SL g306 ( .A(n_251), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_251), .B(n_275), .Y(n_307) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_279), .A2(n_259), .B1(n_274), .B2(n_266), .Y(n_308) );
OAI21xp5_ASAP7_75t_SL g309 ( .A1(n_259), .A2(n_266), .B(n_271), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_257), .B(n_263), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_257), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_300), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_291), .Y(n_314) );
AOI21xp33_ASAP7_75t_L g315 ( .A1(n_287), .A2(n_248), .B(n_265), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_303), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_303), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_303), .Y(n_318) );
A2O1A1Ixp33_ASAP7_75t_L g319 ( .A1(n_287), .A2(n_268), .B(n_285), .C(n_284), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_303), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_301), .A2(n_248), .B1(n_282), .B2(n_284), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_303), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_301), .B(n_284), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_295), .B(n_274), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_291), .B(n_282), .Y(n_325) );
AOI211xp5_ASAP7_75t_L g326 ( .A1(n_288), .A2(n_285), .B(n_268), .C(n_260), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_307), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_295), .A2(n_282), .B1(n_265), .B2(n_285), .Y(n_328) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_300), .B(n_260), .C(n_271), .D(n_275), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_305), .B(n_265), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_307), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_293), .B(n_282), .Y(n_332) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_303), .B(n_286), .Y(n_333) );
OAI21xp33_ASAP7_75t_L g334 ( .A1(n_305), .A2(n_268), .B(n_266), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_294), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_289), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_325), .B(n_297), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_318), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_325), .B(n_308), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_332), .B(n_297), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_332), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_319), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_321), .B(n_309), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_321), .B(n_309), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_324), .B(n_308), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_316), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_336), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_314), .B(n_265), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_316), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_323), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_328), .B(n_293), .Y(n_352) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_329), .B(n_306), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_314), .B(n_292), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_330), .B(n_310), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_324), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_326), .B(n_292), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_327), .B(n_292), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_315), .B(n_331), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_313), .B(n_310), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_334), .B(n_310), .Y(n_361) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_327), .B(n_312), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_318), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_335), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_318), .B(n_312), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_318), .Y(n_366) );
INVx4_ASAP7_75t_L g367 ( .A(n_318), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_363), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_364), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_364), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_364), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_337), .B(n_331), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_337), .B(n_335), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_367), .Y(n_375) );
AND2x4_ASAP7_75t_SL g376 ( .A(n_358), .B(n_296), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_337), .B(n_340), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_346), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_337), .B(n_322), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_350), .Y(n_380) );
OAI31xp33_ASAP7_75t_L g381 ( .A1(n_353), .A2(n_288), .A3(n_292), .B(n_275), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
AO21x2_ASAP7_75t_L g383 ( .A1(n_342), .A2(n_317), .B(n_322), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_342), .B(n_269), .C(n_333), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_351), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_347), .B(n_299), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_351), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_357), .B(n_320), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_341), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_341), .B(n_255), .Y(n_392) );
CKINVDCx11_ASAP7_75t_R g393 ( .A(n_365), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_341), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_346), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_348), .B(n_255), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_347), .B(n_299), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_348), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_363), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_359), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_346), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_349), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_355), .B(n_255), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_340), .B(n_320), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_359), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_361), .A2(n_317), .B(n_333), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_340), .B(n_255), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_359), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_349), .Y(n_411) );
NAND2xp33_ASAP7_75t_L g412 ( .A(n_375), .B(n_362), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_393), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_370), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_387), .B(n_356), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_371), .Y(n_417) );
AOI211x1_ASAP7_75t_L g418 ( .A1(n_377), .A2(n_357), .B(n_343), .C(n_344), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_409), .A2(n_353), .B1(n_356), .B2(n_352), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_401), .Y(n_420) );
AOI211xp5_ASAP7_75t_L g421 ( .A1(n_381), .A2(n_345), .B(n_357), .C(n_343), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_391), .A2(n_342), .B1(n_344), .B2(n_343), .C(n_352), .Y(n_423) );
NOR2x1_ASAP7_75t_SL g424 ( .A(n_375), .B(n_345), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_398), .B(n_344), .Y(n_425) );
OAI32xp33_ASAP7_75t_SL g426 ( .A1(n_385), .A2(n_360), .A3(n_345), .B1(n_339), .B2(n_352), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_398), .B(n_339), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_391), .B(n_355), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_394), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_377), .B(n_358), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_397), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
INVx3_ASAP7_75t_L g433 ( .A(n_375), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_373), .B(n_354), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_409), .A2(n_354), .B1(n_358), .B2(n_362), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_376), .A2(n_354), .B1(n_362), .B2(n_310), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_373), .B(n_360), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_372), .Y(n_438) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_400), .A2(n_361), .B(n_360), .Y(n_439) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_381), .A2(n_273), .B(n_272), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_372), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_380), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_374), .B(n_349), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_380), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_400), .A2(n_349), .B1(n_283), .B2(n_247), .C(n_252), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_401), .Y(n_446) );
OAI22xp33_ASAP7_75t_L g447 ( .A1(n_369), .A2(n_290), .B1(n_304), .B2(n_367), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_369), .A2(n_367), .B1(n_365), .B2(n_290), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_376), .A2(n_367), .B1(n_365), .B2(n_304), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g450 ( .A(n_385), .B(n_269), .C(n_367), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_382), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_392), .A2(n_307), .B(n_263), .C(n_247), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_374), .B(n_367), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_382), .B(n_365), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_379), .B(n_366), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_405), .B(n_365), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_379), .B(n_366), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_384), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_376), .A2(n_296), .B1(n_311), .B2(n_273), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_390), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_384), .B(n_338), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_386), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_413), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_457), .B(n_406), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_430), .B(n_410), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_410), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_415), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_425), .B(n_406), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_423), .B(n_407), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_414), .B(n_386), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_420), .Y(n_472) );
XOR2xp5_ASAP7_75t_L g473 ( .A(n_414), .B(n_405), .Y(n_473) );
OR2x6_ASAP7_75t_L g474 ( .A(n_448), .B(n_390), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_417), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_422), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_427), .B(n_407), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_429), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_431), .B(n_388), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_453), .A2(n_392), .B(n_273), .Y(n_480) );
INVx3_ASAP7_75t_SL g481 ( .A(n_433), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_432), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_427), .B(n_388), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_438), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_412), .B(n_411), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_463), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_454), .B(n_389), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_443), .B(n_389), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_416), .B(n_390), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_434), .B(n_404), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_456), .B(n_402), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_441), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_444), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_452), .B(n_389), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_459), .B(n_389), .Y(n_496) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_433), .B(n_411), .Y(n_497) );
INVx2_ASAP7_75t_SL g498 ( .A(n_446), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_418), .B(n_404), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_428), .B(n_396), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_428), .B(n_396), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_437), .B(n_378), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_461), .B(n_368), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_455), .B(n_368), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_424), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_462), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_421), .B(n_395), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_451), .B(n_395), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_435), .B(n_383), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_449), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_510), .A2(n_449), .B(n_440), .C(n_448), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_505), .A2(n_419), .B(n_450), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_473), .B(n_439), .Y(n_513) );
INVxp33_ASAP7_75t_L g514 ( .A(n_473), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_471), .B(n_440), .C(n_436), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g516 ( .A1(n_479), .A2(n_426), .B1(n_447), .B2(n_445), .C(n_458), .Y(n_516) );
AOI221xp5_ASAP7_75t_SL g517 ( .A1(n_499), .A2(n_399), .B1(n_403), .B2(n_395), .C(n_378), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_485), .A2(n_399), .B(n_403), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_474), .A2(n_460), .B1(n_383), .B2(n_403), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_470), .A2(n_378), .B1(n_296), .B2(n_311), .C1(n_408), .C2(n_306), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_467), .B(n_383), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_490), .A2(n_383), .B1(n_311), .B2(n_283), .C(n_252), .Y(n_522) );
OAI211xp5_ASAP7_75t_SL g523 ( .A1(n_507), .A2(n_338), .B(n_264), .C(n_267), .Y(n_523) );
OAI21xp33_ASAP7_75t_SL g524 ( .A1(n_474), .A2(n_408), .B(n_338), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_509), .A2(n_311), .B1(n_264), .B2(n_267), .C(n_338), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g526 ( .A1(n_509), .A2(n_408), .B(n_363), .Y(n_526) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_497), .A2(n_272), .B(n_338), .Y(n_527) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_500), .A2(n_296), .B1(n_363), .B2(n_338), .C1(n_272), .C2(n_298), .Y(n_528) );
AOI222xp33_ASAP7_75t_L g529 ( .A1(n_501), .A2(n_302), .B1(n_298), .B2(n_294), .C1(n_286), .C2(n_256), .Y(n_529) );
OAI211xp5_ASAP7_75t_L g530 ( .A1(n_489), .A2(n_269), .B(n_281), .C(n_298), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_468), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_506), .A2(n_277), .B1(n_294), .B2(n_302), .C(n_280), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_474), .A2(n_269), .B1(n_277), .B2(n_302), .Y(n_533) );
NOR2xp33_ASAP7_75t_R g534 ( .A(n_481), .B(n_280), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_474), .A2(n_269), .B1(n_277), .B2(n_256), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_477), .A2(n_277), .B1(n_254), .B2(n_280), .C(n_255), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_481), .B(n_256), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_491), .A2(n_503), .B1(n_504), .B2(n_469), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_467), .A2(n_254), .B1(n_255), .B2(n_253), .C(n_258), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_487), .A2(n_258), .B1(n_254), .B2(n_253), .Y(n_540) );
AOI211x1_ASAP7_75t_SL g541 ( .A1(n_480), .A2(n_253), .B(n_258), .C(n_483), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_498), .B(n_472), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_495), .A2(n_496), .B1(n_466), .B2(n_465), .Y(n_543) );
OAI21xp33_ASAP7_75t_L g544 ( .A1(n_519), .A2(n_466), .B(n_465), .Y(n_544) );
AO21x1_ASAP7_75t_L g545 ( .A1(n_514), .A2(n_464), .B(n_493), .Y(n_545) );
AOI21xp33_ASAP7_75t_L g546 ( .A1(n_511), .A2(n_486), .B(n_475), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_513), .A2(n_495), .B1(n_496), .B2(n_487), .Y(n_547) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_542), .B(n_491), .Y(n_548) );
NAND3x1_ASAP7_75t_SL g549 ( .A(n_512), .B(n_488), .C(n_498), .Y(n_549) );
OAI211xp5_ASAP7_75t_L g550 ( .A1(n_516), .A2(n_482), .B(n_492), .C(n_502), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_521), .B(n_484), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_543), .B(n_484), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_538), .B(n_488), .Y(n_553) );
NAND4xp25_ASAP7_75t_SL g554 ( .A(n_524), .B(n_468), .C(n_476), .D(n_478), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_531), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_523), .B(n_476), .C(n_478), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_526), .A2(n_494), .B1(n_508), .B2(n_515), .C(n_517), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_523), .B(n_494), .C(n_530), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_537), .A2(n_520), .B(n_528), .C(n_527), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_518), .B(n_533), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_525), .B(n_522), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g562 ( .A(n_536), .B(n_532), .C(n_539), .Y(n_562) );
NAND3x1_ASAP7_75t_SL g563 ( .A(n_534), .B(n_541), .C(n_529), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_548), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_551), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_545), .A2(n_540), .B(n_535), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_555), .Y(n_567) );
NOR2xp33_ASAP7_75t_R g568 ( .A(n_554), .B(n_561), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_553), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_560), .Y(n_570) );
CKINVDCx16_ASAP7_75t_R g571 ( .A(n_549), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_552), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_546), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_547), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_546), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_565), .Y(n_576) );
AND3x2_ASAP7_75t_L g577 ( .A(n_564), .B(n_558), .C(n_556), .Y(n_577) );
NOR3xp33_ASAP7_75t_L g578 ( .A(n_570), .B(n_550), .C(n_563), .Y(n_578) );
OR4x1_ASAP7_75t_L g579 ( .A(n_571), .B(n_559), .C(n_544), .D(n_557), .Y(n_579) );
OA21x2_ASAP7_75t_L g580 ( .A1(n_570), .A2(n_562), .B(n_564), .Y(n_580) );
CKINVDCx16_ASAP7_75t_R g581 ( .A(n_571), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_567), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_581), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_582), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_578), .A2(n_575), .B(n_573), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_580), .A2(n_574), .B1(n_569), .B2(n_572), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_586), .A2(n_577), .B1(n_575), .B2(n_573), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_583), .A2(n_580), .B1(n_576), .B2(n_579), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_588), .A2(n_585), .B1(n_580), .B2(n_584), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_587), .A2(n_576), .B1(n_579), .B2(n_566), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_590), .A2(n_565), .B1(n_568), .B2(n_589), .Y(n_591) );
endmodule