module fake_jpeg_26189_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

MAJIxp5_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_0),
.C(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_0),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_13),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_2),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2x1_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_3),
.B1(n_10),
.B2(n_7),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_8),
.A2(n_3),
.B(n_11),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_11),
.Y(n_23)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_8),
.B(n_11),
.C(n_12),
.D(n_14),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_25),
.B1(n_18),
.B2(n_15),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_26),
.C(n_24),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_13),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_22),
.B(n_25),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.C(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.C(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_30),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_29),
.B2(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_25),
.Y(n_39)
);


endmodule