module real_aes_8494_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_713;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_1), .A2(n_144), .B(n_149), .C(n_186), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_2), .A2(n_139), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g455 ( .A(n_3), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_4), .B(n_163), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_5), .A2(n_15), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_5), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_6), .A2(n_139), .B(n_473), .Y(n_472) );
AND2x6_ASAP7_75t_L g144 ( .A(n_7), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g173 ( .A(n_8), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_9), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_9), .B(n_43), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_10), .A2(n_251), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_11), .B(n_154), .Y(n_190) );
INVx1_ASAP7_75t_L g477 ( .A(n_12), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_13), .B(n_153), .Y(n_525) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_15), .Y(n_716) );
INVx1_ASAP7_75t_L g537 ( .A(n_16), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_17), .A2(n_174), .B(n_199), .C(n_201), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_18), .B(n_163), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_19), .B(n_466), .Y(n_516) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_20), .A2(n_443), .B1(n_715), .B2(n_718), .C1(n_721), .C2(n_725), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_21), .B(n_139), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_22), .B(n_259), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_23), .A2(n_153), .B(n_155), .C(n_159), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_24), .B(n_163), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_25), .B(n_154), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_26), .A2(n_157), .B(n_201), .C(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_27), .B(n_154), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_28), .Y(n_219) );
INVx1_ASAP7_75t_L g233 ( .A(n_29), .Y(n_233) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_30), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_31), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_32), .B(n_154), .Y(n_456) );
INVx1_ASAP7_75t_L g256 ( .A(n_33), .Y(n_256) );
INVx1_ASAP7_75t_L g490 ( .A(n_34), .Y(n_490) );
INVx2_ASAP7_75t_L g142 ( .A(n_35), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_36), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_37), .A2(n_153), .B(n_212), .C(n_214), .Y(n_211) );
INVxp67_ASAP7_75t_L g257 ( .A(n_38), .Y(n_257) );
CKINVDCx14_ASAP7_75t_R g210 ( .A(n_39), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_40), .A2(n_149), .B(n_232), .C(n_238), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_41), .A2(n_144), .B(n_149), .C(n_505), .Y(n_504) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_42), .A2(n_90), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_42), .Y(n_123) );
INVx1_ASAP7_75t_L g113 ( .A(n_43), .Y(n_113) );
INVx1_ASAP7_75t_L g489 ( .A(n_44), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_45), .A2(n_171), .B(n_172), .C(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_46), .B(n_154), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_47), .B(n_440), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_48), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_49), .Y(n_253) );
INVx1_ASAP7_75t_L g147 ( .A(n_50), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_51), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_52), .B(n_139), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_53), .A2(n_149), .B1(n_159), .B2(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_54), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_55), .Y(n_452) );
CKINVDCx14_ASAP7_75t_R g169 ( .A(n_56), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_57), .A2(n_171), .B(n_214), .C(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_58), .Y(n_518) );
INVx1_ASAP7_75t_L g474 ( .A(n_59), .Y(n_474) );
INVx1_ASAP7_75t_L g145 ( .A(n_60), .Y(n_145) );
INVx1_ASAP7_75t_L g136 ( .A(n_61), .Y(n_136) );
INVx1_ASAP7_75t_SL g213 ( .A(n_62), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_63), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_64), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g222 ( .A(n_65), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_SL g465 ( .A1(n_66), .A2(n_214), .B(n_466), .C(n_467), .Y(n_465) );
INVxp67_ASAP7_75t_L g468 ( .A(n_67), .Y(n_468) );
INVx1_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_69), .A2(n_139), .B(n_168), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_70), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_71), .A2(n_139), .B(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_72), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_73), .A2(n_102), .B1(n_114), .B2(n_727), .Y(n_101) );
INVx1_ASAP7_75t_L g512 ( .A(n_74), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_75), .A2(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g197 ( .A(n_76), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_77), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_78), .A2(n_144), .B(n_149), .C(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_79), .A2(n_139), .B(n_146), .Y(n_138) );
INVx1_ASAP7_75t_L g200 ( .A(n_80), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_81), .B(n_234), .Y(n_506) );
INVx2_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g187 ( .A(n_83), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_84), .B(n_466), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_85), .A2(n_144), .B(n_149), .C(n_454), .Y(n_453) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_86), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g435 ( .A(n_86), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g713 ( .A(n_86), .Y(n_713) );
OR2x2_ASAP7_75t_L g714 ( .A(n_86), .B(n_437), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_87), .A2(n_149), .B(n_221), .C(n_224), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_88), .B(n_166), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_89), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_90), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_91), .A2(n_144), .B(n_149), .C(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_92), .Y(n_529) );
INVx1_ASAP7_75t_L g464 ( .A(n_93), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_94), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_95), .B(n_234), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_96), .B(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_97), .B(n_132), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g156 ( .A(n_99), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_100), .A2(n_139), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g727 ( .A(n_102), .Y(n_727) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_111), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g437 ( .A(n_107), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_441), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g726 ( .A(n_117), .Y(n_726) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_432), .B(n_439), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_124), .B1(n_430), .B2(n_431), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_121), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_124), .A2(n_712), .B1(n_722), .B2(n_723), .Y(n_721) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g431 ( .A(n_125), .Y(n_431) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_356), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_298), .C(n_328), .D(n_338), .Y(n_126) );
OAI211xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_203), .B(n_261), .C(n_288), .Y(n_127) );
OAI222xp33_ASAP7_75t_L g383 ( .A1(n_128), .A2(n_303), .B1(n_384), .B2(n_385), .C1(n_386), .C2(n_387), .Y(n_383) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_178), .Y(n_128) );
AOI33xp33_ASAP7_75t_L g309 ( .A1(n_129), .A2(n_296), .A3(n_297), .B1(n_310), .B2(n_315), .B3(n_317), .Y(n_309) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_129), .A2(n_367), .B(n_369), .C(n_371), .Y(n_366) );
OR2x2_ASAP7_75t_L g382 ( .A(n_129), .B(n_368), .Y(n_382) );
INVx1_ASAP7_75t_L g415 ( .A(n_129), .Y(n_415) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
INVx2_ASAP7_75t_L g292 ( .A(n_130), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_130), .B(n_194), .Y(n_308) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_130), .Y(n_343) );
AND2x2_ASAP7_75t_L g372 ( .A(n_130), .B(n_165), .Y(n_372) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_162), .Y(n_130) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_131), .A2(n_195), .B(n_202), .Y(n_194) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_131), .A2(n_208), .B(n_216), .Y(n_207) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_132), .A2(n_462), .B(n_469), .Y(n_461) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g249 ( .A(n_133), .Y(n_249) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_134), .B(n_135), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx2_ASAP7_75t_L g251 ( .A(n_139), .Y(n_251) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_140), .B(n_144), .Y(n_184) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g237 ( .A(n_141), .Y(n_237) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g150 ( .A(n_142), .Y(n_150) );
INVx1_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
INVx1_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
INVx3_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
INVx1_ASAP7_75t_L g466 ( .A(n_143), .Y(n_466) );
INVx4_ASAP7_75t_SL g161 ( .A(n_144), .Y(n_161) );
BUFx3_ASAP7_75t_L g238 ( .A(n_144), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_148), .B(n_152), .C(n_161), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_148), .A2(n_161), .B(n_169), .C(n_170), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g196 ( .A1(n_148), .A2(n_161), .B(n_197), .C(n_198), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_148), .A2(n_161), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_148), .A2(n_161), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_148), .A2(n_161), .B(n_464), .C(n_465), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_148), .A2(n_161), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_148), .A2(n_161), .B(n_534), .C(n_535), .Y(n_533) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
BUFx3_ASAP7_75t_L g176 ( .A(n_150), .Y(n_176) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_153), .B(n_213), .Y(n_212) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_157), .B(n_200), .Y(n_199) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_157), .A2(n_234), .B1(n_256), .B2(n_257), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_157), .B(n_537), .Y(n_536) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g488 ( .A1(n_158), .A2(n_189), .B1(n_489), .B2(n_490), .Y(n_488) );
INVx2_ASAP7_75t_L g457 ( .A(n_159), .Y(n_457) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_161), .A2(n_184), .B1(n_487), .B2(n_491), .Y(n_486) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_163), .A2(n_472), .B(n_478), .Y(n_471) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_164), .B(n_193), .Y(n_192) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_164), .A2(n_218), .B(n_225), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_164), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_SL g508 ( .A(n_164), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g272 ( .A(n_165), .Y(n_272) );
BUFx3_ASAP7_75t_L g280 ( .A(n_165), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_165), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g291 ( .A(n_165), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_165), .B(n_179), .Y(n_320) );
AND2x2_ASAP7_75t_L g389 ( .A(n_165), .B(n_323), .Y(n_389) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_177), .Y(n_165) );
INVx1_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx2_ASAP7_75t_L g227 ( .A(n_166), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_166), .A2(n_184), .B(n_230), .C(n_231), .Y(n_229) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_166), .A2(n_532), .B(n_538), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx5_ASAP7_75t_L g234 ( .A(n_174), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_174), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_174), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
INVx2_ASAP7_75t_SL g283 ( .A(n_178), .Y(n_283) );
OR2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_194), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_179), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g325 ( .A(n_179), .Y(n_325) );
AND2x2_ASAP7_75t_L g336 ( .A(n_179), .B(n_292), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_179), .B(n_321), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_179), .B(n_323), .Y(n_368) );
AND2x2_ASAP7_75t_L g427 ( .A(n_179), .B(n_372), .Y(n_427) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g297 ( .A(n_180), .B(n_194), .Y(n_297) );
AND2x2_ASAP7_75t_L g307 ( .A(n_180), .B(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g329 ( .A(n_180), .Y(n_329) );
AND3x2_ASAP7_75t_L g388 ( .A(n_180), .B(n_389), .C(n_390), .Y(n_388) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_192), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_181), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_181), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_181), .B(n_529), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_184), .A2(n_219), .B(n_220), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_184), .A2(n_452), .B(n_453), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_184), .A2(n_512), .B(n_513), .Y(n_511) );
O2A1O1Ixp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_190), .C(n_191), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_188), .A2(n_191), .B(n_222), .C(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_191), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_191), .A2(n_515), .B(n_516), .Y(n_514) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_194), .Y(n_279) );
INVx1_ASAP7_75t_SL g323 ( .A(n_194), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_194), .B(n_272), .C(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_241), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_204), .A2(n_307), .B(n_359), .C(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_206), .B(n_228), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_206), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_SL g375 ( .A(n_206), .Y(n_375) );
AND2x2_ASAP7_75t_L g396 ( .A(n_206), .B(n_243), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_206), .B(n_305), .Y(n_424) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
AND2x2_ASAP7_75t_L g269 ( .A(n_207), .B(n_260), .Y(n_269) );
INVx2_ASAP7_75t_L g276 ( .A(n_207), .Y(n_276) );
AND2x2_ASAP7_75t_L g296 ( .A(n_207), .B(n_243), .Y(n_296) );
AND2x2_ASAP7_75t_L g346 ( .A(n_207), .B(n_228), .Y(n_346) );
INVx1_ASAP7_75t_L g350 ( .A(n_207), .Y(n_350) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_215), .Y(n_526) );
INVx2_ASAP7_75t_SL g260 ( .A(n_217), .Y(n_260) );
BUFx2_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
AND2x2_ASAP7_75t_L g413 ( .A(n_217), .B(n_228), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g259 ( .A(n_227), .Y(n_259) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_227), .A2(n_521), .B(n_528), .Y(n_520) );
INVx3_ASAP7_75t_SL g243 ( .A(n_228), .Y(n_243) );
AND2x2_ASAP7_75t_L g268 ( .A(n_228), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g275 ( .A(n_228), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g305 ( .A(n_228), .B(n_265), .Y(n_305) );
OR2x2_ASAP7_75t_L g314 ( .A(n_228), .B(n_260), .Y(n_314) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_228), .Y(n_332) );
AND2x2_ASAP7_75t_L g337 ( .A(n_228), .B(n_290), .Y(n_337) );
AND2x2_ASAP7_75t_L g365 ( .A(n_228), .B(n_245), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_228), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g403 ( .A(n_228), .B(n_244), .Y(n_403) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_239), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .C(n_236), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_234), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_237), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g327 ( .A(n_243), .B(n_276), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_243), .B(n_269), .Y(n_355) );
AND2x2_ASAP7_75t_L g373 ( .A(n_243), .B(n_290), .Y(n_373) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_260), .Y(n_244) );
AND2x2_ASAP7_75t_L g274 ( .A(n_245), .B(n_260), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_245), .B(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g312 ( .A(n_245), .Y(n_312) );
OR2x2_ASAP7_75t_L g360 ( .A(n_245), .B(n_280), .Y(n_360) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_250), .B(n_258), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_247), .A2(n_266), .B(n_267), .Y(n_265) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_247), .A2(n_511), .B(n_517), .Y(n_510) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AOI21xp5_ASAP7_75t_SL g502 ( .A1(n_248), .A2(n_503), .B(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_249), .A2(n_451), .B(n_458), .Y(n_450) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_249), .A2(n_486), .B(n_492), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_249), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g266 ( .A(n_250), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_258), .Y(n_267) );
AND2x2_ASAP7_75t_L g295 ( .A(n_260), .B(n_265), .Y(n_295) );
INVx1_ASAP7_75t_L g303 ( .A(n_260), .Y(n_303) );
AND2x2_ASAP7_75t_L g398 ( .A(n_260), .B(n_276), .Y(n_398) );
AOI222xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_270), .B1(n_273), .B2(n_277), .C1(n_281), .C2(n_284), .Y(n_261) );
INVx1_ASAP7_75t_L g393 ( .A(n_262), .Y(n_393) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_268), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_263), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g300 ( .A(n_263), .B(n_269), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_263), .B(n_291), .Y(n_316) );
OAI222xp33_ASAP7_75t_L g338 ( .A1(n_263), .A2(n_339), .B1(n_344), .B2(n_345), .C1(n_353), .C2(n_355), .Y(n_338) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g326 ( .A(n_265), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_265), .B(n_346), .Y(n_386) );
AND2x2_ASAP7_75t_L g397 ( .A(n_265), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g405 ( .A(n_268), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_270), .B(n_321), .Y(n_384) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_272), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g342 ( .A(n_272), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx3_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_275), .A2(n_378), .B(n_381), .C(n_383), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_275), .B(n_312), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_275), .B(n_295), .Y(n_417) );
AND2x2_ASAP7_75t_L g290 ( .A(n_276), .B(n_286), .Y(n_290) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g317 ( .A(n_279), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_280), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g369 ( .A(n_280), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g408 ( .A(n_280), .B(n_308), .Y(n_408) );
INVx1_ASAP7_75t_L g420 ( .A(n_280), .Y(n_420) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_283), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx1_ASAP7_75t_L g401 ( .A(n_286), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_291), .B(n_293), .C(n_297), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_289), .A2(n_319), .B1(n_334), .B2(n_337), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_290), .B(n_304), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_290), .B(n_312), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_291), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g354 ( .A(n_291), .Y(n_354) );
AND2x2_ASAP7_75t_L g361 ( .A(n_291), .B(n_341), .Y(n_361) );
INVx2_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NOR4xp25_ASAP7_75t_L g299 ( .A(n_296), .B(n_300), .C(n_301), .D(n_304), .Y(n_299) );
INVx1_ASAP7_75t_SL g370 ( .A(n_297), .Y(n_370) );
AND2x2_ASAP7_75t_L g414 ( .A(n_297), .B(n_415), .Y(n_414) );
OAI211xp5_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_306), .B(n_309), .C(n_318), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_305), .B(n_375), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_307), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_425) );
INVx1_ASAP7_75t_SL g380 ( .A(n_308), .Y(n_380) );
AND2x2_ASAP7_75t_L g419 ( .A(n_308), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_312), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_316), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_317), .B(n_342), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_324), .B(n_326), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g394 ( .A(n_321), .Y(n_394) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g422 ( .A(n_322), .Y(n_422) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_323), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B(n_333), .Y(n_328) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_329), .Y(n_341) );
OR2x2_ASAP7_75t_L g379 ( .A(n_329), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI21xp33_ASAP7_75t_SL g374 ( .A1(n_332), .A2(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_336), .A2(n_363), .B1(n_366), .B2(n_373), .C(n_374), .Y(n_362) );
INVx1_ASAP7_75t_SL g406 ( .A(n_337), .Y(n_406) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g353 ( .A(n_341), .B(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_350), .B2(n_351), .Y(n_345) );
INVx1_ASAP7_75t_L g385 ( .A(n_346), .Y(n_385) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_349), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR4xp25_ASAP7_75t_L g356 ( .A(n_357), .B(n_391), .C(n_404), .D(n_416), .Y(n_356) );
NAND3xp33_ASAP7_75t_SL g357 ( .A(n_358), .B(n_362), .C(n_377), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_360), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_367), .B(n_372), .Y(n_376) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_379), .A2(n_405), .B1(n_406), .B2(n_407), .C(n_409), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_381), .A2(n_396), .B(n_397), .C(n_399), .Y(n_395) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_382), .A2(n_400), .B1(n_402), .B2(n_403), .Y(n_399) );
INVx2_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_394), .C(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g410 ( .A(n_403), .Y(n_410) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI21xp5_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_411), .B(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B1(n_421), .B2(n_423), .C(n_425), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g443 ( .A1(n_431), .A2(n_444), .B1(n_712), .B2(n_714), .Y(n_443) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g440 ( .A(n_435), .Y(n_440) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_436), .B(n_713), .Y(n_720) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g712 ( .A(n_437), .B(n_713), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_439), .A2(n_442), .B(n_726), .Y(n_441) );
INVx1_ASAP7_75t_L g722 ( .A(n_444), .Y(n_722) );
NAND2x1_ASAP7_75t_L g444 ( .A(n_445), .B(n_628), .Y(n_444) );
NOR5xp2_ASAP7_75t_L g445 ( .A(n_446), .B(n_551), .C(n_583), .D(n_598), .E(n_615), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_479), .B(n_498), .C(n_539), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_460), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_448), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_448), .B(n_603), .Y(n_666) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_449), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_449), .B(n_495), .Y(n_552) );
AND2x2_ASAP7_75t_L g593 ( .A(n_449), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_449), .B(n_562), .Y(n_597) );
OR2x2_ASAP7_75t_L g634 ( .A(n_449), .B(n_485), .Y(n_634) );
INVx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g484 ( .A(n_450), .B(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g542 ( .A(n_450), .Y(n_542) );
OR2x2_ASAP7_75t_L g705 ( .A(n_450), .B(n_545), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_460), .A2(n_608), .B1(n_609), .B2(n_612), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_460), .B(n_542), .Y(n_691) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_470), .Y(n_460) );
AND2x2_ASAP7_75t_L g497 ( .A(n_461), .B(n_485), .Y(n_497) );
AND2x2_ASAP7_75t_L g544 ( .A(n_461), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g549 ( .A(n_461), .Y(n_549) );
INVx3_ASAP7_75t_L g562 ( .A(n_461), .Y(n_562) );
OR2x2_ASAP7_75t_L g582 ( .A(n_461), .B(n_545), .Y(n_582) );
AND2x2_ASAP7_75t_L g601 ( .A(n_461), .B(n_471), .Y(n_601) );
BUFx2_ASAP7_75t_L g633 ( .A(n_461), .Y(n_633) );
AND2x4_ASAP7_75t_L g548 ( .A(n_470), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g483 ( .A(n_471), .Y(n_483) );
INVx2_ASAP7_75t_L g496 ( .A(n_471), .Y(n_496) );
OR2x2_ASAP7_75t_L g564 ( .A(n_471), .B(n_545), .Y(n_564) );
AND2x2_ASAP7_75t_L g594 ( .A(n_471), .B(n_485), .Y(n_594) );
AND2x2_ASAP7_75t_L g611 ( .A(n_471), .B(n_542), .Y(n_611) );
AND2x2_ASAP7_75t_L g651 ( .A(n_471), .B(n_562), .Y(n_651) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_471), .B(n_497), .Y(n_687) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp33_ASAP7_75t_SL g480 ( .A(n_481), .B(n_494), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_482), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_483), .A2(n_497), .B(n_626), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_483), .B(n_485), .Y(n_681) );
AND2x2_ASAP7_75t_L g617 ( .A(n_484), .B(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g545 ( .A(n_485), .Y(n_545) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_485), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_494), .B(n_542), .Y(n_710) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_495), .A2(n_653), .B1(n_654), .B2(n_659), .Y(n_652) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
AND2x2_ASAP7_75t_L g543 ( .A(n_496), .B(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g581 ( .A(n_496), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g618 ( .A(n_496), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_497), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g672 ( .A(n_497), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_519), .Y(n_499) );
INVx4_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
AND2x2_ASAP7_75t_L g636 ( .A(n_500), .B(n_603), .Y(n_636) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
INVx3_ASAP7_75t_L g555 ( .A(n_501), .Y(n_555) );
AND2x2_ASAP7_75t_L g569 ( .A(n_501), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g573 ( .A(n_501), .Y(n_573) );
INVx2_ASAP7_75t_L g587 ( .A(n_501), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_501), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g644 ( .A(n_501), .B(n_639), .Y(n_644) );
AND2x2_ASAP7_75t_L g709 ( .A(n_501), .B(n_679), .Y(n_709) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .Y(n_501) );
AND2x2_ASAP7_75t_L g550 ( .A(n_510), .B(n_531), .Y(n_550) );
INVx2_ASAP7_75t_L g570 ( .A(n_510), .Y(n_570) );
INVx1_ASAP7_75t_L g575 ( .A(n_519), .Y(n_575) );
AND2x2_ASAP7_75t_L g621 ( .A(n_519), .B(n_569), .Y(n_621) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_530), .Y(n_519) );
INVx2_ASAP7_75t_L g560 ( .A(n_520), .Y(n_560) );
INVx1_ASAP7_75t_L g568 ( .A(n_520), .Y(n_568) );
AND2x2_ASAP7_75t_L g586 ( .A(n_520), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_520), .B(n_570), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
AND2x2_ASAP7_75t_L g603 ( .A(n_530), .B(n_560), .Y(n_603) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g556 ( .A(n_531), .Y(n_556) );
AND2x2_ASAP7_75t_L g639 ( .A(n_531), .B(n_570), .Y(n_639) );
OAI21xp5_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_546), .B(n_550), .Y(n_539) );
INVx1_ASAP7_75t_SL g584 ( .A(n_540), .Y(n_584) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_541), .B(n_548), .Y(n_641) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g590 ( .A(n_542), .B(n_545), .Y(n_590) );
AND2x2_ASAP7_75t_L g619 ( .A(n_542), .B(n_563), .Y(n_619) );
OR2x2_ASAP7_75t_L g622 ( .A(n_542), .B(n_582), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_543), .A2(n_635), .B1(n_687), .B2(n_688), .C1(n_690), .C2(n_692), .Y(n_686) );
BUFx2_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g589 ( .A(n_548), .B(n_590), .Y(n_589) );
INVx3_ASAP7_75t_SL g606 ( .A(n_548), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_548), .B(n_600), .Y(n_660) );
AND2x2_ASAP7_75t_L g595 ( .A(n_550), .B(n_555), .Y(n_595) );
INVx1_ASAP7_75t_L g614 ( .A(n_550), .Y(n_614) );
OAI221xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_553), .B1(n_557), .B2(n_561), .C(n_565), .Y(n_551) );
OR2x2_ASAP7_75t_L g623 ( .A(n_553), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g608 ( .A(n_555), .B(n_578), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_555), .B(n_568), .Y(n_648) );
AND2x2_ASAP7_75t_L g653 ( .A(n_555), .B(n_603), .Y(n_653) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_555), .Y(n_663) );
NAND2x1_ASAP7_75t_SL g674 ( .A(n_555), .B(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g559 ( .A(n_556), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g579 ( .A(n_556), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_556), .B(n_574), .Y(n_605) );
INVx1_ASAP7_75t_L g671 ( .A(n_556), .Y(n_671) );
INVx1_ASAP7_75t_L g646 ( .A(n_557), .Y(n_646) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g658 ( .A(n_558), .Y(n_658) );
NOR2xp67_ASAP7_75t_L g670 ( .A(n_558), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g675 ( .A(n_559), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_559), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g578 ( .A(n_560), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_560), .B(n_570), .Y(n_591) );
INVx1_ASAP7_75t_L g657 ( .A(n_560), .Y(n_657) );
INVx1_ASAP7_75t_L g678 ( .A(n_561), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_571), .B(n_580), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g711 ( .A(n_567), .B(n_644), .Y(n_711) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g679 ( .A(n_568), .B(n_639), .Y(n_679) );
AOI32xp33_ASAP7_75t_L g592 ( .A1(n_569), .A2(n_575), .A3(n_593), .B1(n_595), .B2(n_596), .Y(n_592) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_569), .A2(n_601), .A3(n_684), .B1(n_695), .B2(n_696), .C1(n_697), .C2(n_699), .Y(n_694) );
INVx2_ASAP7_75t_L g574 ( .A(n_570), .Y(n_574) );
INVx1_ASAP7_75t_L g684 ( .A(n_570), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_572), .B(n_578), .Y(n_627) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_573), .B(n_639), .Y(n_689) );
INVx1_ASAP7_75t_L g576 ( .A(n_574), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_574), .B(n_603), .Y(n_693) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_582), .B(n_677), .Y(n_676) );
OAI221xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_585), .B1(n_588), .B2(n_591), .C(n_592), .Y(n_583) );
OR2x2_ASAP7_75t_L g604 ( .A(n_585), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g613 ( .A(n_585), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g638 ( .A(n_586), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g642 ( .A(n_596), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B1(n_604), .B2(n_606), .C(n_607), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_600), .A2(n_631), .B1(n_635), .B2(n_636), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_601), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_601), .Y(n_706) );
INVx1_ASAP7_75t_L g700 ( .A(n_603), .Y(n_700) );
INVx1_ASAP7_75t_SL g635 ( .A(n_604), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_606), .B(n_634), .Y(n_696) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_611), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g677 ( .A(n_611), .Y(n_677) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_620), .B1(n_622), .B2(n_623), .C(n_625), .Y(n_615) );
NOR2xp33_ASAP7_75t_SL g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_617), .A2(n_635), .B1(n_681), .B2(n_682), .Y(n_680) );
CKINVDCx14_ASAP7_75t_R g620 ( .A(n_621), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g699 ( .A1(n_622), .A2(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR3xp33_ASAP7_75t_SL g628 ( .A(n_629), .B(n_661), .C(n_685), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g629 ( .A(n_630), .B(n_637), .C(n_645), .D(n_652), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g708 ( .A(n_633), .Y(n_708) );
INVx3_ASAP7_75t_SL g702 ( .A(n_634), .Y(n_702) );
OR2x2_ASAP7_75t_L g707 ( .A(n_634), .B(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B1(n_642), .B2(n_644), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_639), .B(n_657), .Y(n_698) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_647), .B(n_649), .Y(n_645) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g661 ( .A1(n_662), .A2(n_664), .B(n_667), .C(n_680), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g695 ( .A(n_666), .Y(n_695) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_672), .B1(n_673), .B2(n_676), .C1(n_678), .C2(n_679), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND4xp25_ASAP7_75t_SL g704 ( .A(n_677), .B(n_705), .C(n_706), .D(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND3xp33_ASAP7_75t_SL g685 ( .A(n_686), .B(n_694), .C(n_703), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_703) );
INVx1_ASAP7_75t_L g724 ( .A(n_714), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_715), .Y(n_725) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx3_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
endmodule