module fake_jpeg_1503_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_45),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g104 ( 
.A(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_58),
.Y(n_87)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

CKINVDCx9p33_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_52),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_53),
.Y(n_106)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_64),
.Y(n_105)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_34),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_74),
.Y(n_116)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_29),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_21),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_19),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_22),
.B(n_12),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_27),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_83),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_95),
.B1(n_56),
.B2(n_55),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_24),
.B1(n_16),
.B2(n_18),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_90),
.A2(n_111),
.B1(n_69),
.B2(n_46),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_83),
.B1(n_82),
.B2(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_99),
.B1(n_70),
.B2(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_94),
.B(n_96),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_42),
.B1(n_41),
.B2(n_37),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_18),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_24),
.B1(n_18),
.B2(n_16),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g175 ( 
.A1(n_100),
.A2(n_102),
.B(n_115),
.C(n_5),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_53),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_16),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_108),
.B(n_123),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_112),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_34),
.B1(n_27),
.B2(n_25),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_25),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_64),
.A2(n_39),
.B1(n_35),
.B2(n_32),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_23),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_23),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_21),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_51),
.B(n_19),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_63),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_19),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_136),
.B(n_149),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_138),
.A2(n_152),
.B1(n_105),
.B2(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_159),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_146),
.A2(n_153),
.B1(n_154),
.B2(n_165),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_46),
.B(n_29),
.C(n_48),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_147),
.A2(n_172),
.B(n_10),
.C(n_11),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_87),
.B(n_54),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_66),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_66),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_62),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_160),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_90),
.A2(n_62),
.B1(n_61),
.B2(n_60),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_61),
.B1(n_60),
.B2(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_0),
.Y(n_156)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_0),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_104),
.A2(n_0),
.B(n_1),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_0),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_1),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_167),
.Y(n_190)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

OAI22x1_ASAP7_75t_L g165 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_131),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_2),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_3),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_183),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_173),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_100),
.A2(n_3),
.B(n_5),
.C(n_7),
.Y(n_172)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_93),
.A2(n_102),
.B1(n_135),
.B2(n_92),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_185),
.B1(n_91),
.B2(n_113),
.Y(n_202)
);

NAND2x1_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_9),
.Y(n_222)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_178),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_7),
.B(n_8),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_179),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_120),
.B(n_7),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_181),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_118),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_91),
.B1(n_113),
.B2(n_119),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_92),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_116),
.B(n_114),
.C(n_125),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_188),
.B(n_182),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_105),
.B1(n_135),
.B2(n_84),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_198),
.B1(n_202),
.B2(n_208),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_152),
.A2(n_175),
.B1(n_140),
.B2(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_142),
.B(n_116),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_213),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_139),
.B(n_122),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_138),
.A2(n_124),
.B1(n_122),
.B2(n_89),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_228),
.B1(n_167),
.B2(n_147),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_141),
.B(n_89),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_219),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_137),
.B(n_97),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_175),
.A2(n_97),
.B1(n_101),
.B2(n_119),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_136),
.B(n_101),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_223),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_9),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_155),
.B(n_11),
.C(n_149),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_231),
.C(n_181),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_175),
.A2(n_11),
.B1(n_174),
.B2(n_161),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_145),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_175),
.A2(n_185),
.B1(n_165),
.B2(n_173),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_186),
.B(n_176),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_207),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_171),
.C(n_159),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_170),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_233),
.B(n_234),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_183),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_237),
.B1(n_241),
.B2(n_220),
.Y(n_272)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_167),
.B1(n_172),
.B2(n_166),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_144),
.B(n_157),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_238),
.A2(n_265),
.B(n_257),
.Y(n_301)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_242),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_187),
.B(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_262),
.B(n_215),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_196),
.B(n_158),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_254),
.B(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_248),
.A2(n_222),
.B(n_215),
.Y(n_281)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_200),
.B(n_164),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_253),
.B(n_217),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_196),
.B(n_179),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_216),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_193),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_205),
.B(n_204),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_260),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_195),
.B(n_221),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_187),
.A2(n_192),
.B(n_188),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_205),
.B(n_204),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_264),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_195),
.B(n_225),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_193),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_267),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_208),
.Y(n_266)
);

NOR2x1_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_222),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_223),
.B(n_188),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_209),
.B(n_215),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_199),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_210),
.C(n_209),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_275),
.C(n_297),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_272),
.A2(n_284),
.B1(n_300),
.B2(n_240),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_219),
.C(n_207),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_281),
.B(n_286),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_235),
.B1(n_241),
.B2(n_266),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_280),
.B1(n_285),
.B2(n_295),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_283),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_232),
.A2(n_228),
.B1(n_202),
.B2(n_191),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_234),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_248),
.A2(n_198),
.B1(n_211),
.B2(n_214),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_241),
.A2(n_237),
.B1(n_240),
.B2(n_243),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_261),
.A2(n_190),
.B(n_203),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_262),
.A2(n_211),
.B(n_190),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_294),
.B(n_298),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_301),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_268),
.A2(n_199),
.B(n_197),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_241),
.A2(n_189),
.B1(n_227),
.B2(n_197),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_267),
.A2(n_189),
.B(n_217),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_252),
.A2(n_212),
.B(n_227),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_247),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_238),
.A2(n_212),
.B1(n_255),
.B2(n_242),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_240),
.B1(n_251),
.B2(n_259),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_303),
.A2(n_305),
.B1(n_328),
.B2(n_279),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_280),
.A2(n_240),
.B1(n_263),
.B2(n_236),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_253),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_307),
.B(n_290),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_309),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_277),
.B(n_254),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_239),
.C(n_233),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_310),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_273),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_326),
.Y(n_349)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_239),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_314),
.C(n_319),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_264),
.C(n_247),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_290),
.B(n_244),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_316),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_246),
.C(n_249),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_327),
.B1(n_271),
.B2(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_272),
.A2(n_256),
.B1(n_260),
.B2(n_245),
.Y(n_328)
);

FAx1_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_304),
.CI(n_276),
.CON(n_329),
.SN(n_329)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_322),
.B(n_304),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_303),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_311),
.B1(n_285),
.B2(n_326),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_332),
.B1(n_334),
.B2(n_343),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_327),
.A2(n_292),
.B1(n_282),
.B2(n_271),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_269),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_337),
.B(n_347),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_320),
.C(n_315),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_293),
.C(n_274),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_348),
.C(n_319),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_302),
.A2(n_284),
.B1(n_300),
.B2(n_288),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_287),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_274),
.C(n_287),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_331),
.A2(n_302),
.B1(n_305),
.B2(n_328),
.Y(n_350)
);

OAI31xp33_ASAP7_75t_L g380 ( 
.A1(n_350),
.A2(n_358),
.A3(n_361),
.B(n_364),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_354),
.Y(n_375)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_349),
.Y(n_353)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_314),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_317),
.C(n_312),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_367),
.C(n_337),
.Y(n_376)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_349),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_363),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_359),
.B(n_362),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_344),
.A2(n_315),
.B1(n_325),
.B2(n_324),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_360),
.B(n_345),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_318),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_318),
.B1(n_292),
.B2(n_321),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_333),
.B(n_256),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_365),
.B(n_347),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g366 ( 
.A(n_329),
.B(n_294),
.CI(n_298),
.CON(n_366),
.SN(n_366)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_366),
.A2(n_338),
.B1(n_330),
.B2(n_346),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_289),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_358),
.A2(n_329),
.B(n_335),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_368),
.A2(n_370),
.B(n_372),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_366),
.A2(n_335),
.B(n_364),
.Y(n_370)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_373),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_374),
.B(n_342),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_378),
.C(n_381),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_355),
.A2(n_301),
.B(n_299),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_286),
.B(n_281),
.Y(n_379)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_379),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_362),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_386),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_375),
.B(n_354),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_383),
.B(n_388),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_380),
.B(n_351),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_352),
.C(n_367),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_352),
.C(n_370),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_391),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_387),
.A2(n_368),
.B(n_377),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_392),
.A2(n_394),
.B(n_398),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_369),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_389),
.C(n_384),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_387),
.A2(n_371),
.B(n_379),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_400),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_385),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_340),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_402),
.A2(n_396),
.B(n_397),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_401),
.B(n_384),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_404),
.Y(n_407)
);

OAI321xp33_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_341),
.A3(n_372),
.B1(n_366),
.B2(n_286),
.C(n_295),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_406),
.A2(n_403),
.B(n_341),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_407),
.Y(n_409)
);


endmodule