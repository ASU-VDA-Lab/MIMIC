module real_jpeg_29736_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx11_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_0),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_54),
.B1(n_61),
.B2(n_62),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_54),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_44),
.B1(n_45),
.B2(n_63),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_63),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_4),
.A2(n_33),
.B1(n_35),
.B2(n_63),
.Y(n_199)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_6),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_137),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_137),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_6),
.A2(n_33),
.B1(n_35),
.B2(n_137),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_51),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_8),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_186),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_186),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_186),
.Y(n_273)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_10),
.A2(n_38),
.B1(n_61),
.B2(n_62),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_38),
.B1(n_44),
.B2(n_45),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_11),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_165),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_165),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_11),
.A2(n_33),
.B1(n_35),
.B2(n_165),
.Y(n_265)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_48)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_13),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_14),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_57),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_14),
.B(n_44),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_14),
.A2(n_44),
.B(n_225),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_184),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_14),
.A2(n_30),
.B(n_33),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_14),
.B(n_133),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_14),
.A2(n_84),
.B1(n_158),
.B2(n_273),
.Y(n_275)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_114),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_113),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_20),
.B(n_97),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_81),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_21),
.A2(n_22),
.B1(n_71),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_69),
.B2(n_70),
.Y(n_22)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_24),
.A2(n_25),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_40),
.C(n_55),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_36),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_26),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_26),
.A2(n_32),
.B1(n_92),
.B2(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_26),
.A2(n_36),
.B(n_93),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_26),
.A2(n_32),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_26),
.A2(n_76),
.B(n_233),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_26),
.A2(n_32),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_26),
.A2(n_32),
.B1(n_232),
.B2(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_28),
.A2(n_45),
.A3(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g226 ( 
.A(n_29),
.B(n_223),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_29),
.A2(n_31),
.B(n_184),
.C(n_252),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_32),
.A2(n_78),
.B(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_32),
.B(n_184),
.Y(n_271)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_35),
.B(n_277),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_37),
.B(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B(n_52),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_41),
.A2(n_52),
.B(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_41),
.A2(n_107),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_48),
.B1(n_50),
.B2(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_42),
.B(n_53),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_42),
.A2(n_48),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_42),
.A2(n_48),
.B1(n_180),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_42),
.A2(n_48),
.B1(n_208),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_45),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_44),
.B(n_58),
.Y(n_197)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_45),
.A2(n_66),
.B1(n_183),
.B2(n_197),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_48),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_70),
.B1(n_99),
.B2(n_111),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_64),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_68),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_60),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_56),
.A2(n_101),
.B1(n_136),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_56),
.A2(n_101),
.B1(n_164),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_58),
.B(n_62),
.C(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_57),
.B(n_95),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_57),
.A2(n_65),
.B1(n_183),
.B2(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_62),
.Y(n_66)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g183 ( 
.A(n_62),
.B(n_184),
.CON(n_183),
.SN(n_183)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_109),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_82),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_90),
.B(n_94),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_94),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_83),
.A2(n_91),
.B1(n_120),
.B2(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B(n_88),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_84),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_84),
.A2(n_87),
.B1(n_155),
.B2(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_84),
.A2(n_129),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_84),
.A2(n_158),
.B1(n_265),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_85),
.A2(n_89),
.B(n_157),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_85),
.A2(n_86),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_89),
.Y(n_129)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_91),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_94),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_112),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_110),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_100),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_143),
.B(n_317),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_139),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_116),
.B(n_139),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_121),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_122),
.A2(n_123),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_132),
.C(n_134),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_125),
.B(n_130),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_126),
.A2(n_199),
.B(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_169),
.B(n_316),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_166),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_145),
.B(n_166),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_152),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_150),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_152),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.C(n_162),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_153),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_159),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_158),
.B(n_184),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_160),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_310),
.B(n_315),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_213),
.B(n_296),
.C(n_309),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_200),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_172),
.B(n_200),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_187),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_174),
.B(n_175),
.C(n_187),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_182),
.B(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_185),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_189),
.B(n_193),
.C(n_195),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.C(n_206),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_201),
.A2(n_202),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_206),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_211),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_295),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_288),
.B(n_294),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_243),
.B(n_287),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_234),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_217),
.B(n_234),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_227),
.C(n_230),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_218),
.A2(n_219),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_221),
.Y(n_241)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_235),
.B(n_241),
.C(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_281),
.B(n_286),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_261),
.B(n_280),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_246),
.B(n_253),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_251),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_258),
.C(n_259),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_260),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_269),
.B(n_279),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_267),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_274),
.B(n_278),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_290),
.Y(n_294)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_291),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_298),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_307),
.B2(n_308),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_304),
.C(n_308),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_307),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);


endmodule