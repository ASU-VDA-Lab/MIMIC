module fake_ibex_85_n_4595 (n_151, n_1084, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1079, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_1080, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_1077, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_343, n_310, n_714, n_1076, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_1075, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_1081, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_1083, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_1082, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_1089, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1078, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_1086, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_1087, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_1073, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_1085, n_361, n_455, n_419, n_774, n_72, n_1048, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_1088, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_4595);

input n_151;
input n_1084;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1079;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_1080;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_1077;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_343;
input n_310;
input n_714;
input n_1076;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_1075;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_1081;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_1083;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_1082;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_1089;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1078;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_1086;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_1087;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_1073;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_1085;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_1088;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_4595;

wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_2201;
wire n_1582;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_3319;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_4514;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_4372;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4353;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4343;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_4418;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_4403;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_2918;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1910;
wire n_2333;
wire n_1496;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3699;
wire n_1955;
wire n_3668;
wire n_4312;
wire n_4567;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_1326;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_4499;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_3777;
wire n_1799;
wire n_3293;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_4505;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3963;
wire n_3887;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4549;
wire n_4105;
wire n_4573;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4523;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3694;
wire n_3147;
wire n_2052;
wire n_3690;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_3448;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3634;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_1987;
wire n_4571;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4501;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_4230;
wire n_3849;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_4180;
wire n_4131;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_2063;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4485;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_3364;
wire n_1236;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_2080;
wire n_1477;
wire n_1184;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1990;
wire n_1179;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_3205;
wire n_3872;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_2935;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1566;
wire n_1464;
wire n_4362;
wire n_3568;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_4559;
wire n_1395;
wire n_1729;
wire n_1115;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_2197;
wire n_1523;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_4552;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_3719;
wire n_3390;
wire n_3948;
wire n_4425;
wire n_1599;
wire n_1806;
wire n_1539;
wire n_1400;
wire n_2711;
wire n_3070;
wire n_2842;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_3495;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_4117;
wire n_3999;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1683;
wire n_1185;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_3772;
wire n_2728;
wire n_2948;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_3955;
wire n_3867;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_4276;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_3902;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_4185;
wire n_2422;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_3784;
wire n_4142;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1694;
wire n_1458;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1858;
wire n_1537;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1962;
wire n_1225;
wire n_2346;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1860;
wire n_1491;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_4149;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_1396;
wire n_2916;
wire n_1923;
wire n_1224;
wire n_3206;
wire n_4021;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_3736;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_3162;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_4436;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_2059;
wire n_1278;
wire n_3276;
wire n_4366;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3959;
wire n_3743;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_2592;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1642;
wire n_1455;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_3273;
wire n_4367;
wire n_3139;
wire n_2700;
wire n_1222;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_4029;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1102;
wire n_3648;
wire n_3234;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_1275;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_4032;
wire n_3121;
wire n_2232;
wire n_2898;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_2278;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1809;
wire n_2367;
wire n_1206;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_1586;
wire n_1542;
wire n_1362;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3561;
wire n_2381;
wire n_2313;
wire n_3368;
wire n_3586;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_4555;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_4562;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_4281;
wire n_4345;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_3539;
wire n_1892;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_3989;
wire n_2119;
wire n_3844;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_4415;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1912;
wire n_1369;
wire n_1297;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_1285;
wire n_3042;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1824;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4528;
wire n_1486;
wire n_4363;
wire n_4502;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_4147;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_2005;
wire n_1284;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_2928;
wire n_3225;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_2169;
wire n_1398;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_4207;
wire n_4412;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_3286;
wire n_4038;
wire n_1092;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_4274;
wire n_4395;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_2148;
wire n_2104;
wire n_2303;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_3938;
wire n_4354;
wire n_4448;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_1450;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_3189;
wire n_2443;
wire n_3052;
wire n_4544;
wire n_2797;
wire n_2279;
wire n_1536;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_4275;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3550;
wire n_3261;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_1414;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_2619;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_4506;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_3792;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3988;
wire n_3758;
wire n_4327;
wire n_2656;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_3654;
wire n_3980;
wire n_2673;
wire n_2676;
wire n_2430;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_841),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_537),
.Y(n_1091)
);

CKINVDCx11_ASAP7_75t_R g1092 ( 
.A(n_142),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_683),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_163),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_185),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_189),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_337),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_602),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_544),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_495),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_787),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_187),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_977),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1043),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_871),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_92),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_607),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_583),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_559),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_256),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_628),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_698),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_832),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_457),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_824),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_288),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_839),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_447),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_85),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_203),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_610),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_656),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_657),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_216),
.Y(n_1124)
);

BUFx10_ASAP7_75t_L g1125 ( 
.A(n_115),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_131),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_823),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_431),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_737),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_110),
.Y(n_1130)
);

BUFx10_ASAP7_75t_L g1131 ( 
.A(n_671),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_554),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1041),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_949),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_522),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_843),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_813),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_380),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_9),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_71),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1009),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_248),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_136),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_861),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_620),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1026),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_1063),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_543),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_546),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_469),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_214),
.Y(n_1151)
);

BUFx2_ASAP7_75t_SL g1152 ( 
.A(n_452),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_209),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_858),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_433),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_306),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_324),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_914),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_941),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_101),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_330),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_134),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1071),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_852),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_791),
.Y(n_1165)
);

CKINVDCx16_ASAP7_75t_R g1166 ( 
.A(n_117),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_388),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_605),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_241),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1058),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_28),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_407),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_551),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1002),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1062),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_975),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_80),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_992),
.Y(n_1178)
);

BUFx2_ASAP7_75t_SL g1179 ( 
.A(n_261),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_427),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_202),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_173),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_1049),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_739),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_443),
.Y(n_1185)
);

BUFx5_ASAP7_75t_L g1186 ( 
.A(n_266),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1035),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_808),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_839),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_252),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_463),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_708),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_367),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_665),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_454),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_809),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_359),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_98),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_680),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_413),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_684),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_414),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_429),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_506),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_793),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_293),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_337),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_841),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_886),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_247),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1051),
.Y(n_1211)
);

CKINVDCx16_ASAP7_75t_R g1212 ( 
.A(n_874),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_918),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_455),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_782),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_194),
.Y(n_1216)
);

BUFx8_ASAP7_75t_SL g1217 ( 
.A(n_20),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1005),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_500),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_327),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_122),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1056),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_485),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_668),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_620),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_665),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_963),
.Y(n_1227)
);

CKINVDCx14_ASAP7_75t_R g1228 ( 
.A(n_563),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_715),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_31),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_525),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_480),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1045),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_199),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_87),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_553),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1088),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_22),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_689),
.Y(n_1239)
);

BUFx5_ASAP7_75t_L g1240 ( 
.A(n_466),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_696),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_342),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_876),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1033),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_939),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_768),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_894),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_128),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_430),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_243),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_151),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1003),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_112),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_470),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_580),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_221),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_873),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_769),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_172),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_270),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_242),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_239),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_233),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_136),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_8),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_186),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_141),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_69),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_38),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_259),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_369),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_444),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_137),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_619),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_677),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_490),
.Y(n_1276)
);

BUFx5_ASAP7_75t_L g1277 ( 
.A(n_493),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_544),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_301),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_317),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_283),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_39),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_945),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_373),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_561),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_659),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_659),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_94),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_150),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_244),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_755),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1044),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_250),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_914),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_562),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_157),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_805),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_535),
.Y(n_1298)
);

CKINVDCx14_ASAP7_75t_R g1299 ( 
.A(n_371),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_173),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_956),
.Y(n_1301)
);

BUFx5_ASAP7_75t_L g1302 ( 
.A(n_368),
.Y(n_1302)
);

CKINVDCx16_ASAP7_75t_R g1303 ( 
.A(n_784),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_138),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_810),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_403),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1000),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_729),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_286),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_185),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_692),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_703),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_698),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_443),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_891),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_538),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_314),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_989),
.Y(n_1318)
);

BUFx10_ASAP7_75t_L g1319 ( 
.A(n_1061),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_638),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1046),
.Y(n_1321)
);

BUFx10_ASAP7_75t_L g1322 ( 
.A(n_20),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_168),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_245),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_310),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_813),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1087),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1017),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_61),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_896),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_236),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_874),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_149),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_855),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_833),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1036),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_473),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_119),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_58),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_576),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_901),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_581),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_871),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_960),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1039),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_195),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_156),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_603),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_742),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_291),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_192),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_1001),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_652),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1006),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_916),
.Y(n_1355)
);

CKINVDCx14_ASAP7_75t_R g1356 ( 
.A(n_960),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_618),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_184),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_490),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_782),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1006),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1010),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_309),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1067),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_63),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_69),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_149),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_486),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_141),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_765),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_754),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_408),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_553),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_976),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_450),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1029),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_8),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_49),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_627),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_501),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_977),
.Y(n_1381)
);

CKINVDCx14_ASAP7_75t_R g1382 ( 
.A(n_762),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_51),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_240),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1050),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1011),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_463),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1041),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_566),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_391),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_398),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1057),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_505),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_314),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1059),
.Y(n_1395)
);

BUFx2_ASAP7_75t_SL g1396 ( 
.A(n_104),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_536),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_987),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_619),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_708),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_487),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_526),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_531),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_930),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_864),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_248),
.Y(n_1406)
);

BUFx10_ASAP7_75t_L g1407 ( 
.A(n_165),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1052),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_182),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_265),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_671),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_803),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_5),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_318),
.Y(n_1414)
);

BUFx10_ASAP7_75t_L g1415 ( 
.A(n_763),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_883),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_252),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1000),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_411),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_135),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_567),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1076),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_168),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_863),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_357),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_866),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_99),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_159),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_525),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1042),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_540),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_476),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_605),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_67),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_776),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_682),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_328),
.Y(n_1437)
);

BUFx10_ASAP7_75t_L g1438 ( 
.A(n_890),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_685),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_465),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_974),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_127),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_238),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_273),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_615),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_82),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1040),
.Y(n_1447)
);

BUFx10_ASAP7_75t_L g1448 ( 
.A(n_373),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1049),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1048),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_957),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_579),
.Y(n_1452)
);

CKINVDCx16_ASAP7_75t_R g1453 ( 
.A(n_794),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1062),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_450),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_628),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_889),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_856),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_224),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_448),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_125),
.Y(n_1461)
);

BUFx10_ASAP7_75t_L g1462 ( 
.A(n_425),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_348),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_272),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_87),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1054),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_571),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_235),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_730),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1038),
.Y(n_1470)
);

BUFx8_ASAP7_75t_SL g1471 ( 
.A(n_786),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_851),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_661),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_245),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1081),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_19),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_110),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_903),
.Y(n_1478)
);

BUFx5_ASAP7_75t_L g1479 ( 
.A(n_798),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_77),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_44),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_820),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_582),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1055),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1076),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_569),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_71),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_555),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1053),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_815),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_237),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_825),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_764),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_26),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_957),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_818),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_971),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_532),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_731),
.Y(n_1499)
);

BUFx10_ASAP7_75t_L g1500 ( 
.A(n_650),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_506),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_499),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_821),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1034),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_723),
.Y(n_1505)
);

CKINVDCx16_ASAP7_75t_R g1506 ( 
.A(n_870),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_259),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_753),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_871),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_108),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_32),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_872),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_346),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_188),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_923),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_769),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_323),
.Y(n_1517)
);

BUFx10_ASAP7_75t_L g1518 ( 
.A(n_283),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_899),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_88),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1001),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_112),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1060),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_456),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_234),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_958),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_890),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_92),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_342),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_115),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_559),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_864),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_375),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_419),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1039),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_260),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_845),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_294),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_535),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_367),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_332),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1037),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1047),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_249),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_2),
.Y(n_1545)
);

INVx4_ASAP7_75t_R g1546 ( 
.A(n_312),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_691),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_276),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_760),
.Y(n_1549)
);

BUFx5_ASAP7_75t_L g1550 ( 
.A(n_960),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_757),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_115),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_80),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_922),
.Y(n_1554)
);

BUFx5_ASAP7_75t_L g1555 ( 
.A(n_246),
.Y(n_1555)
);

CKINVDCx14_ASAP7_75t_R g1556 ( 
.A(n_360),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_993),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_766),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_359),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_258),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1085),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1016),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_739),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_172),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_735),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_53),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1077),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_326),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_319),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1049),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_825),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_251),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1064),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_382),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_823),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_194),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_43),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_296),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_347),
.Y(n_1579)
);

BUFx5_ASAP7_75t_L g1580 ( 
.A(n_1065),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_930),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1015),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_32),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_225),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_903),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_781),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1069),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_714),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_283),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_65),
.Y(n_1590)
);

BUFx10_ASAP7_75t_L g1591 ( 
.A(n_101),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_300),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_232),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_130),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_101),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_268),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_650),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_138),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1092),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1094),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1125),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1130),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1322),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1092),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1125),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1423),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1094),
.Y(n_1607)
);

CKINVDCx20_ASAP7_75t_R g1608 ( 
.A(n_1217),
.Y(n_1608)
);

INVx4_ASAP7_75t_R g1609 ( 
.A(n_1310),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1125),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1338),
.Y(n_1611)
);

INVxp33_ASAP7_75t_L g1612 ( 
.A(n_1217),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1228),
.Y(n_1613)
);

INVxp33_ASAP7_75t_SL g1614 ( 
.A(n_1261),
.Y(n_1614)
);

BUFx2_ASAP7_75t_SL g1615 ( 
.A(n_1407),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_1310),
.Y(n_1616)
);

CKINVDCx16_ASAP7_75t_R g1617 ( 
.A(n_1166),
.Y(n_1617)
);

INVxp33_ASAP7_75t_SL g1618 ( 
.A(n_1226),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1407),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1591),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1228),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1591),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1555),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1555),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1299),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1511),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1356),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1131),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1584),
.Y(n_1629)
);

CKINVDCx14_ASAP7_75t_R g1630 ( 
.A(n_1356),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1555),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1382),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1598),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1102),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1095),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1106),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1382),
.Y(n_1637)
);

INVxp67_ASAP7_75t_SL g1638 ( 
.A(n_1525),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1556),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1556),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1555),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1131),
.Y(n_1642)
);

INVxp33_ASAP7_75t_SL g1643 ( 
.A(n_1454),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1120),
.Y(n_1644)
);

CKINVDCx20_ASAP7_75t_R g1645 ( 
.A(n_1102),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1124),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1384),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1471),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1143),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1160),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1471),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1555),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1555),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1162),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1169),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1181),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1525),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1182),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1190),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1096),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1221),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1230),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_1590),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1248),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1265),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1594),
.Y(n_1666)
);

INVxp33_ASAP7_75t_SL g1667 ( 
.A(n_1119),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1090),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1329),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1186),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1234),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1331),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1333),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1358),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1377),
.Y(n_1675)
);

INVxp33_ASAP7_75t_SL g1676 ( 
.A(n_1126),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1268),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1383),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1406),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1428),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1459),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1461),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1474),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1476),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1186),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1139),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1140),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1142),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1480),
.Y(n_1689)
);

CKINVDCx14_ASAP7_75t_R g1690 ( 
.A(n_1131),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1186),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1186),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1276),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1481),
.Y(n_1694)
);

INVxp67_ASAP7_75t_SL g1695 ( 
.A(n_1210),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1487),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1520),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1530),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1186),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1268),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1544),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1545),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1296),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1157),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1564),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1577),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1151),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1595),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1576),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1258),
.Y(n_1710)
);

INVxp33_ASAP7_75t_SL g1711 ( 
.A(n_1153),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1215),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1210),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1171),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

OA21x2_ASAP7_75t_L g1716 ( 
.A1(n_1685),
.A2(n_1256),
.B(n_1251),
.Y(n_1716)
);

INVx4_ASAP7_75t_L g1717 ( 
.A(n_1628),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1606),
.B(n_1314),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1602),
.B(n_1335),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1623),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1616),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1641),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1693),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1602),
.B(n_1376),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1616),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1693),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1652),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1693),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1638),
.Y(n_1729)
);

OA21x2_ASAP7_75t_L g1730 ( 
.A1(n_1691),
.A2(n_1256),
.B(n_1251),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1653),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1642),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1606),
.B(n_1489),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1647),
.B(n_1557),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1638),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1635),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1636),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1642),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1644),
.A2(n_1572),
.B(n_1293),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1624),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1660),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_L g1742 ( 
.A(n_1613),
.B(n_1186),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1631),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1695),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1666),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1692),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_SL g1747 ( 
.A(n_1614),
.B(n_1667),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1699),
.A2(n_1572),
.B(n_1293),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1646),
.Y(n_1749)
);

INVx5_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1649),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1676),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1709),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1713),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1657),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1650),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1600),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1607),
.Y(n_1758)
);

OA21x2_ASAP7_75t_L g1759 ( 
.A1(n_1654),
.A2(n_1117),
.B(n_1100),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1655),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1656),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1663),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1711),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1658),
.A2(n_1117),
.B(n_1100),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1704),
.A2(n_1177),
.B1(n_1235),
.B2(n_1198),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1668),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1710),
.B(n_1238),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1659),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1714),
.Y(n_1769)
);

OA21x2_ASAP7_75t_L g1770 ( 
.A1(n_1661),
.A2(n_1144),
.B(n_1138),
.Y(n_1770)
);

INVx3_ASAP7_75t_L g1771 ( 
.A(n_1603),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1686),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1605),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1662),
.Y(n_1774)
);

BUFx6f_ASAP7_75t_L g1775 ( 
.A(n_1664),
.Y(n_1775)
);

AND2x6_ASAP7_75t_L g1776 ( 
.A(n_1610),
.B(n_1098),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1626),
.B(n_1098),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1634),
.A2(n_1109),
.B1(n_1132),
.B2(n_1108),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1615),
.B(n_1319),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1665),
.A2(n_1144),
.B(n_1138),
.Y(n_1780)
);

INVx6_ASAP7_75t_L g1781 ( 
.A(n_1618),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1669),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1672),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1673),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1687),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1611),
.B(n_1196),
.Y(n_1786)
);

BUFx8_ASAP7_75t_SL g1787 ( 
.A(n_1645),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1674),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1688),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1619),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1620),
.B(n_1622),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1675),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1678),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1629),
.B(n_1319),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1679),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1633),
.B(n_1183),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1680),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1681),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1682),
.Y(n_1799)
);

OA21x2_ASAP7_75t_L g1800 ( 
.A1(n_1683),
.A2(n_1203),
.B(n_1158),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1684),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1689),
.B(n_1250),
.Y(n_1802)
);

OA21x2_ASAP7_75t_L g1803 ( 
.A1(n_1694),
.A2(n_1203),
.B(n_1158),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1621),
.B(n_1625),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1696),
.Y(n_1805)
);

INVx6_ASAP7_75t_L g1806 ( 
.A(n_1643),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1697),
.Y(n_1807)
);

INVx5_ASAP7_75t_L g1808 ( 
.A(n_1609),
.Y(n_1808)
);

AND2x6_ASAP7_75t_L g1809 ( 
.A(n_1698),
.B(n_1183),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1701),
.B(n_1253),
.Y(n_1810)
);

INVx4_ASAP7_75t_L g1811 ( 
.A(n_1707),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1702),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1630),
.B(n_1212),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1705),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1706),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1708),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1627),
.B(n_1259),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1599),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1632),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1604),
.Y(n_1820)
);

INVx5_ASAP7_75t_L g1821 ( 
.A(n_1612),
.Y(n_1821)
);

BUFx2_ASAP7_75t_L g1822 ( 
.A(n_1637),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1639),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1640),
.B(n_1229),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1648),
.B(n_1262),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1651),
.Y(n_1826)
);

CKINVDCx14_ASAP7_75t_R g1827 ( 
.A(n_1671),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1677),
.Y(n_1828)
);

OA21x2_ASAP7_75t_L g1829 ( 
.A1(n_1700),
.A2(n_1275),
.B(n_1214),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1703),
.B(n_1303),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1628),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1628),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_1634),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1628),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1617),
.A2(n_1263),
.B1(n_1266),
.B2(n_1264),
.Y(n_1835)
);

BUFx8_ASAP7_75t_SL g1836 ( 
.A(n_1608),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1635),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1606),
.B(n_1362),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1616),
.Y(n_1839)
);

CKINVDCx11_ASAP7_75t_R g1840 ( 
.A(n_1608),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_L g1841 ( 
.A(n_1628),
.B(n_1362),
.Y(n_1841)
);

OA21x2_ASAP7_75t_L g1842 ( 
.A1(n_1685),
.A2(n_1275),
.B(n_1214),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1693),
.Y(n_1843)
);

CKINVDCx11_ASAP7_75t_R g1844 ( 
.A(n_1608),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1635),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1670),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1616),
.Y(n_1847)
);

BUFx6f_ASAP7_75t_L g1848 ( 
.A(n_1693),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1606),
.B(n_1371),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1693),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1685),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1685),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1685),
.Y(n_1853)
);

OAI22x1_ASAP7_75t_R g1854 ( 
.A1(n_1634),
.A2(n_1109),
.B1(n_1132),
.B2(n_1108),
.Y(n_1854)
);

BUFx6f_ASAP7_75t_L g1855 ( 
.A(n_1693),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1635),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1616),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1616),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1606),
.B(n_1269),
.Y(n_1859)
);

BUFx8_ASAP7_75t_L g1860 ( 
.A(n_1668),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1628),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1606),
.B(n_1426),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1616),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1670),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1693),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1693),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1628),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1635),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1614),
.A2(n_1514),
.B1(n_1453),
.B2(n_1506),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1670),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1628),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1690),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1693),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1670),
.Y(n_1874)
);

OA21x2_ASAP7_75t_L g1875 ( 
.A1(n_1685),
.A2(n_1350),
.B(n_1315),
.Y(n_1875)
);

OA21x2_ASAP7_75t_L g1876 ( 
.A1(n_1685),
.A2(n_1350),
.B(n_1315),
.Y(n_1876)
);

INVx5_ASAP7_75t_L g1877 ( 
.A(n_1628),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1606),
.B(n_1426),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1616),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1616),
.Y(n_1880)
);

INVx5_ASAP7_75t_L g1881 ( 
.A(n_1628),
.Y(n_1881)
);

OAI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1636),
.A2(n_1395),
.B(n_1354),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1693),
.Y(n_1883)
);

INVxp33_ASAP7_75t_SL g1884 ( 
.A(n_1647),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1693),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1670),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1616),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1628),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1606),
.B(n_1282),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1670),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1693),
.Y(n_1891)
);

AND2x6_ASAP7_75t_L g1892 ( 
.A(n_1601),
.B(n_1534),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1837),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1802),
.B(n_1288),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1837),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1845),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1845),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1882),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1736),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1754),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1856),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_R g1902 ( 
.A(n_1872),
.B(n_1593),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1868),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1739),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1787),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1717),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1836),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1840),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1844),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1753),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_R g1911 ( 
.A(n_1827),
.B(n_1136),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1759),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1884),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1797),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1833),
.Y(n_1915)
);

AOI21x1_ASAP7_75t_L g1916 ( 
.A1(n_1764),
.A2(n_1093),
.B(n_1091),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1860),
.Y(n_1917)
);

CKINVDCx16_ASAP7_75t_R g1918 ( 
.A(n_1752),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1810),
.B(n_1290),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1814),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1763),
.Y(n_1921)
);

BUFx3_ASAP7_75t_L g1922 ( 
.A(n_1745),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1779),
.Y(n_1923)
);

CKINVDCx20_ASAP7_75t_R g1924 ( 
.A(n_1745),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_1772),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1772),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1762),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1785),
.Y(n_1928)
);

BUFx10_ASAP7_75t_L g1929 ( 
.A(n_1781),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_R g1930 ( 
.A(n_1826),
.B(n_1149),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1764),
.Y(n_1931)
);

CKINVDCx20_ASAP7_75t_R g1932 ( 
.A(n_1854),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1781),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1770),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1780),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1766),
.Y(n_1936)
);

BUFx10_ASAP7_75t_L g1937 ( 
.A(n_1806),
.Y(n_1937)
);

INVxp67_ASAP7_75t_SL g1938 ( 
.A(n_1780),
.Y(n_1938)
);

CKINVDCx20_ASAP7_75t_R g1939 ( 
.A(n_1806),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1800),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1794),
.B(n_1300),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1778),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1835),
.Y(n_1943)
);

BUFx10_ASAP7_75t_L g1944 ( 
.A(n_1734),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1803),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1803),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1765),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1794),
.B(n_1304),
.Y(n_1948)
);

BUFx10_ASAP7_75t_L g1949 ( 
.A(n_1804),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1741),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1811),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1769),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1842),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1818),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1808),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1842),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1875),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1820),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1820),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1721),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1725),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_1869),
.Y(n_1962)
);

CKINVDCx20_ASAP7_75t_R g1963 ( 
.A(n_1822),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1729),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1875),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_1822),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1823),
.Y(n_1967)
);

CKINVDCx20_ASAP7_75t_R g1968 ( 
.A(n_1823),
.Y(n_1968)
);

NAND2x1_ASAP7_75t_L g1969 ( 
.A(n_1809),
.B(n_1546),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1735),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_R g1971 ( 
.A(n_1789),
.B(n_1149),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1732),
.B(n_1116),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1716),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1821),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1821),
.Y(n_1975)
);

CKINVDCx5p33_ASAP7_75t_R g1976 ( 
.A(n_1828),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1771),
.Y(n_1977)
);

AND3x2_ASAP7_75t_L g1978 ( 
.A(n_1719),
.B(n_1724),
.C(n_1813),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1817),
.B(n_1323),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1859),
.B(n_1324),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1876),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1718),
.Y(n_1982)
);

BUFx8_ASAP7_75t_L g1983 ( 
.A(n_1733),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1747),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_1825),
.Y(n_1985)
);

CKINVDCx20_ASAP7_75t_R g1986 ( 
.A(n_1889),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1767),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1716),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1839),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1819),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1847),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1830),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1838),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1730),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_R g1995 ( 
.A(n_1809),
.B(n_1218),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_R g1996 ( 
.A(n_1809),
.B(n_1218),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1857),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1748),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1858),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1849),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1862),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1863),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1878),
.Y(n_2003)
);

NAND2xp33_ASAP7_75t_R g2004 ( 
.A(n_1829),
.B(n_1339),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1750),
.Y(n_2005)
);

CKINVDCx20_ASAP7_75t_R g2006 ( 
.A(n_1829),
.Y(n_2006)
);

BUFx10_ASAP7_75t_L g2007 ( 
.A(n_1824),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1879),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1880),
.Y(n_2009)
);

CKINVDCx20_ASAP7_75t_R g2010 ( 
.A(n_1786),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1777),
.B(n_1796),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_R g2012 ( 
.A(n_1790),
.B(n_1742),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1887),
.Y(n_2013)
);

NOR2xp67_ASAP7_75t_L g2014 ( 
.A(n_1877),
.B(n_0),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1757),
.Y(n_2015)
);

CKINVDCx20_ASAP7_75t_R g2016 ( 
.A(n_1877),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1758),
.Y(n_2017)
);

CKINVDCx20_ASAP7_75t_R g2018 ( 
.A(n_1881),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1776),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1776),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1773),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_R g2022 ( 
.A(n_1738),
.B(n_1239),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1892),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1892),
.Y(n_2024)
);

CKINVDCx20_ASAP7_75t_R g2025 ( 
.A(n_1881),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1737),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1892),
.Y(n_2027)
);

CKINVDCx20_ASAP7_75t_R g2028 ( 
.A(n_1755),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1831),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1832),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1834),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1861),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1867),
.Y(n_2033)
);

NAND2xp33_ASAP7_75t_R g2034 ( 
.A(n_1871),
.B(n_1346),
.Y(n_2034)
);

NOR2x1p5_ASAP7_75t_L g2035 ( 
.A(n_1888),
.B(n_1347),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1805),
.B(n_1352),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1791),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1749),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1749),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_R g2040 ( 
.A(n_1783),
.B(n_1239),
.Y(n_2040)
);

AND3x2_ASAP7_75t_L g2041 ( 
.A(n_1783),
.B(n_1246),
.C(n_1245),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1751),
.Y(n_2042)
);

INVx3_ASAP7_75t_L g2043 ( 
.A(n_1751),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1756),
.Y(n_2044)
);

BUFx10_ASAP7_75t_L g2045 ( 
.A(n_1756),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1760),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1761),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_1768),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1768),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_1774),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1775),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1782),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1784),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_SL g2054 ( 
.A(n_1784),
.B(n_1351),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1795),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1795),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1799),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1799),
.Y(n_2058)
);

CKINVDCx20_ASAP7_75t_R g2059 ( 
.A(n_1801),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1816),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1816),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1812),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1841),
.A2(n_1395),
.B(n_1354),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1792),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1793),
.Y(n_2065)
);

INVxp67_ASAP7_75t_SL g2066 ( 
.A(n_1788),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1798),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1807),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1815),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1851),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_1851),
.A2(n_1853),
.B(n_1852),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_1852),
.Y(n_2072)
);

CKINVDCx16_ASAP7_75t_R g2073 ( 
.A(n_1853),
.Y(n_2073)
);

INVxp67_ASAP7_75t_L g2074 ( 
.A(n_1746),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_R g2075 ( 
.A(n_1740),
.B(n_1246),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1743),
.Y(n_2076)
);

NOR2xp67_ASAP7_75t_L g2077 ( 
.A(n_1723),
.B(n_1),
.Y(n_2077)
);

BUFx2_ASAP7_75t_L g2078 ( 
.A(n_1715),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1846),
.B(n_1352),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_SL g2080 ( 
.A1(n_1864),
.A2(n_1342),
.B1(n_1419),
.B2(n_1270),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1870),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1720),
.Y(n_2082)
);

AND2x6_ASAP7_75t_L g2083 ( 
.A(n_1874),
.B(n_1534),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1722),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1886),
.Y(n_2085)
);

CKINVDCx16_ASAP7_75t_R g2086 ( 
.A(n_1890),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1727),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_1731),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1726),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_1726),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1728),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1728),
.B(n_1352),
.Y(n_2092)
);

AND3x1_ASAP7_75t_L g2093 ( 
.A(n_1843),
.B(n_1342),
.C(n_1270),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1843),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_1848),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1848),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1850),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1891),
.Y(n_2098)
);

CKINVDCx20_ASAP7_75t_R g2099 ( 
.A(n_1855),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1865),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1866),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1873),
.Y(n_2102)
);

CKINVDCx20_ASAP7_75t_R g2103 ( 
.A(n_1873),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1883),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1885),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1885),
.B(n_1365),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1744),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1837),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_1929),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_1987),
.B(n_1165),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2037),
.B(n_1366),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2066),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2071),
.Y(n_2113)
);

OAI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2073),
.A2(n_1498),
.B1(n_1517),
.B2(n_1419),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1999),
.Y(n_2115)
);

CKINVDCx20_ASAP7_75t_R g2116 ( 
.A(n_1893),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_1923),
.B(n_1129),
.Y(n_2117)
);

NAND3x1_ASAP7_75t_L g2118 ( 
.A(n_1932),
.B(n_1517),
.C(n_1498),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_1901),
.B(n_1527),
.Y(n_2119)
);

NAND2xp33_ASAP7_75t_L g2120 ( 
.A(n_1950),
.B(n_1367),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_1899),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_1895),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_1896),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1912),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1922),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1894),
.B(n_1378),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_1897),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1927),
.Y(n_2128)
);

INVxp33_ASAP7_75t_L g2129 ( 
.A(n_2075),
.Y(n_2129)
);

BUFx10_ASAP7_75t_L g2130 ( 
.A(n_1917),
.Y(n_2130)
);

AND2x6_ASAP7_75t_L g2131 ( 
.A(n_1960),
.B(n_1538),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1931),
.Y(n_2132)
);

BUFx2_ASAP7_75t_L g2133 ( 
.A(n_2108),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1919),
.B(n_1409),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_2064),
.B(n_1413),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1900),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2072),
.B(n_1417),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1913),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2107),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1973),
.Y(n_2140)
);

AND3x4_ASAP7_75t_L g2141 ( 
.A(n_1908),
.B(n_1585),
.C(n_1579),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2079),
.B(n_1420),
.Y(n_2142)
);

INVx5_ASAP7_75t_L g2143 ( 
.A(n_2045),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_2006),
.A2(n_1396),
.B1(n_1538),
.B2(n_1579),
.Y(n_2144)
);

INVxp33_ASAP7_75t_L g2145 ( 
.A(n_2040),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1961),
.Y(n_2146)
);

BUFx10_ASAP7_75t_L g2147 ( 
.A(n_1909),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_1924),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1964),
.Y(n_2149)
);

AND2x6_ASAP7_75t_L g2150 ( 
.A(n_1970),
.B(n_1276),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1937),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1973),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1934),
.Y(n_2153)
);

INVx6_ASAP7_75t_L g2154 ( 
.A(n_1937),
.Y(n_2154)
);

AND2x6_ASAP7_75t_L g2155 ( 
.A(n_1989),
.B(n_1276),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1991),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1973),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_2065),
.B(n_1427),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_1921),
.B(n_1585),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1997),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_L g2161 ( 
.A(n_2045),
.Y(n_2161)
);

INVx2_ASAP7_75t_SL g2162 ( 
.A(n_1944),
.Y(n_2162)
);

AND2x6_ASAP7_75t_L g2163 ( 
.A(n_2002),
.B(n_1276),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1935),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2008),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2009),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2013),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2062),
.B(n_1434),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2067),
.B(n_1442),
.Y(n_2169)
);

CKINVDCx14_ASAP7_75t_R g2170 ( 
.A(n_1930),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1940),
.Y(n_2171)
);

AND2x6_ASAP7_75t_L g2172 ( 
.A(n_2069),
.B(n_1387),
.Y(n_2172)
);

BUFx2_ASAP7_75t_L g2173 ( 
.A(n_2022),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2021),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2076),
.B(n_1443),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_1963),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1944),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1945),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_2068),
.B(n_1903),
.Y(n_2179)
);

NOR2x1p5_ASAP7_75t_L g2180 ( 
.A(n_1905),
.B(n_1446),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2082),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_1985),
.B(n_1307),
.Y(n_2182)
);

BUFx6f_ASAP7_75t_L g2183 ( 
.A(n_1955),
.Y(n_2183)
);

BUFx3_ASAP7_75t_L g2184 ( 
.A(n_2103),
.Y(n_2184)
);

BUFx8_ASAP7_75t_SL g2185 ( 
.A(n_1907),
.Y(n_2185)
);

BUFx2_ASAP7_75t_L g2186 ( 
.A(n_1968),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1946),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1988),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1951),
.B(n_1465),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2084),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_2007),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2084),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1994),
.Y(n_2193)
);

AND2x4_ASAP7_75t_SL g2194 ( 
.A(n_2059),
.B(n_1415),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2070),
.Y(n_2195)
);

INVx3_ASAP7_75t_L g2196 ( 
.A(n_1949),
.Y(n_2196)
);

NOR3xp33_ASAP7_75t_L g2197 ( 
.A(n_2080),
.B(n_1539),
.C(n_1421),
.Y(n_2197)
);

BUFx3_ASAP7_75t_L g2198 ( 
.A(n_1939),
.Y(n_2198)
);

BUFx6f_ASAP7_75t_L g2199 ( 
.A(n_1998),
.Y(n_2199)
);

BUFx6f_ASAP7_75t_L g2200 ( 
.A(n_2050),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2078),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2063),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1904),
.Y(n_2203)
);

INVxp67_ASAP7_75t_L g2204 ( 
.A(n_2034),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_1941),
.B(n_1470),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1953),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1977),
.B(n_1468),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_1949),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_2007),
.Y(n_2209)
);

INVx2_ASAP7_75t_SL g2210 ( 
.A(n_1983),
.Y(n_2210)
);

CKINVDCx16_ASAP7_75t_R g2211 ( 
.A(n_1902),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_1948),
.B(n_1986),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_2035),
.B(n_1170),
.Y(n_2213)
);

OR2x6_ASAP7_75t_L g2214 ( 
.A(n_1969),
.B(n_1152),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_1918),
.B(n_1353),
.Y(n_2215)
);

BUFx2_ASAP7_75t_L g2216 ( 
.A(n_2093),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1982),
.B(n_1560),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_1925),
.B(n_1444),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2074),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1956),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1957),
.Y(n_2221)
);

BUFx10_ASAP7_75t_L g2222 ( 
.A(n_1933),
.Y(n_2222)
);

BUFx3_ASAP7_75t_L g2223 ( 
.A(n_1983),
.Y(n_2223)
);

AND2x6_ASAP7_75t_L g2224 ( 
.A(n_1965),
.B(n_1387),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1914),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1926),
.B(n_1596),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2015),
.A2(n_1491),
.B1(n_1510),
.B2(n_1477),
.Y(n_2227)
);

INVx1_ASAP7_75t_SL g2228 ( 
.A(n_1928),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_2017),
.B(n_1099),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1981),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_2016),
.Y(n_2231)
);

INVx5_ASAP7_75t_L g2232 ( 
.A(n_2083),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1920),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_1980),
.A2(n_1979),
.B1(n_1947),
.B2(n_1972),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_2090),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_2091),
.Y(n_2236)
);

BUFx6f_ASAP7_75t_L g2237 ( 
.A(n_2095),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2092),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1898),
.Y(n_2239)
);

CKINVDCx20_ASAP7_75t_R g2240 ( 
.A(n_1911),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2086),
.B(n_1101),
.Y(n_2241)
);

NOR2x1p5_ASAP7_75t_L g2242 ( 
.A(n_1966),
.B(n_1522),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_1910),
.B(n_1906),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_2018),
.Y(n_2244)
);

INVx2_ASAP7_75t_SL g2245 ( 
.A(n_1995),
.Y(n_2245)
);

OR2x2_ASAP7_75t_L g2246 ( 
.A(n_1952),
.B(n_1484),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2085),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2014),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1915),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1906),
.B(n_1528),
.Y(n_2250)
);

AO22x2_ASAP7_75t_L g2251 ( 
.A1(n_1938),
.A2(n_1179),
.B1(n_1586),
.B2(n_1369),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1938),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_1990),
.B(n_1103),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2081),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2106),
.Y(n_2255)
);

BUFx3_ASAP7_75t_L g2256 ( 
.A(n_2025),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2011),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1916),
.Y(n_2258)
);

BUFx3_ASAP7_75t_L g2259 ( 
.A(n_1954),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_1974),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2043),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_1978),
.B(n_1176),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_1975),
.Y(n_2263)
);

BUFx2_ASAP7_75t_L g2264 ( 
.A(n_1996),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_2100),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_1967),
.B(n_1260),
.Y(n_2266)
);

AND2x2_ASAP7_75t_SL g2267 ( 
.A(n_2041),
.B(n_1401),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_1993),
.B(n_1104),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1943),
.B(n_1438),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_2102),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2083),
.Y(n_2271)
);

OR2x6_ASAP7_75t_L g2272 ( 
.A(n_1958),
.B(n_1271),
.Y(n_2272)
);

AOI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_2083),
.A2(n_2028),
.B1(n_2054),
.B2(n_1978),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2019),
.B(n_1552),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2005),
.B(n_1309),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_1959),
.Y(n_2276)
);

INVx3_ASAP7_75t_L g2277 ( 
.A(n_2038),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2087),
.B(n_1553),
.Y(n_2278)
);

INVx2_ASAP7_75t_SL g2279 ( 
.A(n_2039),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_2088),
.B(n_1547),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2083),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2046),
.B(n_1566),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_2020),
.B(n_1289),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2048),
.B(n_2049),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2029),
.B(n_1097),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2023),
.B(n_1105),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2083),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2042),
.Y(n_2288)
);

NAND3x1_ASAP7_75t_L g2289 ( 
.A(n_1942),
.B(n_1112),
.C(n_1110),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2000),
.B(n_1438),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2001),
.B(n_1107),
.Y(n_2291)
);

AND2x6_ASAP7_75t_L g2292 ( 
.A(n_2043),
.B(n_2044),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_2003),
.B(n_1111),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2047),
.Y(n_2294)
);

BUFx2_ASAP7_75t_L g2295 ( 
.A(n_2051),
.Y(n_2295)
);

CKINVDCx16_ASAP7_75t_R g2296 ( 
.A(n_1962),
.Y(n_2296)
);

BUFx4f_ASAP7_75t_L g2297 ( 
.A(n_2057),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_2104),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_2052),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2026),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2030),
.B(n_1448),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2010),
.B(n_1113),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2053),
.B(n_1114),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2055),
.B(n_1115),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_2056),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2058),
.B(n_1118),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_2105),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1976),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_1984),
.B(n_1121),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2031),
.B(n_1448),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_2060),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_SL g2312 ( 
.A(n_2024),
.B(n_1122),
.Y(n_2312)
);

OR2x2_ASAP7_75t_L g2313 ( 
.A(n_1992),
.B(n_1123),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2061),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2077),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2032),
.B(n_1135),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_2033),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2012),
.B(n_1137),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2027),
.B(n_1462),
.Y(n_2319)
);

INVx4_ASAP7_75t_L g2320 ( 
.A(n_2089),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2089),
.Y(n_2321)
);

BUFx6f_ASAP7_75t_L g2322 ( 
.A(n_2089),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2004),
.B(n_1462),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_2094),
.Y(n_2324)
);

INVx1_ASAP7_75t_SL g2325 ( 
.A(n_2096),
.Y(n_2325)
);

INVx2_ASAP7_75t_SL g2326 ( 
.A(n_2097),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2101),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2098),
.B(n_1462),
.Y(n_2328)
);

BUFx3_ASAP7_75t_L g2329 ( 
.A(n_2099),
.Y(n_2329)
);

AND2x6_ASAP7_75t_L g2330 ( 
.A(n_2036),
.B(n_1387),
.Y(n_2330)
);

INVx2_ASAP7_75t_SL g2331 ( 
.A(n_1929),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_L g2332 ( 
.A1(n_2006),
.A2(n_1518),
.B1(n_1500),
.B2(n_1216),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_1922),
.B(n_1141),
.Y(n_2333)
);

INVx1_ASAP7_75t_SL g2334 ( 
.A(n_1893),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2071),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2066),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1922),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2037),
.B(n_1146),
.Y(n_2338)
);

BUFx4f_ASAP7_75t_L g2339 ( 
.A(n_1936),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2066),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_1899),
.B(n_1147),
.Y(n_2341)
);

AND2x6_ASAP7_75t_L g2342 ( 
.A(n_2036),
.B(n_1387),
.Y(n_2342)
);

BUFx10_ASAP7_75t_L g2343 ( 
.A(n_1917),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_1901),
.B(n_1500),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2071),
.Y(n_2345)
);

INVx4_ASAP7_75t_L g2346 ( 
.A(n_1899),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2066),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2066),
.Y(n_2348)
);

BUFx2_ASAP7_75t_L g2349 ( 
.A(n_1893),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_1971),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2071),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_1929),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2066),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2071),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2071),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2071),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2071),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2066),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2037),
.B(n_1154),
.Y(n_2359)
);

NAND2x1p5_ASAP7_75t_L g2360 ( 
.A(n_1922),
.B(n_1127),
.Y(n_2360)
);

AND2x6_ASAP7_75t_L g2361 ( 
.A(n_2036),
.B(n_1399),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_1899),
.B(n_1155),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2071),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_1899),
.B(n_1156),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2071),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2066),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2066),
.Y(n_2367)
);

AND3x2_ASAP7_75t_L g2368 ( 
.A(n_1936),
.B(n_1133),
.C(n_1128),
.Y(n_2368)
);

OR2x2_ASAP7_75t_L g2369 ( 
.A(n_1899),
.B(n_1164),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2037),
.A2(n_1172),
.B1(n_1173),
.B2(n_1168),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_1922),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_2099),
.Y(n_2372)
);

INVx4_ASAP7_75t_SL g2373 ( 
.A(n_1922),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_2099),
.Y(n_2374)
);

AND2x4_ASAP7_75t_L g2375 ( 
.A(n_1923),
.B(n_1134),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2066),
.Y(n_2376)
);

INVxp33_ASAP7_75t_L g2377 ( 
.A(n_1901),
.Y(n_2377)
);

AO22x2_ASAP7_75t_L g2378 ( 
.A1(n_1938),
.A2(n_1148),
.B1(n_1150),
.B2(n_1145),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2112),
.B(n_1174),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2128),
.B(n_1175),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2197),
.A2(n_1518),
.B1(n_1180),
.B2(n_1184),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_2339),
.B(n_1185),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2360),
.B(n_1187),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_2143),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2377),
.B(n_1188),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2143),
.B(n_1189),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2190),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2192),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2252),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2110),
.B(n_1193),
.Y(n_2390)
);

A2O1A1Ixp33_ASAP7_75t_L g2391 ( 
.A1(n_2126),
.A2(n_1408),
.B(n_1431),
.C(n_1401),
.Y(n_2391)
);

OAI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2132),
.A2(n_1161),
.B(n_1159),
.Y(n_2392)
);

O2A1O1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2134),
.A2(n_1167),
.B(n_1178),
.C(n_1163),
.Y(n_2393)
);

NOR3xp33_ASAP7_75t_L g2394 ( 
.A(n_2182),
.B(n_1192),
.C(n_1191),
.Y(n_2394)
);

INVx1_ASAP7_75t_SL g2395 ( 
.A(n_2116),
.Y(n_2395)
);

CKINVDCx16_ASAP7_75t_R g2396 ( 
.A(n_2211),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2336),
.B(n_2340),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2153),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2111),
.B(n_1204),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2347),
.B(n_2348),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2164),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2121),
.B(n_1207),
.Y(n_2402)
);

OAI22xp5_ASAP7_75t_L g2403 ( 
.A1(n_2378),
.A2(n_2353),
.B1(n_2366),
.B2(n_2358),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2205),
.A2(n_1211),
.B1(n_1219),
.B2(n_1213),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2161),
.B(n_2125),
.Y(n_2405)
);

INVx3_ASAP7_75t_L g2406 ( 
.A(n_2161),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2334),
.B(n_1223),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2344),
.B(n_1225),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_2145),
.B(n_1227),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2367),
.B(n_1231),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2376),
.B(n_1233),
.Y(n_2411)
);

BUFx4_ASAP7_75t_L g2412 ( 
.A(n_2284),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2122),
.B(n_1237),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2136),
.Y(n_2414)
);

AOI22xp33_ASAP7_75t_L g2415 ( 
.A1(n_2267),
.A2(n_1242),
.B1(n_1243),
.B2(n_1241),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_2127),
.B(n_1244),
.Y(n_2416)
);

BUFx6f_ASAP7_75t_L g2417 ( 
.A(n_2140),
.Y(n_2417)
);

OAI21xp5_ASAP7_75t_L g2418 ( 
.A1(n_2171),
.A2(n_1195),
.B(n_1194),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2125),
.B(n_1249),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2139),
.B(n_1252),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2146),
.B(n_1254),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2269),
.B(n_1255),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2149),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2129),
.B(n_1257),
.Y(n_2424)
);

BUFx3_ASAP7_75t_L g2425 ( 
.A(n_2337),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2203),
.A2(n_1199),
.B(n_1197),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2178),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_SL g2428 ( 
.A1(n_2114),
.A2(n_2216),
.B1(n_2170),
.B2(n_2173),
.Y(n_2428)
);

AOI21xp5_ASAP7_75t_L g2429 ( 
.A1(n_2239),
.A2(n_1201),
.B(n_1200),
.Y(n_2429)
);

NOR2x1p5_ASAP7_75t_L g2430 ( 
.A(n_2223),
.B(n_1283),
.Y(n_2430)
);

AOI22xp33_ASAP7_75t_L g2431 ( 
.A1(n_2144),
.A2(n_1291),
.B1(n_1295),
.B2(n_1286),
.Y(n_2431)
);

INVx1_ASAP7_75t_SL g2432 ( 
.A(n_2246),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_SL g2433 ( 
.A(n_2130),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2156),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2349),
.B(n_1297),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2349),
.B(n_1298),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2160),
.B(n_1301),
.Y(n_2437)
);

OR2x2_ASAP7_75t_L g2438 ( 
.A(n_2148),
.B(n_1305),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2165),
.Y(n_2439)
);

OAI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2378),
.A2(n_1408),
.B1(n_1432),
.B2(n_1431),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_L g2441 ( 
.A(n_2228),
.B(n_1306),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2166),
.B(n_1311),
.Y(n_2442)
);

AND2x6_ASAP7_75t_SL g2443 ( 
.A(n_2159),
.B(n_1202),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2341),
.B(n_1313),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2167),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2362),
.B(n_1317),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2364),
.B(n_1318),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2218),
.B(n_1320),
.Y(n_2448)
);

INVx6_ASAP7_75t_L g2449 ( 
.A(n_2343),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_2369),
.B(n_1325),
.Y(n_2450)
);

BUFx5_ASAP7_75t_L g2451 ( 
.A(n_2224),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2123),
.Y(n_2452)
);

INVx2_ASAP7_75t_SL g2453 ( 
.A(n_2222),
.Y(n_2453)
);

NAND2x1p5_ASAP7_75t_L g2454 ( 
.A(n_2232),
.B(n_1399),
.Y(n_2454)
);

INVx8_ASAP7_75t_L g2455 ( 
.A(n_2131),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2375),
.B(n_2323),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2251),
.A2(n_1437),
.B1(n_1439),
.B2(n_1432),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2375),
.B(n_1330),
.Y(n_2458)
);

INVxp67_ASAP7_75t_L g2459 ( 
.A(n_2133),
.Y(n_2459)
);

NOR3xp33_ASAP7_75t_L g2460 ( 
.A(n_2179),
.B(n_1206),
.C(n_1205),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2371),
.B(n_1334),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2187),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2308),
.B(n_1343),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2333),
.B(n_1345),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2251),
.A2(n_1439),
.B1(n_1482),
.B2(n_1437),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2227),
.B(n_1349),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2137),
.B(n_1355),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2212),
.B(n_1357),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2174),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2142),
.B(n_1359),
.Y(n_2470)
);

AOI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_2229),
.A2(n_1363),
.B1(n_1364),
.B2(n_1361),
.Y(n_2471)
);

NOR3xp33_ASAP7_75t_L g2472 ( 
.A(n_2216),
.B(n_1209),
.C(n_1208),
.Y(n_2472)
);

AOI21xp5_ASAP7_75t_L g2473 ( 
.A1(n_2113),
.A2(n_1222),
.B(n_1220),
.Y(n_2473)
);

NAND3xp33_ASAP7_75t_L g2474 ( 
.A(n_2332),
.B(n_2248),
.C(n_2273),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2195),
.B(n_1368),
.Y(n_2475)
);

BUFx5_ASAP7_75t_L g2476 ( 
.A(n_2224),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_2338),
.B(n_1370),
.Y(n_2477)
);

OR2x2_ASAP7_75t_L g2478 ( 
.A(n_2226),
.B(n_1372),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2255),
.B(n_2370),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2188),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_2359),
.B(n_1375),
.Y(n_2481)
);

OAI22xp5_ASAP7_75t_SL g2482 ( 
.A1(n_2141),
.A2(n_2240),
.B1(n_2296),
.B2(n_2350),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2219),
.Y(n_2483)
);

AOI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_2302),
.A2(n_1385),
.B1(n_1386),
.B2(n_1381),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_L g2485 ( 
.A(n_2313),
.B(n_1391),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2168),
.B(n_1397),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2175),
.B(n_1400),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2238),
.B(n_1402),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2234),
.B(n_1404),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2311),
.B(n_1410),
.Y(n_2490)
);

AND2x4_ASAP7_75t_L g2491 ( 
.A(n_2373),
.B(n_1224),
.Y(n_2491)
);

INVxp67_ASAP7_75t_L g2492 ( 
.A(n_2176),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2257),
.B(n_1412),
.Y(n_2493)
);

BUFx5_ASAP7_75t_L g2494 ( 
.A(n_2224),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2115),
.B(n_1418),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2206),
.Y(n_2496)
);

OAI221xp5_ASAP7_75t_L g2497 ( 
.A1(n_2278),
.A2(n_1429),
.B1(n_1430),
.B2(n_1424),
.C(n_1422),
.Y(n_2497)
);

NOR2xp33_ASAP7_75t_L g2498 ( 
.A(n_2309),
.B(n_1440),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2207),
.B(n_1441),
.Y(n_2499)
);

OAI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2220),
.A2(n_1515),
.B1(n_1524),
.B2(n_1507),
.Y(n_2500)
);

AOI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2335),
.A2(n_1236),
.B(n_1232),
.Y(n_2501)
);

NOR2xp67_ASAP7_75t_L g2502 ( 
.A(n_2210),
.B(n_254),
.Y(n_2502)
);

BUFx3_ASAP7_75t_L g2503 ( 
.A(n_2184),
.Y(n_2503)
);

NOR3xp33_ASAP7_75t_L g2504 ( 
.A(n_2217),
.B(n_1589),
.C(n_1578),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2131),
.B(n_1449),
.Y(n_2505)
);

BUFx8_ASAP7_75t_L g2506 ( 
.A(n_2176),
.Y(n_2506)
);

NOR3xp33_ASAP7_75t_L g2507 ( 
.A(n_2253),
.B(n_1597),
.C(n_1247),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2247),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2201),
.Y(n_2509)
);

NAND2xp33_ASAP7_75t_L g2510 ( 
.A(n_2131),
.B(n_1478),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2280),
.B(n_1450),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2250),
.B(n_1452),
.Y(n_2512)
);

A2O1A1Ixp33_ASAP7_75t_L g2513 ( 
.A1(n_2225),
.A2(n_1567),
.B(n_1587),
.C(n_1524),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2280),
.B(n_1460),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2285),
.B(n_1463),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2221),
.B(n_1466),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2328),
.B(n_2262),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_2301),
.B(n_1469),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2310),
.B(n_1472),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2285),
.B(n_1473),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2230),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2117),
.B(n_1483),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2330),
.B(n_1488),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2135),
.B(n_1490),
.Y(n_2524)
);

OAI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2272),
.A2(n_1497),
.B1(n_1499),
.B2(n_1496),
.Y(n_2525)
);

AOI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2242),
.A2(n_2213),
.B1(n_2266),
.B2(n_2241),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2233),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2330),
.B(n_2342),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2330),
.B(n_1503),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2342),
.B(n_1508),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2361),
.B(n_2120),
.Y(n_2531)
);

INVx2_ASAP7_75t_SL g2532 ( 
.A(n_2329),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_2158),
.B(n_1516),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2254),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2202),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2290),
.B(n_1521),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_2282),
.B(n_1523),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2361),
.B(n_1529),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2361),
.B(n_1531),
.Y(n_2539)
);

NOR2xp67_ASAP7_75t_L g2540 ( 
.A(n_2138),
.B(n_254),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2243),
.B(n_1532),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2373),
.B(n_1533),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2243),
.B(n_1536),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_SL g2544 ( 
.A(n_2295),
.B(n_1537),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2288),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2345),
.Y(n_2546)
);

OAI22xp5_ASAP7_75t_SL g2547 ( 
.A1(n_2249),
.A2(n_1542),
.B1(n_1543),
.B2(n_1540),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_SL g2548 ( 
.A(n_2295),
.B(n_1554),
.Y(n_2548)
);

INVx3_ASAP7_75t_L g2549 ( 
.A(n_2232),
.Y(n_2549)
);

INVx5_ASAP7_75t_L g2550 ( 
.A(n_2172),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2294),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2368),
.B(n_1562),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_2235),
.B(n_1563),
.Y(n_2553)
);

INVx8_ASAP7_75t_L g2554 ( 
.A(n_2272),
.Y(n_2554)
);

NAND3xp33_ASAP7_75t_L g2555 ( 
.A(n_2315),
.B(n_1414),
.C(n_1399),
.Y(n_2555)
);

BUFx5_ASAP7_75t_L g2556 ( 
.A(n_2150),
.Y(n_2556)
);

NAND2x1p5_ASAP7_75t_L g2557 ( 
.A(n_2232),
.B(n_1399),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2169),
.B(n_1565),
.Y(n_2558)
);

BUFx6f_ASAP7_75t_L g2559 ( 
.A(n_2140),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2351),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2374),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2268),
.B(n_1568),
.Y(n_2562)
);

BUFx3_ASAP7_75t_L g2563 ( 
.A(n_2372),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2194),
.B(n_1571),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2291),
.B(n_1573),
.Y(n_2565)
);

INVxp67_ASAP7_75t_L g2566 ( 
.A(n_2186),
.Y(n_2566)
);

CKINVDCx11_ASAP7_75t_R g2567 ( 
.A(n_2147),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2213),
.B(n_2293),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2319),
.B(n_1575),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2152),
.Y(n_2570)
);

OAI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2354),
.A2(n_1587),
.B1(n_1456),
.B2(n_1457),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2327),
.Y(n_2572)
);

AOI22xp33_ASAP7_75t_L g2573 ( 
.A1(n_2264),
.A2(n_1582),
.B1(n_1588),
.B2(n_1581),
.Y(n_2573)
);

O2A1O1Ixp33_ASAP7_75t_L g2574 ( 
.A1(n_2303),
.A2(n_1274),
.B(n_1278),
.C(n_1272),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2214),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2304),
.B(n_1592),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2324),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2235),
.B(n_1216),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2306),
.B(n_1279),
.Y(n_2579)
);

OAI22xp5_ASAP7_75t_SL g2580 ( 
.A1(n_2186),
.A2(n_1281),
.B1(n_1284),
.B2(n_1280),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2204),
.B(n_1285),
.Y(n_2581)
);

AND2x4_ASAP7_75t_L g2582 ( 
.A(n_2307),
.B(n_1287),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2355),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2356),
.A2(n_1294),
.B(n_1292),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2200),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2152),
.Y(n_2586)
);

NOR3xp33_ASAP7_75t_L g2587 ( 
.A(n_2283),
.B(n_1312),
.C(n_1308),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2318),
.B(n_1316),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2200),
.Y(n_2589)
);

INVx2_ASAP7_75t_SL g2590 ( 
.A(n_2236),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2316),
.B(n_1321),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2189),
.B(n_1326),
.Y(n_2592)
);

OA22x2_ASAP7_75t_L g2593 ( 
.A1(n_2264),
.A2(n_1328),
.B1(n_1332),
.B2(n_1327),
.Y(n_2593)
);

INVx2_ASAP7_75t_SL g2594 ( 
.A(n_2237),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2275),
.B(n_1336),
.Y(n_2595)
);

OAI22xp33_ASAP7_75t_L g2596 ( 
.A1(n_2259),
.A2(n_1340),
.B1(n_1341),
.B2(n_1337),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2275),
.B(n_1344),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2198),
.B(n_1348),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2245),
.B(n_1360),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2314),
.B(n_1373),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2277),
.B(n_1374),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2162),
.B(n_1379),
.Y(n_2602)
);

OR2x6_ASAP7_75t_L g2603 ( 
.A(n_2231),
.B(n_1380),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2261),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2177),
.B(n_1388),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2299),
.B(n_1389),
.Y(n_2606)
);

AND2x6_ASAP7_75t_L g2607 ( 
.A(n_2157),
.B(n_1267),
.Y(n_2607)
);

OAI22xp33_ASAP7_75t_L g2608 ( 
.A1(n_2276),
.A2(n_1392),
.B1(n_1393),
.B2(n_1390),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2305),
.B(n_1394),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2317),
.A2(n_1277),
.B1(n_1302),
.B2(n_1240),
.Y(n_2610)
);

AOI22xp5_ASAP7_75t_L g2611 ( 
.A1(n_2289),
.A2(n_1403),
.B1(n_1405),
.B2(n_1398),
.Y(n_2611)
);

NAND3xp33_ASAP7_75t_L g2612 ( 
.A(n_2357),
.B(n_1456),
.C(n_1414),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2279),
.B(n_1411),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2265),
.B(n_1267),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2363),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2274),
.B(n_1416),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2365),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2300),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_SL g2619 ( 
.A(n_2270),
.B(n_1273),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2286),
.B(n_1425),
.Y(n_2620)
);

AOI22xp5_ASAP7_75t_L g2621 ( 
.A1(n_2118),
.A2(n_1435),
.B1(n_1436),
.B2(n_1433),
.Y(n_2621)
);

AOI221xp5_ASAP7_75t_L g2622 ( 
.A1(n_2191),
.A2(n_1445),
.B1(n_1455),
.B2(n_1451),
.C(n_1447),
.Y(n_2622)
);

AOI22xp5_ASAP7_75t_L g2623 ( 
.A1(n_2109),
.A2(n_1464),
.B1(n_1467),
.B2(n_1458),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2193),
.A2(n_1456),
.B1(n_1457),
.B2(n_1414),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_2270),
.B(n_1273),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2199),
.B(n_1475),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2196),
.B(n_1485),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_2208),
.B(n_1486),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2209),
.B(n_1492),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2180),
.A2(n_1277),
.B1(n_1302),
.B2(n_1240),
.Y(n_2630)
);

OAI21xp5_ASAP7_75t_L g2631 ( 
.A1(n_2258),
.A2(n_1495),
.B(n_1493),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2298),
.B(n_1273),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2297),
.B(n_1273),
.Y(n_2633)
);

AO221x1_ASAP7_75t_L g2634 ( 
.A1(n_2271),
.A2(n_1457),
.B1(n_1505),
.B2(n_1456),
.C(n_1414),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2271),
.B(n_1501),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2312),
.B(n_1502),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2331),
.B(n_1504),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2287),
.Y(n_2638)
);

INVxp67_ASAP7_75t_L g2639 ( 
.A(n_2151),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2325),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2352),
.B(n_1509),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2281),
.B(n_1512),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_2260),
.B(n_1513),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_L g2644 ( 
.A(n_2263),
.B(n_1526),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2281),
.B(n_1548),
.Y(n_2645)
);

INVx2_ASAP7_75t_SL g2646 ( 
.A(n_2244),
.Y(n_2646)
);

A2O1A1Ixp33_ASAP7_75t_L g2647 ( 
.A1(n_2326),
.A2(n_1551),
.B(n_1558),
.C(n_1549),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2320),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_SL g2649 ( 
.A(n_2183),
.B(n_2256),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_SL g2650 ( 
.A(n_2183),
.B(n_1494),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_L g2651 ( 
.A(n_2292),
.B(n_1559),
.Y(n_2651)
);

OR2x2_ASAP7_75t_L g2652 ( 
.A(n_2321),
.B(n_1561),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2292),
.B(n_1569),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2292),
.B(n_1570),
.Y(n_2654)
);

NAND2x1_ASAP7_75t_L g2655 ( 
.A(n_2150),
.B(n_1457),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2150),
.B(n_1479),
.Y(n_2656)
);

NOR3xp33_ASAP7_75t_L g2657 ( 
.A(n_2185),
.B(n_1277),
.C(n_1240),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2155),
.Y(n_2658)
);

NOR3x1_ASAP7_75t_L g2659 ( 
.A(n_2172),
.B(n_254),
.C(n_253),
.Y(n_2659)
);

OR2x2_ASAP7_75t_L g2660 ( 
.A(n_2155),
.B(n_253),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2163),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2163),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_L g2663 ( 
.A(n_2163),
.B(n_255),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_SL g2664 ( 
.A(n_2339),
.B(n_1494),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2252),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2373),
.B(n_255),
.Y(n_2666)
);

NOR3xp33_ASAP7_75t_L g2667 ( 
.A(n_2110),
.B(n_1277),
.C(n_1240),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2128),
.B(n_1550),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2339),
.B(n_1494),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2339),
.B(n_1494),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2128),
.B(n_1550),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2128),
.B(n_1550),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2252),
.Y(n_2673)
);

OR2x6_ASAP7_75t_L g2674 ( 
.A(n_2210),
.B(n_1535),
.Y(n_2674)
);

INVxp33_ASAP7_75t_L g2675 ( 
.A(n_2215),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2128),
.B(n_1550),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2128),
.B(n_1550),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2252),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2252),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2128),
.B(n_1550),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2128),
.B(n_1550),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2128),
.B(n_1580),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_SL g2683 ( 
.A(n_2339),
.B(n_1583),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_SL g2684 ( 
.A(n_2339),
.B(n_1583),
.Y(n_2684)
);

AOI22xp33_ASAP7_75t_L g2685 ( 
.A1(n_2197),
.A2(n_1302),
.B1(n_1479),
.B2(n_1277),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2339),
.B(n_1583),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2377),
.B(n_256),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2181),
.Y(n_2688)
);

OAI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2114),
.A2(n_1519),
.B1(n_1535),
.B2(n_1505),
.Y(n_2689)
);

OAI21xp33_ASAP7_75t_L g2690 ( 
.A1(n_2126),
.A2(n_1519),
.B(n_1505),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2119),
.B(n_1302),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2143),
.Y(n_2692)
);

OR2x6_ASAP7_75t_L g2693 ( 
.A(n_2210),
.B(n_1519),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2339),
.B(n_1479),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_L g2695 ( 
.A(n_2377),
.B(n_256),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2119),
.B(n_1479),
.Y(n_2696)
);

AOI22xp33_ASAP7_75t_L g2697 ( 
.A1(n_2197),
.A2(n_1580),
.B1(n_1479),
.B2(n_1535),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2119),
.B(n_1580),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2252),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2110),
.A2(n_1580),
.B1(n_1574),
.B2(n_1541),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2339),
.B(n_1580),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_SL g2702 ( 
.A(n_2339),
.B(n_1541),
.Y(n_2702)
);

AOI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2110),
.A2(n_1574),
.B1(n_1541),
.B2(n_258),
.Y(n_2703)
);

BUFx6f_ASAP7_75t_L g2704 ( 
.A(n_2322),
.Y(n_2704)
);

NOR2x2_ASAP7_75t_L g2705 ( 
.A(n_2272),
.B(n_1085),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2339),
.B(n_257),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2252),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2252),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2128),
.B(n_2),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2181),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_2197),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_2143),
.Y(n_2712)
);

INVx2_ASAP7_75t_SL g2713 ( 
.A(n_2154),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2252),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2110),
.A2(n_261),
.B1(n_262),
.B2(n_260),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2143),
.Y(n_2716)
);

AOI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2110),
.A2(n_261),
.B1(n_262),
.B2(n_260),
.Y(n_2717)
);

AND2x6_ASAP7_75t_SL g2718 ( 
.A(n_2159),
.B(n_3),
.Y(n_2718)
);

INVx2_ASAP7_75t_SL g2719 ( 
.A(n_2154),
.Y(n_2719)
);

CKINVDCx20_ASAP7_75t_R g2720 ( 
.A(n_2116),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2252),
.Y(n_2721)
);

NAND2xp33_ASAP7_75t_L g2722 ( 
.A(n_2322),
.B(n_4),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2128),
.B(n_4),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2128),
.B(n_4),
.Y(n_2724)
);

OR2x2_ASAP7_75t_L g2725 ( 
.A(n_2114),
.B(n_263),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2181),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2252),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2181),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_SL g2729 ( 
.A(n_2339),
.B(n_263),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2339),
.B(n_264),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2112),
.B(n_5),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2128),
.B(n_6),
.Y(n_2732)
);

INVx3_ASAP7_75t_L g2733 ( 
.A(n_2143),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2128),
.B(n_6),
.Y(n_2734)
);

AOI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2203),
.A2(n_6),
.B(n_7),
.Y(n_2735)
);

INVx2_ASAP7_75t_SL g2736 ( 
.A(n_2154),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2252),
.Y(n_2737)
);

AOI22xp33_ASAP7_75t_L g2738 ( 
.A1(n_2197),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2128),
.B(n_7),
.Y(n_2739)
);

NOR2xp33_ASAP7_75t_L g2740 ( 
.A(n_2377),
.B(n_264),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2181),
.Y(n_2741)
);

NAND3xp33_ASAP7_75t_L g2742 ( 
.A(n_2144),
.B(n_266),
.C(n_265),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2197),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2181),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2339),
.B(n_267),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2128),
.B(n_9),
.Y(n_2746)
);

INVx3_ASAP7_75t_L g2747 ( 
.A(n_2143),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2181),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2339),
.B(n_267),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2181),
.Y(n_2750)
);

OAI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2124),
.A2(n_10),
.B(n_11),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2128),
.B(n_10),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_SL g2753 ( 
.A(n_2252),
.B(n_268),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2128),
.B(n_11),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_SL g2755 ( 
.A(n_2339),
.B(n_268),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2128),
.B(n_11),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2128),
.B(n_12),
.Y(n_2757)
);

NOR2xp67_ASAP7_75t_L g2758 ( 
.A(n_2346),
.B(n_273),
.Y(n_2758)
);

INVx4_ASAP7_75t_L g2759 ( 
.A(n_2143),
.Y(n_2759)
);

AOI22xp33_ASAP7_75t_L g2760 ( 
.A1(n_2197),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2181),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_SL g2762 ( 
.A(n_2252),
.B(n_269),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2181),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2128),
.B(n_13),
.Y(n_2764)
);

AND2x6_ASAP7_75t_SL g2765 ( 
.A(n_2159),
.B(n_13),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2339),
.B(n_269),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2128),
.B(n_14),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2119),
.B(n_1076),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2373),
.B(n_269),
.Y(n_2769)
);

OAI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2124),
.A2(n_14),
.B(n_15),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2128),
.B(n_14),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_R g2772 ( 
.A(n_2116),
.B(n_15),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2128),
.B(n_15),
.Y(n_2773)
);

INVxp67_ASAP7_75t_L g2774 ( 
.A(n_2246),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2128),
.B(n_15),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_2339),
.B(n_271),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2119),
.B(n_1080),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_SL g2778 ( 
.A(n_2339),
.B(n_271),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2128),
.B(n_16),
.Y(n_2779)
);

NAND2xp33_ASAP7_75t_L g2780 ( 
.A(n_2322),
.B(n_16),
.Y(n_2780)
);

NOR2x1p5_ASAP7_75t_L g2781 ( 
.A(n_2223),
.B(n_272),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2128),
.B(n_16),
.Y(n_2782)
);

AND2x6_ASAP7_75t_L g2783 ( 
.A(n_2252),
.B(n_272),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2252),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2128),
.B(n_17),
.Y(n_2785)
);

INVx4_ASAP7_75t_L g2786 ( 
.A(n_2143),
.Y(n_2786)
);

INVx5_ASAP7_75t_L g2787 ( 
.A(n_2161),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2339),
.B(n_273),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2377),
.B(n_274),
.Y(n_2789)
);

OR2x2_ASAP7_75t_SL g2790 ( 
.A(n_2211),
.B(n_1086),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2128),
.B(n_18),
.Y(n_2791)
);

BUFx4f_ASAP7_75t_L g2792 ( 
.A(n_2210),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2181),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2128),
.B(n_19),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2128),
.B(n_19),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2181),
.Y(n_2796)
);

OR2x6_ASAP7_75t_L g2797 ( 
.A(n_2210),
.B(n_274),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2181),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_2128),
.B(n_20),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2252),
.A2(n_276),
.B1(n_277),
.B2(n_275),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_SL g2801 ( 
.A(n_2223),
.Y(n_2801)
);

AO221x1_ASAP7_75t_L g2802 ( 
.A1(n_2251),
.A2(n_278),
.B1(n_279),
.B2(n_277),
.C(n_275),
.Y(n_2802)
);

AOI22xp33_ASAP7_75t_L g2803 ( 
.A1(n_2197),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2803)
);

INVxp67_ASAP7_75t_L g2804 ( 
.A(n_2246),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_SL g2805 ( 
.A(n_2339),
.B(n_277),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2339),
.B(n_278),
.Y(n_2806)
);

AOI22xp33_ASAP7_75t_L g2807 ( 
.A1(n_2197),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2128),
.B(n_23),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2128),
.B(n_23),
.Y(n_2809)
);

NOR2x1_ASAP7_75t_L g2810 ( 
.A(n_2223),
.B(n_278),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2181),
.Y(n_2811)
);

O2A1O1Ixp33_ASAP7_75t_L g2812 ( 
.A1(n_2126),
.A2(n_280),
.B(n_281),
.C(n_279),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_L g2813 ( 
.A(n_2377),
.B(n_279),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_SL g2814 ( 
.A(n_2339),
.B(n_281),
.Y(n_2814)
);

INVx4_ASAP7_75t_L g2815 ( 
.A(n_2143),
.Y(n_2815)
);

NOR2x1p5_ASAP7_75t_L g2816 ( 
.A(n_2223),
.B(n_280),
.Y(n_2816)
);

OR2x2_ASAP7_75t_L g2817 ( 
.A(n_2114),
.B(n_280),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_SL g2818 ( 
.A(n_2339),
.B(n_284),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_SL g2819 ( 
.A(n_2339),
.B(n_284),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2181),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2181),
.Y(n_2821)
);

AOI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2110),
.A2(n_285),
.B1(n_286),
.B2(n_282),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2181),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2377),
.B(n_282),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2112),
.B(n_24),
.Y(n_2825)
);

NOR2xp33_ASAP7_75t_SL g2826 ( 
.A(n_2252),
.B(n_285),
.Y(n_2826)
);

AOI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2110),
.A2(n_287),
.B1(n_288),
.B2(n_286),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2112),
.B(n_24),
.Y(n_2828)
);

AOI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2612),
.A2(n_288),
.B(n_287),
.Y(n_2829)
);

NAND3xp33_ASAP7_75t_L g2830 ( 
.A(n_2457),
.B(n_289),
.C(n_287),
.Y(n_2830)
);

AOI21xp5_ASAP7_75t_L g2831 ( 
.A1(n_2612),
.A2(n_290),
.B(n_289),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2546),
.A2(n_291),
.B(n_290),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_R g2833 ( 
.A(n_2720),
.B(n_2567),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2432),
.B(n_2479),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2389),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2675),
.B(n_292),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2456),
.B(n_292),
.Y(n_2837)
);

O2A1O1Ixp33_ASAP7_75t_L g2838 ( 
.A1(n_2457),
.A2(n_295),
.B(n_296),
.C(n_293),
.Y(n_2838)
);

AND2x4_ASAP7_75t_L g2839 ( 
.A(n_2787),
.B(n_295),
.Y(n_2839)
);

AOI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2394),
.A2(n_297),
.B1(n_298),
.B2(n_295),
.Y(n_2840)
);

AOI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2560),
.A2(n_298),
.B(n_297),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2414),
.B(n_299),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_2753),
.B(n_300),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2665),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2583),
.A2(n_301),
.B(n_300),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2673),
.Y(n_2846)
);

AOI21xp5_ASAP7_75t_L g2847 ( 
.A1(n_2615),
.A2(n_303),
.B(n_302),
.Y(n_2847)
);

AOI21xp5_ASAP7_75t_L g2848 ( 
.A1(n_2617),
.A2(n_303),
.B(n_302),
.Y(n_2848)
);

OAI21xp33_ASAP7_75t_L g2849 ( 
.A1(n_2753),
.A2(n_24),
.B(n_25),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2678),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2509),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_2762),
.B(n_304),
.Y(n_2852)
);

OAI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2393),
.A2(n_24),
.B(n_25),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2568),
.B(n_304),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2535),
.A2(n_306),
.B(n_305),
.Y(n_2855)
);

AOI33xp33_ASAP7_75t_L g2856 ( 
.A1(n_2381),
.A2(n_308),
.A3(n_306),
.B1(n_309),
.B2(n_307),
.B3(n_305),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2762),
.B(n_307),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2571),
.A2(n_308),
.B(n_307),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2423),
.B(n_308),
.Y(n_2859)
);

OAI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2392),
.A2(n_25),
.B(n_26),
.Y(n_2860)
);

AND2x4_ASAP7_75t_L g2861 ( 
.A(n_2787),
.B(n_309),
.Y(n_2861)
);

BUFx4f_ASAP7_75t_L g2862 ( 
.A(n_2554),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2434),
.B(n_311),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2440),
.A2(n_312),
.B1(n_313),
.B2(n_311),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2679),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2690),
.A2(n_313),
.B(n_312),
.Y(n_2866)
);

INVx3_ASAP7_75t_L g2867 ( 
.A(n_2759),
.Y(n_2867)
);

AOI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2631),
.A2(n_316),
.B(n_315),
.Y(n_2868)
);

AOI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2668),
.A2(n_316),
.B(n_315),
.Y(n_2869)
);

INVx1_ASAP7_75t_SL g2870 ( 
.A(n_2412),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2671),
.A2(n_318),
.B(n_317),
.Y(n_2871)
);

BUFx2_ASAP7_75t_L g2872 ( 
.A(n_2693),
.Y(n_2872)
);

INVx3_ASAP7_75t_L g2873 ( 
.A(n_2786),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2387),
.Y(n_2874)
);

A2O1A1Ixp33_ASAP7_75t_L g2875 ( 
.A1(n_2574),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2672),
.A2(n_319),
.B(n_318),
.Y(n_2876)
);

AOI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_2676),
.A2(n_320),
.B(n_319),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2677),
.A2(n_321),
.B(n_320),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2680),
.A2(n_2682),
.B(n_2681),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2388),
.Y(n_2880)
);

AOI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2774),
.A2(n_321),
.B1(n_322),
.B2(n_320),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_2674),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2439),
.B(n_322),
.Y(n_2883)
);

AOI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2516),
.A2(n_2707),
.B(n_2699),
.Y(n_2884)
);

AO21x2_ASAP7_75t_L g2885 ( 
.A1(n_2634),
.A2(n_323),
.B(n_322),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2445),
.B(n_323),
.Y(n_2886)
);

A2O1A1Ixp33_ASAP7_75t_L g2887 ( 
.A1(n_2812),
.A2(n_30),
.B(n_27),
.C(n_29),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2516),
.A2(n_325),
.B(n_324),
.Y(n_2888)
);

OAI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2440),
.A2(n_325),
.B1(n_326),
.B2(n_324),
.Y(n_2889)
);

OAI21xp5_ASAP7_75t_L g2890 ( 
.A1(n_2418),
.A2(n_27),
.B(n_29),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2826),
.B(n_325),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2784),
.A2(n_2714),
.B(n_2708),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2721),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2727),
.Y(n_2894)
);

OAI21xp33_ASAP7_75t_L g2895 ( 
.A1(n_2465),
.A2(n_29),
.B(n_30),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2737),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2815),
.Y(n_2897)
);

AOI21xp5_ASAP7_75t_L g2898 ( 
.A1(n_2473),
.A2(n_328),
.B(n_327),
.Y(n_2898)
);

NAND2x1p5_ASAP7_75t_L g2899 ( 
.A(n_2787),
.B(n_328),
.Y(n_2899)
);

AOI21x1_ASAP7_75t_L g2900 ( 
.A1(n_2403),
.A2(n_330),
.B(n_329),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_SL g2901 ( 
.A(n_2525),
.B(n_329),
.Y(n_2901)
);

AOI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2804),
.A2(n_330),
.B1(n_331),
.B2(n_329),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2688),
.B(n_331),
.Y(n_2903)
);

AO21x1_ASAP7_75t_L g2904 ( 
.A1(n_2800),
.A2(n_2770),
.B(n_2751),
.Y(n_2904)
);

OR2x2_ASAP7_75t_L g2905 ( 
.A(n_2448),
.B(n_332),
.Y(n_2905)
);

INVxp67_ASAP7_75t_L g2906 ( 
.A(n_2797),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2710),
.B(n_333),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2501),
.A2(n_334),
.B(n_333),
.Y(n_2908)
);

AOI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2584),
.A2(n_334),
.B(n_333),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2492),
.B(n_2566),
.Y(n_2910)
);

HB1xp67_ASAP7_75t_L g2911 ( 
.A(n_2674),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2428),
.B(n_335),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2786),
.Y(n_2913)
);

O2A1O1Ixp33_ASAP7_75t_L g2914 ( 
.A1(n_2391),
.A2(n_336),
.B(n_337),
.C(n_335),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2693),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2726),
.B(n_2728),
.Y(n_2916)
);

AND2x4_ASAP7_75t_L g2917 ( 
.A(n_2815),
.B(n_338),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2741),
.B(n_338),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2744),
.B(n_339),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_L g2920 ( 
.A(n_2417),
.Y(n_2920)
);

A2O1A1Ixp33_ASAP7_75t_L g2921 ( 
.A1(n_2742),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2748),
.B(n_340),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2397),
.A2(n_341),
.B(n_340),
.Y(n_2923)
);

NAND2x1_ASAP7_75t_L g2924 ( 
.A(n_2607),
.B(n_2693),
.Y(n_2924)
);

OAI21xp33_ASAP7_75t_L g2925 ( 
.A1(n_2477),
.A2(n_31),
.B(n_32),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2750),
.B(n_341),
.Y(n_2926)
);

OAI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2652),
.A2(n_343),
.B1(n_344),
.B2(n_342),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2761),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2763),
.B(n_343),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2793),
.B(n_343),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2796),
.B(n_344),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2798),
.B(n_345),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2811),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2820),
.B(n_345),
.Y(n_2934)
);

OAI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2647),
.A2(n_33),
.B(n_34),
.Y(n_2935)
);

AOI21xp5_ASAP7_75t_L g2936 ( 
.A1(n_2400),
.A2(n_349),
.B(n_348),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2821),
.B(n_348),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2398),
.Y(n_2938)
);

OAI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2379),
.A2(n_33),
.B(n_34),
.Y(n_2939)
);

OR2x2_ASAP7_75t_L g2940 ( 
.A(n_2478),
.B(n_2395),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2797),
.A2(n_351),
.B1(n_352),
.B2(n_350),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_SL g2942 ( 
.A(n_2452),
.B(n_350),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2823),
.B(n_351),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2401),
.Y(n_2944)
);

AOI21xp5_ASAP7_75t_L g2945 ( 
.A1(n_2635),
.A2(n_352),
.B(n_351),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2459),
.B(n_352),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2635),
.A2(n_354),
.B(n_353),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2399),
.B(n_353),
.Y(n_2948)
);

OR2x6_ASAP7_75t_L g2949 ( 
.A(n_2554),
.B(n_355),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2469),
.B(n_355),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2588),
.A2(n_357),
.B(n_356),
.Y(n_2951)
);

INVx4_ASAP7_75t_L g2952 ( 
.A(n_2455),
.Y(n_2952)
);

BUFx6f_ASAP7_75t_L g2953 ( 
.A(n_2417),
.Y(n_2953)
);

AND2x4_ASAP7_75t_L g2954 ( 
.A(n_2384),
.B(n_356),
.Y(n_2954)
);

OAI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2379),
.A2(n_33),
.B(n_34),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2427),
.A2(n_359),
.B(n_358),
.Y(n_2956)
);

NOR3xp33_ASAP7_75t_L g2957 ( 
.A(n_2474),
.B(n_360),
.C(n_358),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2390),
.B(n_358),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2511),
.B(n_361),
.Y(n_2959)
);

AOI221x1_ASAP7_75t_L g2960 ( 
.A1(n_2800),
.A2(n_2667),
.B1(n_2770),
.B2(n_2624),
.C(n_2555),
.Y(n_2960)
);

INVx4_ASAP7_75t_L g2961 ( 
.A(n_2455),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2508),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2462),
.A2(n_363),
.B(n_362),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_SL g2964 ( 
.A(n_2758),
.B(n_364),
.Y(n_2964)
);

NOR3xp33_ASAP7_75t_L g2965 ( 
.A(n_2580),
.B(n_2565),
.C(n_2562),
.Y(n_2965)
);

O2A1O1Ixp33_ASAP7_75t_L g2966 ( 
.A1(n_2497),
.A2(n_365),
.B(n_366),
.C(n_364),
.Y(n_2966)
);

INVx2_ASAP7_75t_SL g2967 ( 
.A(n_2449),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2534),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2527),
.Y(n_2969)
);

AOI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2480),
.A2(n_365),
.B(n_364),
.Y(n_2970)
);

OR2x2_ASAP7_75t_L g2971 ( 
.A(n_2438),
.B(n_365),
.Y(n_2971)
);

O2A1O1Ixp5_ASAP7_75t_L g2972 ( 
.A1(n_2531),
.A2(n_368),
.B(n_369),
.C(n_366),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2514),
.B(n_2422),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2517),
.B(n_368),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_L g2975 ( 
.A(n_2464),
.B(n_369),
.Y(n_2975)
);

OAI21xp5_ASAP7_75t_L g2976 ( 
.A1(n_2512),
.A2(n_35),
.B(n_36),
.Y(n_2976)
);

AOI22xp5_ASAP7_75t_L g2977 ( 
.A1(n_2444),
.A2(n_371),
.B1(n_372),
.B2(n_370),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2515),
.B(n_370),
.Y(n_2978)
);

AOI21xp33_ASAP7_75t_L g2979 ( 
.A1(n_2485),
.A2(n_2498),
.B(n_2447),
.Y(n_2979)
);

BUFx6f_ASAP7_75t_L g2980 ( 
.A(n_2417),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_SL g2981 ( 
.A(n_2502),
.B(n_370),
.Y(n_2981)
);

INVx4_ASAP7_75t_L g2982 ( 
.A(n_2455),
.Y(n_2982)
);

BUFx6f_ASAP7_75t_L g2983 ( 
.A(n_2559),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2768),
.B(n_2777),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_SL g2985 ( 
.A(n_2554),
.B(n_373),
.Y(n_2985)
);

INVx4_ASAP7_75t_L g2986 ( 
.A(n_2433),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2496),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2521),
.Y(n_2988)
);

NOR2xp33_ASAP7_75t_L g2989 ( 
.A(n_2468),
.B(n_374),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2483),
.B(n_374),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2638),
.A2(n_375),
.B(n_374),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2731),
.Y(n_2992)
);

BUFx3_ASAP7_75t_L g2993 ( 
.A(n_2449),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2731),
.Y(n_2994)
);

AO21x1_ASAP7_75t_L g2995 ( 
.A1(n_2500),
.A2(n_2557),
.B(n_2454),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_SL g2996 ( 
.A(n_2640),
.B(n_375),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2408),
.B(n_376),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2518),
.B(n_376),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2691),
.B(n_377),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2696),
.B(n_377),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2825),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2579),
.A2(n_2591),
.B(n_2642),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2698),
.B(n_378),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2545),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2825),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2507),
.B(n_378),
.Y(n_3006)
);

AOI21x1_ASAP7_75t_L g3007 ( 
.A1(n_2626),
.A2(n_379),
.B(n_378),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2828),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2645),
.A2(n_380),
.B(n_379),
.Y(n_3009)
);

NAND3xp33_ASAP7_75t_L g3010 ( 
.A(n_2700),
.B(n_382),
.C(n_381),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2550),
.B(n_381),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2828),
.Y(n_3012)
);

O2A1O1Ixp33_ASAP7_75t_SL g3013 ( 
.A1(n_2578),
.A2(n_384),
.B(n_385),
.C(n_383),
.Y(n_3013)
);

A2O1A1Ixp33_ASAP7_75t_L g3014 ( 
.A1(n_2735),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2551),
.Y(n_3015)
);

HB1xp67_ASAP7_75t_L g3016 ( 
.A(n_2603),
.Y(n_3016)
);

NOR3xp33_ASAP7_75t_L g3017 ( 
.A(n_2706),
.B(n_384),
.C(n_383),
.Y(n_3017)
);

AOI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_2446),
.A2(n_384),
.B1(n_385),
.B2(n_383),
.Y(n_3018)
);

AOI21x1_ASAP7_75t_L g3019 ( 
.A1(n_2500),
.A2(n_386),
.B(n_385),
.Y(n_3019)
);

BUFx3_ASAP7_75t_L g3020 ( 
.A(n_2503),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2519),
.B(n_386),
.Y(n_3021)
);

OAI21xp33_ASAP7_75t_L g3022 ( 
.A1(n_2481),
.A2(n_36),
.B(n_37),
.Y(n_3022)
);

AOI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2722),
.A2(n_387),
.B(n_386),
.Y(n_3023)
);

AOI33xp33_ASAP7_75t_L g3024 ( 
.A1(n_2711),
.A2(n_390),
.A3(n_388),
.B1(n_391),
.B2(n_389),
.B3(n_387),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_SL g3025 ( 
.A(n_2550),
.B(n_2556),
.Y(n_3025)
);

AOI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2780),
.A2(n_388),
.B(n_387),
.Y(n_3026)
);

AOI21xp33_ASAP7_75t_L g3027 ( 
.A1(n_2450),
.A2(n_390),
.B(n_389),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_2426),
.A2(n_390),
.B(n_389),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2572),
.Y(n_3029)
);

OAI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2499),
.A2(n_38),
.B(n_39),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2431),
.B(n_391),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2622),
.B(n_392),
.Y(n_3032)
);

INVx5_ASAP7_75t_L g3033 ( 
.A(n_2607),
.Y(n_3033)
);

INVxp67_ASAP7_75t_L g3034 ( 
.A(n_2797),
.Y(n_3034)
);

A2O1A1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2429),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_3035)
);

OAI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_2611),
.A2(n_394),
.B1(n_395),
.B2(n_393),
.Y(n_3036)
);

AOI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_2559),
.A2(n_394),
.B(n_393),
.Y(n_3037)
);

NOR2xp67_ASAP7_75t_L g3038 ( 
.A(n_2692),
.B(n_394),
.Y(n_3038)
);

AOI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2520),
.A2(n_397),
.B1(n_398),
.B2(n_396),
.Y(n_3039)
);

AO21x1_ASAP7_75t_L g3040 ( 
.A1(n_2557),
.A2(n_400),
.B(n_399),
.Y(n_3040)
);

AOI21x1_ASAP7_75t_L g3041 ( 
.A1(n_2528),
.A2(n_2661),
.B(n_2658),
.Y(n_3041)
);

AOI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2570),
.A2(n_2586),
.B(n_2510),
.Y(n_3042)
);

AOI21x1_ASAP7_75t_L g3043 ( 
.A1(n_2651),
.A2(n_400),
.B(n_399),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2536),
.B(n_400),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2383),
.B(n_401),
.Y(n_3045)
);

HB1xp67_ASAP7_75t_L g3046 ( 
.A(n_2603),
.Y(n_3046)
);

OAI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2467),
.A2(n_41),
.B(n_42),
.Y(n_3047)
);

AOI21xp33_ASAP7_75t_L g3048 ( 
.A1(n_2575),
.A2(n_2505),
.B(n_2489),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2563),
.Y(n_3049)
);

O2A1O1Ixp33_ASAP7_75t_L g3050 ( 
.A1(n_2504),
.A2(n_403),
.B(n_404),
.C(n_402),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_2484),
.B(n_2435),
.Y(n_3051)
);

NOR3xp33_ASAP7_75t_L g3052 ( 
.A(n_2729),
.B(n_405),
.C(n_404),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2436),
.B(n_406),
.Y(n_3053)
);

INVx4_ASAP7_75t_L g3054 ( 
.A(n_2801),
.Y(n_3054)
);

BUFx6f_ASAP7_75t_L g3055 ( 
.A(n_2607),
.Y(n_3055)
);

INVx2_ASAP7_75t_SL g3056 ( 
.A(n_2792),
.Y(n_3056)
);

AOI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2709),
.A2(n_410),
.B(n_409),
.Y(n_3057)
);

AND2x4_ASAP7_75t_L g3058 ( 
.A(n_2692),
.B(n_409),
.Y(n_3058)
);

BUFx3_ASAP7_75t_L g3059 ( 
.A(n_2425),
.Y(n_3059)
);

CKINVDCx5p33_ASAP7_75t_R g3060 ( 
.A(n_2801),
.Y(n_3060)
);

O2A1O1Ixp33_ASAP7_75t_L g3061 ( 
.A1(n_2596),
.A2(n_414),
.B(n_415),
.C(n_412),
.Y(n_3061)
);

AOI21xp5_ASAP7_75t_L g3062 ( 
.A1(n_2723),
.A2(n_414),
.B(n_412),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2550),
.B(n_416),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2470),
.B(n_416),
.Y(n_3064)
);

NOR2xp67_ASAP7_75t_L g3065 ( 
.A(n_2712),
.B(n_416),
.Y(n_3065)
);

AOI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2724),
.A2(n_2734),
.B(n_2732),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2739),
.A2(n_418),
.B(n_417),
.Y(n_3067)
);

O2A1O1Ixp5_ASAP7_75t_L g3068 ( 
.A1(n_2614),
.A2(n_418),
.B(n_419),
.C(n_417),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_L g3069 ( 
.A(n_2413),
.B(n_418),
.Y(n_3069)
);

AND2x4_ASAP7_75t_L g3070 ( 
.A(n_2712),
.B(n_420),
.Y(n_3070)
);

O2A1O1Ixp33_ASAP7_75t_L g3071 ( 
.A1(n_2608),
.A2(n_2819),
.B(n_2818),
.C(n_2730),
.Y(n_3071)
);

OAI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2486),
.A2(n_41),
.B(n_42),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2460),
.B(n_421),
.Y(n_3073)
);

INVx3_ASAP7_75t_L g3074 ( 
.A(n_2716),
.Y(n_3074)
);

OAI21xp33_ASAP7_75t_L g3075 ( 
.A1(n_2599),
.A2(n_43),
.B(n_44),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_SL g3076 ( 
.A(n_2556),
.B(n_422),
.Y(n_3076)
);

AOI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2746),
.A2(n_423),
.B(n_422),
.Y(n_3077)
);

BUFx6f_ASAP7_75t_L g3078 ( 
.A(n_2704),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2752),
.A2(n_2809),
.B(n_2808),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2556),
.B(n_423),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2404),
.B(n_424),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2458),
.B(n_424),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2754),
.A2(n_2757),
.B(n_2756),
.Y(n_3083)
);

AOI21xp5_ASAP7_75t_L g3084 ( 
.A1(n_2764),
.A2(n_2771),
.B(n_2767),
.Y(n_3084)
);

OAI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2487),
.A2(n_43),
.B(n_44),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2716),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2493),
.B(n_425),
.Y(n_3087)
);

OAI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2703),
.A2(n_426),
.B1(n_427),
.B2(n_425),
.Y(n_3088)
);

AOI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2773),
.A2(n_427),
.B(n_426),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2775),
.A2(n_428),
.B(n_426),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_L g3091 ( 
.A(n_2704),
.Y(n_3091)
);

HB1xp67_ASAP7_75t_L g3092 ( 
.A(n_2783),
.Y(n_3092)
);

AOI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_2779),
.A2(n_429),
.B(n_428),
.Y(n_3093)
);

OAI21xp33_ASAP7_75t_L g3094 ( 
.A1(n_2613),
.A2(n_45),
.B(n_46),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2782),
.Y(n_3095)
);

AOI21xp5_ASAP7_75t_L g3096 ( 
.A1(n_2785),
.A2(n_429),
.B(n_428),
.Y(n_3096)
);

O2A1O1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2745),
.A2(n_431),
.B(n_432),
.C(n_430),
.Y(n_3097)
);

AOI21xp5_ASAP7_75t_L g3098 ( 
.A1(n_2791),
.A2(n_433),
.B(n_432),
.Y(n_3098)
);

HB1xp67_ASAP7_75t_L g3099 ( 
.A(n_2783),
.Y(n_3099)
);

INVx1_ASAP7_75t_SL g3100 ( 
.A(n_2542),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2600),
.B(n_434),
.Y(n_3101)
);

O2A1O1Ixp5_ASAP7_75t_L g3102 ( 
.A1(n_2619),
.A2(n_435),
.B(n_436),
.C(n_434),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_SL g3103 ( 
.A(n_2556),
.B(n_435),
.Y(n_3103)
);

AO21x1_ASAP7_75t_L g3104 ( 
.A1(n_2663),
.A2(n_438),
.B(n_437),
.Y(n_3104)
);

AND2x6_ASAP7_75t_L g3105 ( 
.A(n_2659),
.B(n_437),
.Y(n_3105)
);

O2A1O1Ixp33_ASAP7_75t_SL g3106 ( 
.A1(n_2625),
.A2(n_438),
.B(n_439),
.C(n_437),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2618),
.Y(n_3107)
);

OAI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2415),
.A2(n_439),
.B1(n_440),
.B2(n_438),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2738),
.B(n_439),
.Y(n_3109)
);

O2A1O1Ixp33_ASAP7_75t_SL g3110 ( 
.A1(n_2632),
.A2(n_441),
.B(n_442),
.C(n_440),
.Y(n_3110)
);

OAI22xp5_ASAP7_75t_L g3111 ( 
.A1(n_2725),
.A2(n_441),
.B1(n_442),
.B2(n_440),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_2733),
.B(n_441),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2743),
.B(n_442),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2760),
.B(n_443),
.Y(n_3114)
);

OAI21xp33_ASAP7_75t_L g3115 ( 
.A1(n_2643),
.A2(n_45),
.B(n_46),
.Y(n_3115)
);

INVx3_ASAP7_75t_L g3116 ( 
.A(n_2733),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2794),
.A2(n_445),
.B(n_444),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2795),
.A2(n_445),
.B(n_444),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2799),
.A2(n_447),
.B(n_446),
.Y(n_3119)
);

BUFx2_ASAP7_75t_SL g3120 ( 
.A(n_2430),
.Y(n_3120)
);

OAI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_2817),
.A2(n_448),
.B1(n_449),
.B2(n_446),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2416),
.B(n_448),
.Y(n_3122)
);

NOR3xp33_ASAP7_75t_L g3123 ( 
.A(n_2749),
.B(n_451),
.C(n_449),
.Y(n_3123)
);

HB1xp67_ASAP7_75t_L g3124 ( 
.A(n_2783),
.Y(n_3124)
);

INVxp67_ASAP7_75t_SL g3125 ( 
.A(n_2704),
.Y(n_3125)
);

AOI21x1_ASAP7_75t_L g3126 ( 
.A1(n_2653),
.A2(n_452),
.B(n_451),
.Y(n_3126)
);

INVx2_ASAP7_75t_SL g3127 ( 
.A(n_2792),
.Y(n_3127)
);

OAI21xp33_ASAP7_75t_L g3128 ( 
.A1(n_2644),
.A2(n_46),
.B(n_47),
.Y(n_3128)
);

OAI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2715),
.A2(n_454),
.B1(n_455),
.B2(n_453),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_L g3130 ( 
.A(n_2441),
.B(n_453),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2747),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2803),
.B(n_455),
.Y(n_3132)
);

AOI21x1_ASAP7_75t_L g3133 ( 
.A1(n_2654),
.A2(n_457),
.B(n_456),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2807),
.B(n_456),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2582),
.B(n_457),
.Y(n_3135)
);

NAND3xp33_ASAP7_75t_L g3136 ( 
.A(n_2630),
.B(n_459),
.C(n_458),
.Y(n_3136)
);

INVx4_ASAP7_75t_L g3137 ( 
.A(n_2783),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2488),
.B(n_458),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2689),
.B(n_459),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2601),
.Y(n_3140)
);

AND2x4_ASAP7_75t_L g3141 ( 
.A(n_2406),
.B(n_460),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2581),
.B(n_460),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2537),
.A2(n_462),
.B(n_461),
.Y(n_3143)
);

NAND3xp33_ASAP7_75t_L g3144 ( 
.A(n_2657),
.B(n_463),
.C(n_462),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2623),
.B(n_462),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2380),
.B(n_464),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_2547),
.B(n_2472),
.Y(n_3147)
);

BUFx6f_ASAP7_75t_L g3148 ( 
.A(n_2648),
.Y(n_3148)
);

OAI22xp5_ASAP7_75t_L g3149 ( 
.A1(n_2717),
.A2(n_467),
.B1(n_468),
.B2(n_466),
.Y(n_3149)
);

AOI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_2555),
.A2(n_2475),
.B(n_2513),
.Y(n_3150)
);

AOI21xp33_ASAP7_75t_L g3151 ( 
.A1(n_2605),
.A2(n_467),
.B(n_466),
.Y(n_3151)
);

INVx1_ASAP7_75t_SL g3152 ( 
.A(n_2406),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_L g3153 ( 
.A(n_2407),
.B(n_467),
.Y(n_3153)
);

AOI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_2576),
.A2(n_469),
.B(n_468),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2569),
.B(n_2561),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2420),
.B(n_469),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2421),
.A2(n_471),
.B(n_470),
.Y(n_3157)
);

O2A1O1Ixp5_ASAP7_75t_L g3158 ( 
.A1(n_2405),
.A2(n_471),
.B(n_472),
.C(n_470),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2437),
.A2(n_472),
.B(n_471),
.Y(n_3159)
);

OR2x6_ASAP7_75t_L g3160 ( 
.A(n_2781),
.B(n_472),
.Y(n_3160)
);

HB1xp67_ASAP7_75t_L g3161 ( 
.A(n_2506),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2442),
.B(n_473),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2604),
.A2(n_475),
.B(n_474),
.Y(n_3163)
);

AOI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_2656),
.A2(n_475),
.B(n_474),
.Y(n_3164)
);

AO21x1_ASAP7_75t_L g3165 ( 
.A1(n_2660),
.A2(n_475),
.B(n_474),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2410),
.B(n_2411),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2595),
.B(n_476),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2597),
.B(n_477),
.Y(n_3168)
);

NOR3xp33_ASAP7_75t_L g3169 ( 
.A(n_2755),
.B(n_478),
.C(n_477),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_SL g3170 ( 
.A(n_2648),
.B(n_478),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_L g3171 ( 
.A(n_2466),
.B(n_478),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2662),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2655),
.Y(n_3173)
);

AO21x1_ASAP7_75t_L g3174 ( 
.A1(n_2666),
.A2(n_480),
.B(n_479),
.Y(n_3174)
);

AOI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_2650),
.A2(n_482),
.B(n_481),
.Y(n_3175)
);

O2A1O1Ixp33_ASAP7_75t_L g3176 ( 
.A1(n_2766),
.A2(n_482),
.B(n_483),
.C(n_481),
.Y(n_3176)
);

BUFx2_ASAP7_75t_L g3177 ( 
.A(n_2772),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2606),
.Y(n_3178)
);

NOR2xp67_ASAP7_75t_SL g3179 ( 
.A(n_2396),
.B(n_481),
.Y(n_3179)
);

AOI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2633),
.A2(n_483),
.B(n_482),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_2544),
.B(n_484),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2802),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2523),
.A2(n_485),
.B(n_484),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2529),
.A2(n_486),
.B(n_485),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2685),
.B(n_486),
.Y(n_3185)
);

NOR2xp33_ASAP7_75t_L g3186 ( 
.A(n_2548),
.B(n_487),
.Y(n_3186)
);

O2A1O1Ixp33_ASAP7_75t_L g3187 ( 
.A1(n_2776),
.A2(n_488),
.B(n_489),
.C(n_487),
.Y(n_3187)
);

OAI321xp33_ASAP7_75t_L g3188 ( 
.A1(n_2822),
.A2(n_49),
.A3(n_51),
.B1(n_47),
.B2(n_48),
.C(n_50),
.Y(n_3188)
);

A2O1A1Ixp33_ASAP7_75t_L g3189 ( 
.A1(n_2827),
.A2(n_2695),
.B(n_2740),
.C(n_2687),
.Y(n_3189)
);

OAI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2616),
.A2(n_47),
.B(n_48),
.Y(n_3190)
);

INVx5_ASAP7_75t_L g3191 ( 
.A(n_2666),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_2522),
.B(n_488),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2609),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2549),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2587),
.B(n_488),
.Y(n_3195)
);

AOI21xp5_ASAP7_75t_L g3196 ( 
.A1(n_2530),
.A2(n_490),
.B(n_489),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2540),
.B(n_489),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2549),
.Y(n_3198)
);

OAI22xp5_ASAP7_75t_L g3199 ( 
.A1(n_2526),
.A2(n_492),
.B1(n_493),
.B2(n_491),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2697),
.B(n_491),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2471),
.B(n_493),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2816),
.B(n_494),
.Y(n_3202)
);

INVx3_ASAP7_75t_L g3203 ( 
.A(n_2769),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2602),
.B(n_495),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2629),
.B(n_495),
.Y(n_3205)
);

AOI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_2385),
.A2(n_497),
.B1(n_498),
.B2(n_496),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2769),
.Y(n_3207)
);

NOR3xp33_ASAP7_75t_L g3208 ( 
.A(n_2778),
.B(n_497),
.C(n_496),
.Y(n_3208)
);

OAI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_2620),
.A2(n_49),
.B(n_50),
.Y(n_3209)
);

O2A1O1Ixp5_ASAP7_75t_L g3210 ( 
.A1(n_2702),
.A2(n_499),
.B(n_500),
.C(n_498),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2627),
.B(n_499),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2641),
.Y(n_3212)
);

AND2x4_ASAP7_75t_L g3213 ( 
.A(n_2585),
.B(n_501),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2628),
.B(n_501),
.Y(n_3214)
);

AOI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2538),
.A2(n_503),
.B(n_502),
.Y(n_3215)
);

NOR2x1p5_ASAP7_75t_L g3216 ( 
.A(n_2705),
.B(n_502),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2592),
.B(n_502),
.Y(n_3217)
);

AOI21xp5_ASAP7_75t_L g3218 ( 
.A1(n_2539),
.A2(n_2495),
.B(n_2637),
.Y(n_3218)
);

AOI21xp33_ASAP7_75t_L g3219 ( 
.A1(n_2424),
.A2(n_504),
.B(n_503),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_2694),
.A2(n_507),
.B(n_504),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_2701),
.A2(n_508),
.B(n_507),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_2482),
.B(n_508),
.Y(n_3222)
);

O2A1O1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_2788),
.A2(n_509),
.B(n_510),
.C(n_508),
.Y(n_3223)
);

HB1xp67_ASAP7_75t_L g3224 ( 
.A(n_2590),
.Y(n_3224)
);

O2A1O1Ixp33_ASAP7_75t_L g3225 ( 
.A1(n_3189),
.A2(n_2805),
.B(n_2814),
.C(n_2806),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2851),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_3055),
.Y(n_3227)
);

OAI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_3137),
.A2(n_2790),
.B1(n_2593),
.B2(n_2621),
.Y(n_3228)
);

INVxp67_ASAP7_75t_SL g3229 ( 
.A(n_3092),
.Y(n_3229)
);

BUFx2_ASAP7_75t_R g3230 ( 
.A(n_3120),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3140),
.B(n_2598),
.Y(n_3231)
);

AND2x4_ASAP7_75t_L g3232 ( 
.A(n_3191),
.B(n_2589),
.Y(n_3232)
);

AOI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_2965),
.A2(n_2789),
.B1(n_2824),
.B2(n_2813),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2916),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_3066),
.A2(n_2669),
.B(n_2664),
.Y(n_3235)
);

BUFx6f_ASAP7_75t_L g3236 ( 
.A(n_3055),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3178),
.B(n_2577),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_3191),
.B(n_2491),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3193),
.B(n_2594),
.Y(n_3239)
);

INVxp33_ASAP7_75t_SL g3240 ( 
.A(n_2833),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3079),
.A2(n_2683),
.B(n_2670),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3083),
.A2(n_2686),
.B(n_2684),
.Y(n_3242)
);

BUFx6f_ASAP7_75t_L g3243 ( 
.A(n_3055),
.Y(n_3243)
);

AOI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_3051),
.A2(n_2564),
.B1(n_2409),
.B2(n_2533),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_SL g3245 ( 
.A(n_2915),
.B(n_2451),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_3084),
.A2(n_2386),
.B(n_2610),
.Y(n_3246)
);

A2O1A1Ixp33_ASAP7_75t_L g3247 ( 
.A1(n_2849),
.A2(n_3002),
.B(n_2966),
.C(n_2860),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3150),
.A2(n_2476),
.B(n_2451),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2879),
.A2(n_2476),
.B(n_2451),
.Y(n_3249)
);

OAI221xp5_ASAP7_75t_L g3250 ( 
.A1(n_2979),
.A2(n_2552),
.B1(n_2810),
.B2(n_2573),
.C(n_2524),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_SL g3251 ( 
.A(n_2872),
.B(n_2476),
.Y(n_3251)
);

BUFx6f_ASAP7_75t_L g3252 ( 
.A(n_2924),
.Y(n_3252)
);

INVx3_ASAP7_75t_L g3253 ( 
.A(n_3033),
.Y(n_3253)
);

BUFx6f_ASAP7_75t_L g3254 ( 
.A(n_3033),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_2882),
.B(n_2476),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_2835),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_SL g3257 ( 
.A(n_3191),
.B(n_2476),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_3147),
.B(n_2443),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_SL g3259 ( 
.A(n_3033),
.B(n_2494),
.Y(n_3259)
);

BUFx3_ASAP7_75t_L g3260 ( 
.A(n_2993),
.Y(n_3260)
);

AO21x2_ASAP7_75t_L g3261 ( 
.A1(n_2995),
.A2(n_2461),
.B(n_2419),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3212),
.B(n_2541),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2874),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_2884),
.A2(n_2494),
.B(n_2636),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_2892),
.A2(n_2494),
.B(n_2402),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2834),
.B(n_2543),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2844),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2880),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_2952),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2992),
.B(n_2532),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_2994),
.B(n_3001),
.Y(n_3271)
);

O2A1O1Ixp33_ASAP7_75t_L g3272 ( 
.A1(n_3071),
.A2(n_2558),
.B(n_2553),
.C(n_2490),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2846),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_2850),
.Y(n_3274)
);

BUFx3_ASAP7_75t_L g3275 ( 
.A(n_2862),
.Y(n_3275)
);

NOR3xp33_ASAP7_75t_L g3276 ( 
.A(n_3222),
.B(n_2463),
.C(n_2382),
.Y(n_3276)
);

NOR2x1_ASAP7_75t_L g3277 ( 
.A(n_3160),
.B(n_2649),
.Y(n_3277)
);

HB1xp67_ASAP7_75t_L g3278 ( 
.A(n_3016),
.Y(n_3278)
);

O2A1O1Ixp33_ASAP7_75t_L g3279 ( 
.A1(n_2875),
.A2(n_2639),
.B(n_2646),
.C(n_2453),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2865),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_SL g3281 ( 
.A(n_2911),
.B(n_2713),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_3218),
.A2(n_2736),
.B(n_2719),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2906),
.B(n_2718),
.Y(n_3283)
);

BUFx4f_ASAP7_75t_SL g3284 ( 
.A(n_2870),
.Y(n_3284)
);

INVxp67_ASAP7_75t_L g3285 ( 
.A(n_3046),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_3099),
.B(n_2765),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_3034),
.B(n_509),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2973),
.B(n_509),
.Y(n_3288)
);

AND2x4_ASAP7_75t_L g3289 ( 
.A(n_3203),
.B(n_3207),
.Y(n_3289)
);

OAI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_3124),
.A2(n_3160),
.B1(n_2949),
.B2(n_2830),
.Y(n_3290)
);

AOI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_2843),
.A2(n_511),
.B(n_510),
.Y(n_3291)
);

A2O1A1Ixp33_ASAP7_75t_L g3292 ( 
.A1(n_2890),
.A2(n_511),
.B(n_512),
.C(n_510),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3005),
.B(n_511),
.Y(n_3293)
);

BUFx6f_ASAP7_75t_L g3294 ( 
.A(n_3148),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3008),
.B(n_512),
.Y(n_3295)
);

AND2x6_ASAP7_75t_L g3296 ( 
.A(n_3203),
.B(n_3207),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_2852),
.A2(n_513),
.B(n_512),
.Y(n_3297)
);

AOI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_2857),
.A2(n_514),
.B(n_513),
.Y(n_3298)
);

CKINVDCx5p33_ASAP7_75t_R g3299 ( 
.A(n_3060),
.Y(n_3299)
);

INVxp67_ASAP7_75t_L g3300 ( 
.A(n_2910),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3012),
.B(n_514),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2891),
.A2(n_515),
.B(n_514),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_3100),
.B(n_515),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2893),
.Y(n_3304)
);

OR2x6_ASAP7_75t_L g3305 ( 
.A(n_2949),
.B(n_515),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3135),
.B(n_1080),
.Y(n_3306)
);

AOI22x1_ASAP7_75t_L g3307 ( 
.A1(n_3182),
.A2(n_517),
.B1(n_518),
.B2(n_516),
.Y(n_3307)
);

AO32x1_ASAP7_75t_L g3308 ( 
.A1(n_2941),
.A2(n_518),
.A3(n_519),
.B1(n_517),
.B2(n_516),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2894),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_2940),
.B(n_516),
.Y(n_3310)
);

AOI21xp5_ASAP7_75t_L g3311 ( 
.A1(n_2829),
.A2(n_518),
.B(n_517),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2831),
.A2(n_520),
.B(n_519),
.Y(n_3312)
);

OAI22xp5_ASAP7_75t_L g3313 ( 
.A1(n_2984),
.A2(n_520),
.B1(n_521),
.B2(n_519),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3042),
.A2(n_2904),
.B(n_3048),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_3148),
.Y(n_3315)
);

AOI21xp5_ASAP7_75t_L g3316 ( 
.A1(n_3095),
.A2(n_522),
.B(n_521),
.Y(n_3316)
);

OAI21xp33_ASAP7_75t_L g3317 ( 
.A1(n_2989),
.A2(n_52),
.B(n_53),
.Y(n_3317)
);

INVx2_ASAP7_75t_SL g3318 ( 
.A(n_3161),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2896),
.Y(n_3319)
);

O2A1O1Ixp33_ASAP7_75t_L g3320 ( 
.A1(n_2912),
.A2(n_524),
.B(n_525),
.C(n_523),
.Y(n_3320)
);

INVx3_ASAP7_75t_L g3321 ( 
.A(n_2961),
.Y(n_3321)
);

AOI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_3155),
.A2(n_524),
.B1(n_526),
.B2(n_523),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2928),
.Y(n_3323)
);

AOI22xp33_ASAP7_75t_L g3324 ( 
.A1(n_3105),
.A2(n_527),
.B1(n_528),
.B2(n_526),
.Y(n_3324)
);

OAI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_2853),
.A2(n_528),
.B1(n_529),
.B2(n_527),
.Y(n_3325)
);

INVx5_ASAP7_75t_L g3326 ( 
.A(n_2920),
.Y(n_3326)
);

BUFx12f_ASAP7_75t_L g3327 ( 
.A(n_2986),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2960),
.A2(n_528),
.B(n_527),
.Y(n_3328)
);

OR2x6_ASAP7_75t_SL g3329 ( 
.A(n_2905),
.B(n_1077),
.Y(n_3329)
);

BUFx2_ASAP7_75t_L g3330 ( 
.A(n_3148),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2933),
.B(n_529),
.Y(n_3331)
);

A2O1A1Ixp33_ASAP7_75t_L g3332 ( 
.A1(n_2958),
.A2(n_531),
.B(n_532),
.C(n_530),
.Y(n_3332)
);

CKINVDCx20_ASAP7_75t_R g3333 ( 
.A(n_3177),
.Y(n_3333)
);

AOI21x1_ASAP7_75t_L g3334 ( 
.A1(n_3041),
.A2(n_532),
.B(n_531),
.Y(n_3334)
);

INVx5_ASAP7_75t_L g3335 ( 
.A(n_2920),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_2978),
.B(n_1081),
.Y(n_3336)
);

AOI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_3053),
.A2(n_534),
.B1(n_535),
.B2(n_533),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_3006),
.B(n_533),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_3069),
.B(n_3122),
.Y(n_3339)
);

OAI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_2977),
.A2(n_536),
.B1(n_537),
.B2(n_534),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_2962),
.B(n_536),
.Y(n_3341)
);

AOI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3130),
.A2(n_3153),
.B1(n_2901),
.B2(n_2854),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3004),
.Y(n_3343)
);

AOI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_3076),
.A2(n_540),
.B(n_539),
.Y(n_3344)
);

BUFx3_ASAP7_75t_L g3345 ( 
.A(n_3020),
.Y(n_3345)
);

O2A1O1Ixp5_ASAP7_75t_L g3346 ( 
.A1(n_3080),
.A2(n_541),
.B(n_542),
.C(n_539),
.Y(n_3346)
);

AOI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_3103),
.A2(n_542),
.B(n_541),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_2969),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_2968),
.Y(n_3349)
);

OAI21x1_ASAP7_75t_L g3350 ( 
.A1(n_3025),
.A2(n_543),
.B(n_542),
.Y(n_3350)
);

O2A1O1Ixp33_ASAP7_75t_L g3351 ( 
.A1(n_2985),
.A2(n_544),
.B(n_545),
.C(n_543),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_2866),
.A2(n_546),
.B(n_545),
.Y(n_3352)
);

OR2x6_ASAP7_75t_L g3353 ( 
.A(n_3054),
.B(n_546),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3015),
.Y(n_3354)
);

AOI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_3125),
.A2(n_548),
.B(n_547),
.Y(n_3355)
);

HB1xp67_ASAP7_75t_L g3356 ( 
.A(n_3224),
.Y(n_3356)
);

OAI22x1_ASAP7_75t_L g3357 ( 
.A1(n_3216),
.A2(n_549),
.B1(n_550),
.B2(n_547),
.Y(n_3357)
);

BUFx3_ASAP7_75t_L g3358 ( 
.A(n_3049),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3032),
.B(n_551),
.Y(n_3359)
);

NOR2x1p5_ASAP7_75t_L g3360 ( 
.A(n_2961),
.B(n_551),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_2885),
.A2(n_3166),
.B(n_3172),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3029),
.B(n_552),
.Y(n_3362)
);

O2A1O1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_2887),
.A2(n_553),
.B(n_554),
.C(n_552),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2974),
.B(n_552),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_2971),
.B(n_554),
.Y(n_3365)
);

OAI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3018),
.A2(n_556),
.B1(n_557),
.B2(n_555),
.Y(n_3366)
);

INVx4_ASAP7_75t_L g3367 ( 
.A(n_2982),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_2867),
.B(n_558),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3192),
.B(n_558),
.Y(n_3369)
);

INVx3_ASAP7_75t_L g3370 ( 
.A(n_2982),
.Y(n_3370)
);

BUFx6f_ASAP7_75t_L g3371 ( 
.A(n_2953),
.Y(n_3371)
);

AOI22xp33_ASAP7_75t_L g3372 ( 
.A1(n_3105),
.A2(n_561),
.B1(n_562),
.B2(n_560),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3013),
.A2(n_561),
.B(n_560),
.Y(n_3373)
);

AND2x4_ASAP7_75t_L g3374 ( 
.A(n_2867),
.B(n_560),
.Y(n_3374)
);

O2A1O1Ixp33_ASAP7_75t_L g3375 ( 
.A1(n_3073),
.A2(n_564),
.B(n_565),
.C(n_563),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3039),
.A2(n_565),
.B1(n_566),
.B2(n_564),
.Y(n_3376)
);

BUFx2_ASAP7_75t_L g3377 ( 
.A(n_2873),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3195),
.B(n_568),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3105),
.A2(n_569),
.B1(n_570),
.B2(n_568),
.Y(n_3379)
);

NOR2x1_ASAP7_75t_L g3380 ( 
.A(n_2873),
.B(n_570),
.Y(n_3380)
);

INVxp67_ASAP7_75t_L g3381 ( 
.A(n_2836),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_2897),
.B(n_571),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_L g3383 ( 
.A(n_2948),
.B(n_572),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3105),
.A2(n_3052),
.B1(n_3123),
.B2(n_3017),
.Y(n_3384)
);

OAI21xp5_ASAP7_75t_L g3385 ( 
.A1(n_3158),
.A2(n_574),
.B(n_573),
.Y(n_3385)
);

A2O1A1Ixp33_ASAP7_75t_L g3386 ( 
.A1(n_2925),
.A2(n_3022),
.B(n_2914),
.C(n_2895),
.Y(n_3386)
);

INVx4_ASAP7_75t_L g3387 ( 
.A(n_2839),
.Y(n_3387)
);

OAI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_3211),
.A2(n_576),
.B1(n_577),
.B2(n_575),
.Y(n_3388)
);

AOI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_3106),
.A2(n_577),
.B(n_575),
.Y(n_3389)
);

OAI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3214),
.A2(n_578),
.B1(n_579),
.B2(n_577),
.Y(n_3390)
);

OAI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_2939),
.A2(n_2955),
.B1(n_3206),
.B2(n_2899),
.Y(n_3391)
);

O2A1O1Ixp33_ASAP7_75t_SL g3392 ( 
.A1(n_2921),
.A2(n_1079),
.B(n_1080),
.C(n_1078),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_L g3393 ( 
.A(n_3044),
.B(n_578),
.Y(n_3393)
);

CKINVDCx11_ASAP7_75t_R g3394 ( 
.A(n_3059),
.Y(n_3394)
);

OAI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_3204),
.A2(n_3205),
.B1(n_2935),
.B2(n_3010),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3107),
.Y(n_3396)
);

O2A1O1Ixp33_ASAP7_75t_L g3397 ( 
.A1(n_3197),
.A2(n_581),
.B(n_582),
.C(n_580),
.Y(n_3397)
);

AOI21xp5_ASAP7_75t_L g3398 ( 
.A1(n_3110),
.A2(n_583),
.B(n_582),
.Y(n_3398)
);

INVx8_ASAP7_75t_L g3399 ( 
.A(n_2839),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3171),
.B(n_583),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_2997),
.B(n_584),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3101),
.B(n_584),
.Y(n_3402)
);

BUFx3_ASAP7_75t_L g3403 ( 
.A(n_2967),
.Y(n_3403)
);

AO21x1_ASAP7_75t_L g3404 ( 
.A1(n_2957),
.A2(n_2889),
.B(n_2864),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_SL g3405 ( 
.A(n_2897),
.B(n_585),
.Y(n_3405)
);

BUFx8_ASAP7_75t_L g3406 ( 
.A(n_3056),
.Y(n_3406)
);

OAI22xp5_ASAP7_75t_L g3407 ( 
.A1(n_3038),
.A2(n_586),
.B1(n_587),
.B2(n_585),
.Y(n_3407)
);

A2O1A1Ixp33_ASAP7_75t_L g3408 ( 
.A1(n_2838),
.A2(n_589),
.B(n_590),
.C(n_588),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_3127),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2903),
.Y(n_3410)
);

INVx5_ASAP7_75t_L g3411 ( 
.A(n_2953),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_2868),
.A2(n_591),
.B(n_589),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2907),
.Y(n_3413)
);

OAI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3065),
.A2(n_592),
.B1(n_593),
.B2(n_591),
.Y(n_3414)
);

INVx4_ASAP7_75t_L g3415 ( 
.A(n_2861),
.Y(n_3415)
);

OAI22x1_ASAP7_75t_L g3416 ( 
.A1(n_2861),
.A2(n_592),
.B1(n_593),
.B2(n_591),
.Y(n_3416)
);

AND2x4_ASAP7_75t_L g3417 ( 
.A(n_2913),
.B(n_592),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2918),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_SL g3419 ( 
.A(n_2954),
.B(n_594),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_2856),
.B(n_595),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3024),
.B(n_596),
.Y(n_3421)
);

O2A1O1Ixp5_ASAP7_75t_L g3422 ( 
.A1(n_2964),
.A2(n_597),
.B(n_598),
.C(n_596),
.Y(n_3422)
);

NOR2xp33_ASAP7_75t_L g3423 ( 
.A(n_3179),
.B(n_596),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_2938),
.Y(n_3424)
);

NOR2xp33_ASAP7_75t_L g3425 ( 
.A(n_2959),
.B(n_2975),
.Y(n_3425)
);

AOI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_2858),
.A2(n_598),
.B(n_597),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2919),
.Y(n_3427)
);

O2A1O1Ixp33_ASAP7_75t_L g3428 ( 
.A1(n_3050),
.A2(n_598),
.B(n_599),
.C(n_597),
.Y(n_3428)
);

AOI21xp5_ASAP7_75t_L g3429 ( 
.A1(n_2944),
.A2(n_600),
.B(n_599),
.Y(n_3429)
);

A2O1A1Ixp33_ASAP7_75t_L g3430 ( 
.A1(n_3115),
.A2(n_600),
.B(n_601),
.C(n_599),
.Y(n_3430)
);

A2O1A1Ixp33_ASAP7_75t_L g3431 ( 
.A1(n_3128),
.A2(n_601),
.B(n_602),
.C(n_600),
.Y(n_3431)
);

O2A1O1Ixp5_ASAP7_75t_L g3432 ( 
.A1(n_3139),
.A2(n_602),
.B(n_603),
.C(n_601),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_SL g3433 ( 
.A(n_2954),
.B(n_603),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_3167),
.B(n_604),
.Y(n_3434)
);

O2A1O1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_3142),
.A2(n_3027),
.B(n_2942),
.C(n_2946),
.Y(n_3435)
);

A2O1A1Ixp33_ASAP7_75t_L g3436 ( 
.A1(n_3023),
.A2(n_606),
.B(n_607),
.C(n_604),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3168),
.B(n_3145),
.Y(n_3437)
);

OAI21xp33_ASAP7_75t_SL g3438 ( 
.A1(n_3011),
.A2(n_608),
.B(n_606),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2837),
.B(n_608),
.Y(n_3439)
);

O2A1O1Ixp33_ASAP7_75t_L g3440 ( 
.A1(n_2981),
.A2(n_610),
.B(n_611),
.C(n_609),
.Y(n_3440)
);

AOI21xp5_ASAP7_75t_L g3441 ( 
.A1(n_2987),
.A2(n_610),
.B(n_609),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3081),
.B(n_611),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_2988),
.A2(n_612),
.B(n_611),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3201),
.B(n_612),
.Y(n_3444)
);

AOI221x1_ASAP7_75t_L g3445 ( 
.A1(n_3094),
.A2(n_614),
.B1(n_615),
.B2(n_613),
.C(n_612),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3082),
.B(n_613),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_2922),
.Y(n_3447)
);

AOI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3169),
.A2(n_614),
.B1(n_615),
.B2(n_613),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3058),
.B(n_614),
.Y(n_3449)
);

A2O1A1Ixp33_ASAP7_75t_L g3450 ( 
.A1(n_3026),
.A2(n_617),
.B(n_618),
.C(n_616),
.Y(n_3450)
);

OAI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_2976),
.A2(n_617),
.B1(n_619),
.B2(n_616),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3217),
.B(n_617),
.Y(n_3452)
);

NOR2xp33_ASAP7_75t_L g3453 ( 
.A(n_2998),
.B(n_620),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3019),
.Y(n_3454)
);

AOI21xp5_ASAP7_75t_L g3455 ( 
.A1(n_3064),
.A2(n_622),
.B(n_621),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3146),
.B(n_621),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3030),
.A2(n_3213),
.B1(n_3047),
.B2(n_3085),
.Y(n_3457)
);

A2O1A1Ixp33_ASAP7_75t_SL g3458 ( 
.A1(n_3072),
.A2(n_55),
.B(n_52),
.C(n_54),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_2926),
.Y(n_3459)
);

OAI21x1_ASAP7_75t_L g3460 ( 
.A1(n_3007),
.A2(n_623),
.B(n_622),
.Y(n_3460)
);

OAI21x1_ASAP7_75t_SL g3461 ( 
.A1(n_3174),
.A2(n_624),
.B(n_623),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_3070),
.B(n_624),
.Y(n_3462)
);

OAI22xp5_ASAP7_75t_L g3463 ( 
.A1(n_3213),
.A2(n_626),
.B1(n_627),
.B2(n_625),
.Y(n_3463)
);

CKINVDCx5p33_ASAP7_75t_R g3464 ( 
.A(n_3202),
.Y(n_3464)
);

BUFx6f_ASAP7_75t_L g3465 ( 
.A(n_2953),
.Y(n_3465)
);

NOR2xp67_ASAP7_75t_L g3466 ( 
.A(n_2917),
.B(n_626),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_R g3467 ( 
.A(n_3074),
.B(n_627),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_2980),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_SL g3469 ( 
.A(n_2980),
.B(n_629),
.Y(n_3469)
);

O2A1O1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_3219),
.A2(n_630),
.B(n_631),
.C(n_629),
.Y(n_3470)
);

BUFx3_ASAP7_75t_L g3471 ( 
.A(n_3141),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_2983),
.Y(n_3472)
);

AO21x1_ASAP7_75t_L g3473 ( 
.A1(n_2900),
.A2(n_632),
.B(n_631),
.Y(n_3473)
);

CKINVDCx20_ASAP7_75t_R g3474 ( 
.A(n_3152),
.Y(n_3474)
);

AOI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3156),
.A2(n_633),
.B(n_632),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_2983),
.Y(n_3476)
);

AOI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_3162),
.A2(n_634),
.B(n_633),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_2929),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_2930),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_2983),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2931),
.Y(n_3481)
);

BUFx6f_ASAP7_75t_L g3482 ( 
.A(n_3078),
.Y(n_3482)
);

AOI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_3208),
.A2(n_634),
.B1(n_635),
.B2(n_633),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3087),
.B(n_634),
.Y(n_3484)
);

OAI21x1_ASAP7_75t_L g3485 ( 
.A1(n_3043),
.A2(n_636),
.B(n_635),
.Y(n_3485)
);

BUFx6f_ASAP7_75t_L g3486 ( 
.A(n_3078),
.Y(n_3486)
);

NOR2xp33_ASAP7_75t_L g3487 ( 
.A(n_3021),
.B(n_636),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3129),
.A2(n_638),
.B1(n_639),
.B2(n_637),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3138),
.B(n_2932),
.Y(n_3489)
);

AOI22xp33_ASAP7_75t_L g3490 ( 
.A1(n_3149),
.A2(n_3075),
.B1(n_3088),
.B2(n_3108),
.Y(n_3490)
);

O2A1O1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_3199),
.A2(n_639),
.B(n_640),
.C(n_638),
.Y(n_3491)
);

BUFx6f_ASAP7_75t_L g3492 ( 
.A(n_3078),
.Y(n_3492)
);

CKINVDCx8_ASAP7_75t_R g3493 ( 
.A(n_3091),
.Y(n_3493)
);

AOI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3063),
.A2(n_640),
.B(n_639),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_L g3495 ( 
.A(n_3045),
.B(n_640),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_2934),
.B(n_641),
.Y(n_3496)
);

INVx3_ASAP7_75t_L g3497 ( 
.A(n_3091),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_2937),
.B(n_641),
.Y(n_3498)
);

AO32x1_ASAP7_75t_L g3499 ( 
.A1(n_3111),
.A2(n_643),
.A3(n_644),
.B1(n_642),
.B2(n_641),
.Y(n_3499)
);

NOR2xp33_ASAP7_75t_L g3500 ( 
.A(n_3181),
.B(n_642),
.Y(n_3500)
);

NOR2xp33_ASAP7_75t_L g3501 ( 
.A(n_3186),
.B(n_642),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_2943),
.B(n_643),
.Y(n_3502)
);

BUFx3_ASAP7_75t_L g3503 ( 
.A(n_3086),
.Y(n_3503)
);

AOI22xp5_ASAP7_75t_L g3504 ( 
.A1(n_3109),
.A2(n_646),
.B1(n_647),
.B2(n_645),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3194),
.A2(n_646),
.B(n_645),
.Y(n_3505)
);

O2A1O1Ixp33_ASAP7_75t_L g3506 ( 
.A1(n_3061),
.A2(n_646),
.B(n_647),
.C(n_645),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3126),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3113),
.B(n_648),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3198),
.A2(n_649),
.B(n_648),
.Y(n_3509)
);

AND2x4_ASAP7_75t_L g3510 ( 
.A(n_3116),
.B(n_648),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_L g3511 ( 
.A1(n_3114),
.A2(n_650),
.B1(n_651),
.B2(n_649),
.Y(n_3511)
);

O2A1O1Ixp33_ASAP7_75t_L g3512 ( 
.A1(n_3151),
.A2(n_3121),
.B(n_3035),
.C(n_3036),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_SL g3513 ( 
.A(n_3040),
.B(n_649),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_2972),
.A2(n_653),
.B(n_651),
.Y(n_3514)
);

OAI22x1_ASAP7_75t_L g3515 ( 
.A1(n_2881),
.A2(n_653),
.B1(n_654),
.B2(n_651),
.Y(n_3515)
);

CKINVDCx5p33_ASAP7_75t_R g3516 ( 
.A(n_2902),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_2840),
.B(n_1072),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_2999),
.A2(n_654),
.B(n_653),
.Y(n_3518)
);

O2A1O1Ixp33_ASAP7_75t_L g3519 ( 
.A1(n_3097),
.A2(n_655),
.B(n_656),
.C(n_654),
.Y(n_3519)
);

BUFx2_ASAP7_75t_L g3520 ( 
.A(n_3116),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3133),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_SL g3522 ( 
.A(n_3131),
.B(n_3165),
.Y(n_3522)
);

OAI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_3210),
.A2(n_656),
.B(n_655),
.Y(n_3523)
);

OAI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3190),
.A2(n_657),
.B1(n_658),
.B2(n_655),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_2842),
.B(n_657),
.Y(n_3525)
);

BUFx2_ASAP7_75t_L g3526 ( 
.A(n_3131),
.Y(n_3526)
);

CKINVDCx5p33_ASAP7_75t_R g3527 ( 
.A(n_2927),
.Y(n_3527)
);

INVxp67_ASAP7_75t_SL g3528 ( 
.A(n_2859),
.Y(n_3528)
);

O2A1O1Ixp5_ASAP7_75t_L g3529 ( 
.A1(n_2996),
.A2(n_659),
.B(n_660),
.C(n_658),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_2863),
.B(n_658),
.Y(n_3530)
);

OAI21xp33_ASAP7_75t_L g3531 ( 
.A1(n_3209),
.A2(n_54),
.B(n_55),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_3000),
.A2(n_661),
.B(n_660),
.Y(n_3532)
);

OAI22xp5_ASAP7_75t_L g3533 ( 
.A1(n_3136),
.A2(n_662),
.B1(n_663),
.B2(n_661),
.Y(n_3533)
);

OAI22xp5_ASAP7_75t_L g3534 ( 
.A1(n_3144),
.A2(n_663),
.B1(n_664),
.B2(n_662),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3132),
.B(n_663),
.Y(n_3535)
);

NAND3xp33_ASAP7_75t_SL g3536 ( 
.A(n_3104),
.B(n_3187),
.C(n_3176),
.Y(n_3536)
);

O2A1O1Ixp33_ASAP7_75t_L g3537 ( 
.A1(n_3223),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3134),
.A2(n_667),
.B1(n_668),
.B2(n_666),
.Y(n_3538)
);

INVx1_ASAP7_75t_SL g3539 ( 
.A(n_3112),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_2883),
.B(n_1070),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3003),
.A2(n_667),
.B(n_666),
.Y(n_3541)
);

NOR2xp67_ASAP7_75t_L g3542 ( 
.A(n_3188),
.B(n_668),
.Y(n_3542)
);

OAI21x1_ASAP7_75t_L g3543 ( 
.A1(n_3173),
.A2(n_3102),
.B(n_3068),
.Y(n_3543)
);

A2O1A1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_2945),
.A2(n_670),
.B(n_671),
.C(n_669),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_2886),
.B(n_669),
.Y(n_3545)
);

AOI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_2869),
.A2(n_672),
.B(n_670),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_2871),
.A2(n_673),
.B(n_672),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_2990),
.B(n_673),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_2876),
.A2(n_674),
.B(n_673),
.Y(n_3549)
);

AOI22xp33_ASAP7_75t_L g3550 ( 
.A1(n_3031),
.A2(n_3154),
.B1(n_2888),
.B2(n_2951),
.Y(n_3550)
);

OAI21xp33_ASAP7_75t_SL g3551 ( 
.A1(n_3170),
.A2(n_675),
.B(n_674),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_2950),
.Y(n_3552)
);

AOI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_2877),
.A2(n_676),
.B(n_675),
.Y(n_3553)
);

AOI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_2878),
.A2(n_677),
.B(n_676),
.Y(n_3554)
);

A2O1A1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_2947),
.A2(n_677),
.B(n_678),
.C(n_676),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3157),
.B(n_1089),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3159),
.B(n_679),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_2923),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_SL g3559 ( 
.A(n_2936),
.B(n_679),
.Y(n_3559)
);

O2A1O1Ixp33_ASAP7_75t_L g3560 ( 
.A1(n_3014),
.A2(n_682),
.B(n_683),
.C(n_681),
.Y(n_3560)
);

AO21x1_ASAP7_75t_L g3561 ( 
.A1(n_2832),
.A2(n_682),
.B(n_681),
.Y(n_3561)
);

OR2x2_ASAP7_75t_L g3562 ( 
.A(n_3057),
.B(n_683),
.Y(n_3562)
);

BUFx6f_ASAP7_75t_L g3563 ( 
.A(n_3200),
.Y(n_3563)
);

AOI21xp33_ASAP7_75t_L g3564 ( 
.A1(n_3185),
.A2(n_687),
.B(n_686),
.Y(n_3564)
);

NOR3xp33_ASAP7_75t_SL g3565 ( 
.A(n_3143),
.B(n_1075),
.C(n_1074),
.Y(n_3565)
);

AOI22xp5_ASAP7_75t_L g3566 ( 
.A1(n_3062),
.A2(n_687),
.B1(n_688),
.B2(n_686),
.Y(n_3566)
);

O2A1O1Ixp5_ASAP7_75t_SL g3567 ( 
.A1(n_3037),
.A2(n_687),
.B(n_688),
.C(n_686),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3067),
.B(n_688),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_2991),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_SL g3570 ( 
.A(n_3180),
.B(n_689),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3077),
.B(n_689),
.Y(n_3571)
);

O2A1O1Ixp33_ASAP7_75t_L g3572 ( 
.A1(n_3089),
.A2(n_691),
.B(n_692),
.C(n_690),
.Y(n_3572)
);

AND2x2_ASAP7_75t_SL g3573 ( 
.A(n_3163),
.B(n_690),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3090),
.B(n_690),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3093),
.Y(n_3575)
);

A2O1A1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_3096),
.A2(n_694),
.B(n_695),
.C(n_693),
.Y(n_3576)
);

OAI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_3009),
.A2(n_694),
.B1(n_695),
.B2(n_693),
.Y(n_3577)
);

AOI21xp5_ASAP7_75t_L g3578 ( 
.A1(n_3098),
.A2(n_696),
.B(n_695),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_3117),
.B(n_696),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3118),
.B(n_697),
.Y(n_3580)
);

AND2x4_ASAP7_75t_L g3581 ( 
.A(n_3119),
.B(n_697),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3028),
.B(n_698),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3183),
.B(n_699),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_SL g3584 ( 
.A(n_2841),
.B(n_699),
.Y(n_3584)
);

CKINVDCx5p33_ASAP7_75t_R g3585 ( 
.A(n_3184),
.Y(n_3585)
);

OAI22xp5_ASAP7_75t_L g3586 ( 
.A1(n_3196),
.A2(n_700),
.B1(n_701),
.B2(n_699),
.Y(n_3586)
);

INVx3_ASAP7_75t_L g3587 ( 
.A(n_3175),
.Y(n_3587)
);

AOI22xp33_ASAP7_75t_L g3588 ( 
.A1(n_3215),
.A2(n_702),
.B1(n_703),
.B2(n_700),
.Y(n_3588)
);

BUFx6f_ASAP7_75t_L g3589 ( 
.A(n_3221),
.Y(n_3589)
);

AOI22xp33_ASAP7_75t_L g3590 ( 
.A1(n_2898),
.A2(n_703),
.B1(n_704),
.B2(n_702),
.Y(n_3590)
);

AOI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_2845),
.A2(n_705),
.B(n_704),
.Y(n_3591)
);

A2O1A1Ixp33_ASAP7_75t_L g3592 ( 
.A1(n_2908),
.A2(n_705),
.B(n_706),
.C(n_704),
.Y(n_3592)
);

O2A1O1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_3164),
.A2(n_706),
.B(n_707),
.C(n_705),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_2909),
.B(n_707),
.Y(n_3594)
);

OAI21x1_ASAP7_75t_L g3595 ( 
.A1(n_2847),
.A2(n_710),
.B(n_709),
.Y(n_3595)
);

NOR2xp67_ASAP7_75t_L g3596 ( 
.A(n_3220),
.B(n_709),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_2848),
.A2(n_710),
.B(n_709),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2956),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_2963),
.Y(n_3599)
);

O2A1O1Ixp33_ASAP7_75t_L g3600 ( 
.A1(n_2970),
.A2(n_711),
.B(n_712),
.C(n_710),
.Y(n_3600)
);

INVx4_ASAP7_75t_L g3601 ( 
.A(n_2855),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3140),
.B(n_713),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_3247),
.A2(n_716),
.B(n_714),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3252),
.B(n_716),
.Y(n_3604)
);

OAI21x1_ASAP7_75t_L g3605 ( 
.A1(n_3248),
.A2(n_718),
.B(n_717),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3336),
.B(n_3306),
.Y(n_3606)
);

INVx2_ASAP7_75t_SL g3607 ( 
.A(n_3406),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3234),
.B(n_717),
.Y(n_3608)
);

AOI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_3339),
.A2(n_1079),
.B1(n_1082),
.B2(n_1078),
.Y(n_3609)
);

AND2x4_ASAP7_75t_L g3610 ( 
.A(n_3387),
.B(n_718),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_SL g3611 ( 
.A1(n_3305),
.A2(n_720),
.B(n_719),
.Y(n_3611)
);

AND2x4_ASAP7_75t_L g3612 ( 
.A(n_3387),
.B(n_719),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3252),
.B(n_719),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3226),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3314),
.A2(n_721),
.B(n_720),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_L g3616 ( 
.A1(n_3249),
.A2(n_722),
.B(n_721),
.Y(n_3616)
);

AO31x2_ASAP7_75t_L g3617 ( 
.A1(n_3454),
.A2(n_723),
.A3(n_724),
.B(n_722),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3271),
.B(n_725),
.Y(n_3618)
);

OAI21x1_ASAP7_75t_L g3619 ( 
.A1(n_3507),
.A2(n_3521),
.B(n_3282),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3231),
.B(n_726),
.Y(n_3620)
);

AO31x2_ASAP7_75t_L g3621 ( 
.A1(n_3601),
.A2(n_727),
.A3(n_728),
.B(n_726),
.Y(n_3621)
);

AOI221xp5_ASAP7_75t_SL g3622 ( 
.A1(n_3357),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_3622)
);

NAND3xp33_ASAP7_75t_L g3623 ( 
.A(n_3328),
.B(n_731),
.C(n_730),
.Y(n_3623)
);

OAI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3422),
.A2(n_733),
.B(n_732),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3263),
.B(n_3268),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3361),
.A2(n_734),
.B(n_733),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_SL g3627 ( 
.A(n_3230),
.B(n_3240),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_SL g3628 ( 
.A(n_3415),
.B(n_736),
.Y(n_3628)
);

A2O1A1Ixp33_ASAP7_75t_L g3629 ( 
.A1(n_3466),
.A2(n_737),
.B(n_738),
.C(n_736),
.Y(n_3629)
);

INVx2_ASAP7_75t_SL g3630 ( 
.A(n_3406),
.Y(n_3630)
);

AO31x2_ASAP7_75t_L g3631 ( 
.A1(n_3601),
.A2(n_738),
.A3(n_739),
.B(n_737),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_L g3632 ( 
.A(n_3258),
.B(n_740),
.Y(n_3632)
);

AOI21xp33_ASAP7_75t_L g3633 ( 
.A1(n_3435),
.A2(n_742),
.B(n_741),
.Y(n_3633)
);

OA21x2_ASAP7_75t_L g3634 ( 
.A1(n_3522),
.A2(n_742),
.B(n_741),
.Y(n_3634)
);

OAI21x1_ASAP7_75t_L g3635 ( 
.A1(n_3264),
.A2(n_744),
.B(n_743),
.Y(n_3635)
);

AO31x2_ASAP7_75t_L g3636 ( 
.A1(n_3473),
.A2(n_744),
.A3(n_745),
.B(n_743),
.Y(n_3636)
);

OAI21x1_ASAP7_75t_L g3637 ( 
.A1(n_3543),
.A2(n_744),
.B(n_743),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_3318),
.B(n_745),
.Y(n_3638)
);

NOR4xp25_ASAP7_75t_L g3639 ( 
.A(n_3228),
.B(n_747),
.C(n_748),
.D(n_746),
.Y(n_3639)
);

AO21x1_ASAP7_75t_L g3640 ( 
.A1(n_3290),
.A2(n_748),
.B(n_747),
.Y(n_3640)
);

NOR4xp25_ASAP7_75t_L g3641 ( 
.A(n_3317),
.B(n_750),
.C(n_751),
.D(n_749),
.Y(n_3641)
);

AOI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_3457),
.A2(n_751),
.B(n_750),
.Y(n_3642)
);

OAI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_3305),
.A2(n_751),
.B1(n_752),
.B2(n_750),
.Y(n_3643)
);

AOI221xp5_ASAP7_75t_SL g3644 ( 
.A1(n_3250),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3323),
.Y(n_3645)
);

AOI21x1_ASAP7_75t_L g3646 ( 
.A1(n_3334),
.A2(n_753),
.B(n_752),
.Y(n_3646)
);

OAI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_3329),
.A2(n_755),
.B1(n_756),
.B2(n_754),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3396),
.Y(n_3648)
);

INVx3_ASAP7_75t_SL g3649 ( 
.A(n_3299),
.Y(n_3649)
);

OA21x2_ASAP7_75t_L g3650 ( 
.A1(n_3460),
.A2(n_759),
.B(n_758),
.Y(n_3650)
);

HB1xp67_ASAP7_75t_L g3651 ( 
.A(n_3356),
.Y(n_3651)
);

INVx3_ASAP7_75t_L g3652 ( 
.A(n_3367),
.Y(n_3652)
);

AOI21x1_ASAP7_75t_L g3653 ( 
.A1(n_3259),
.A2(n_759),
.B(n_758),
.Y(n_3653)
);

AOI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_3235),
.A2(n_760),
.B(n_759),
.Y(n_3654)
);

NAND2x1p5_ASAP7_75t_L g3655 ( 
.A(n_3275),
.B(n_3367),
.Y(n_3655)
);

OAI21x1_ASAP7_75t_L g3656 ( 
.A1(n_3587),
.A2(n_3265),
.B(n_3245),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_3467),
.B(n_761),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3241),
.A2(n_764),
.B(n_763),
.Y(n_3658)
);

AOI21x1_ASAP7_75t_SL g3659 ( 
.A1(n_3420),
.A2(n_766),
.B(n_765),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3348),
.B(n_3349),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3242),
.A2(n_768),
.B(n_767),
.Y(n_3661)
);

OAI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3346),
.A2(n_768),
.B(n_767),
.Y(n_3662)
);

INVx2_ASAP7_75t_SL g3663 ( 
.A(n_3345),
.Y(n_3663)
);

INVx4_ASAP7_75t_L g3664 ( 
.A(n_3284),
.Y(n_3664)
);

AO32x2_ASAP7_75t_L g3665 ( 
.A1(n_3395),
.A2(n_784),
.A3(n_792),
.B1(n_778),
.B2(n_771),
.Y(n_3665)
);

A2O1A1Ixp33_ASAP7_75t_L g3666 ( 
.A1(n_3531),
.A2(n_771),
.B(n_772),
.C(n_770),
.Y(n_3666)
);

AOI22xp5_ASAP7_75t_L g3667 ( 
.A1(n_3516),
.A2(n_1072),
.B1(n_1073),
.B2(n_1071),
.Y(n_3667)
);

NOR2xp33_ASAP7_75t_L g3668 ( 
.A(n_3300),
.B(n_772),
.Y(n_3668)
);

INVx1_ASAP7_75t_SL g3669 ( 
.A(n_3394),
.Y(n_3669)
);

BUFx2_ASAP7_75t_L g3670 ( 
.A(n_3474),
.Y(n_3670)
);

AOI221x1_ASAP7_75t_L g3671 ( 
.A1(n_3416),
.A2(n_775),
.B1(n_776),
.B2(n_774),
.C(n_773),
.Y(n_3671)
);

AND2x6_ASAP7_75t_L g3672 ( 
.A(n_3471),
.B(n_775),
.Y(n_3672)
);

OAI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3529),
.A2(n_778),
.B(n_777),
.Y(n_3673)
);

NAND3xp33_ASAP7_75t_L g3674 ( 
.A(n_3423),
.B(n_778),
.C(n_777),
.Y(n_3674)
);

OAI21x1_ASAP7_75t_L g3675 ( 
.A1(n_3598),
.A2(n_3599),
.B(n_3497),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3286),
.B(n_779),
.Y(n_3676)
);

A2O1A1Ixp33_ASAP7_75t_L g3677 ( 
.A1(n_3506),
.A2(n_780),
.B(n_781),
.C(n_779),
.Y(n_3677)
);

CKINVDCx20_ASAP7_75t_R g3678 ( 
.A(n_3333),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3310),
.B(n_3381),
.Y(n_3679)
);

BUFx6f_ASAP7_75t_L g3680 ( 
.A(n_3358),
.Y(n_3680)
);

INVx4_ASAP7_75t_L g3681 ( 
.A(n_3399),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3558),
.A2(n_785),
.B(n_783),
.Y(n_3682)
);

AOI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3575),
.A2(n_785),
.B(n_783),
.Y(n_3683)
);

OAI21x1_ASAP7_75t_L g3684 ( 
.A1(n_3253),
.A2(n_785),
.B(n_783),
.Y(n_3684)
);

OAI21xp5_ASAP7_75t_L g3685 ( 
.A1(n_3432),
.A2(n_787),
.B(n_786),
.Y(n_3685)
);

AOI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3377),
.A2(n_787),
.B(n_786),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_3283),
.B(n_788),
.Y(n_3687)
);

AOI21x1_ASAP7_75t_L g3688 ( 
.A1(n_3251),
.A2(n_790),
.B(n_789),
.Y(n_3688)
);

OA21x2_ASAP7_75t_L g3689 ( 
.A1(n_3485),
.A2(n_790),
.B(n_789),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3256),
.Y(n_3690)
);

OAI21x1_ASAP7_75t_L g3691 ( 
.A1(n_3253),
.A2(n_791),
.B(n_790),
.Y(n_3691)
);

OAI21x1_ASAP7_75t_L g3692 ( 
.A1(n_3255),
.A2(n_3257),
.B(n_3468),
.Y(n_3692)
);

OAI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3476),
.A2(n_792),
.B(n_791),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_SL g3694 ( 
.A1(n_3360),
.A2(n_794),
.B(n_793),
.Y(n_3694)
);

AND2x4_ASAP7_75t_L g3695 ( 
.A(n_3326),
.B(n_794),
.Y(n_3695)
);

CKINVDCx11_ASAP7_75t_R g3696 ( 
.A(n_3327),
.Y(n_3696)
);

OAI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3480),
.A2(n_796),
.B(n_795),
.Y(n_3697)
);

OAI21xp5_ASAP7_75t_SL g3698 ( 
.A1(n_3277),
.A2(n_1066),
.B(n_1065),
.Y(n_3698)
);

BUFx2_ASAP7_75t_L g3699 ( 
.A(n_3399),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3410),
.B(n_796),
.Y(n_3700)
);

OAI21x1_ASAP7_75t_L g3701 ( 
.A1(n_3246),
.A2(n_798),
.B(n_797),
.Y(n_3701)
);

OAI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3342),
.A2(n_798),
.B(n_797),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_3326),
.B(n_799),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3343),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3354),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3267),
.Y(n_3706)
);

A2O1A1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_3363),
.A2(n_800),
.B(n_801),
.C(n_799),
.Y(n_3707)
);

OAI21x1_ASAP7_75t_L g3708 ( 
.A1(n_3350),
.A2(n_801),
.B(n_800),
.Y(n_3708)
);

BUFx8_ASAP7_75t_L g3709 ( 
.A(n_3260),
.Y(n_3709)
);

AO32x2_ASAP7_75t_L g3710 ( 
.A1(n_3463),
.A2(n_817),
.A3(n_824),
.B1(n_809),
.B2(n_802),
.Y(n_3710)
);

OA21x2_ASAP7_75t_L g3711 ( 
.A1(n_3445),
.A2(n_3569),
.B(n_3513),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3413),
.B(n_801),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3418),
.B(n_802),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3427),
.B(n_802),
.Y(n_3714)
);

NAND2x1_ASAP7_75t_L g3715 ( 
.A(n_3296),
.B(n_804),
.Y(n_3715)
);

NOR2xp67_ASAP7_75t_L g3716 ( 
.A(n_3269),
.B(n_806),
.Y(n_3716)
);

BUFx2_ASAP7_75t_L g3717 ( 
.A(n_3330),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3527),
.A2(n_808),
.B1(n_809),
.B2(n_807),
.Y(n_3718)
);

AO31x2_ASAP7_75t_L g3719 ( 
.A1(n_3404),
.A2(n_810),
.A3(n_811),
.B(n_807),
.Y(n_3719)
);

A2O1A1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_3428),
.A2(n_811),
.B(n_812),
.C(n_810),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3447),
.B(n_813),
.Y(n_3721)
);

OA21x2_ASAP7_75t_L g3722 ( 
.A1(n_3386),
.A2(n_815),
.B(n_814),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_SL g3723 ( 
.A(n_3326),
.B(n_814),
.Y(n_3723)
);

NOR2xp67_ASAP7_75t_L g3724 ( 
.A(n_3269),
.B(n_817),
.Y(n_3724)
);

OAI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3225),
.A2(n_817),
.B(n_816),
.Y(n_3725)
);

AO31x2_ASAP7_75t_L g3726 ( 
.A1(n_3561),
.A2(n_819),
.A3(n_820),
.B(n_818),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3459),
.B(n_819),
.Y(n_3727)
);

AO31x2_ASAP7_75t_L g3728 ( 
.A1(n_3391),
.A2(n_820),
.A3(n_821),
.B(n_819),
.Y(n_3728)
);

OAI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3408),
.A2(n_822),
.B(n_821),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3273),
.Y(n_3730)
);

OAI21x1_ASAP7_75t_L g3731 ( 
.A1(n_3595),
.A2(n_823),
.B(n_822),
.Y(n_3731)
);

AO21x2_ASAP7_75t_L g3732 ( 
.A1(n_3461),
.A2(n_824),
.B(n_822),
.Y(n_3732)
);

OAI21x1_ASAP7_75t_L g3733 ( 
.A1(n_3567),
.A2(n_3385),
.B(n_3523),
.Y(n_3733)
);

AND2x2_ASAP7_75t_SL g3734 ( 
.A(n_3374),
.B(n_826),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3274),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3478),
.B(n_827),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3479),
.B(n_827),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3481),
.B(n_827),
.Y(n_3738)
);

OAI21x1_ASAP7_75t_L g3739 ( 
.A1(n_3550),
.A2(n_3307),
.B(n_3352),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3280),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3584),
.A2(n_829),
.B(n_828),
.Y(n_3741)
);

AND2x4_ASAP7_75t_L g3742 ( 
.A(n_3335),
.B(n_830),
.Y(n_3742)
);

NOR2xp67_ASAP7_75t_SL g3743 ( 
.A(n_3254),
.B(n_831),
.Y(n_3743)
);

OAI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3412),
.A2(n_835),
.B(n_834),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3304),
.A2(n_3319),
.B(n_3309),
.Y(n_3745)
);

AOI221xp5_ASAP7_75t_L g3746 ( 
.A1(n_3338),
.A2(n_838),
.B1(n_840),
.B2(n_837),
.C(n_836),
.Y(n_3746)
);

AOI21xp5_ASAP7_75t_L g3747 ( 
.A1(n_3528),
.A2(n_838),
.B(n_837),
.Y(n_3747)
);

CKINVDCx14_ASAP7_75t_R g3748 ( 
.A(n_3353),
.Y(n_3748)
);

A2O1A1Ixp33_ASAP7_75t_L g3749 ( 
.A1(n_3560),
.A2(n_842),
.B(n_843),
.C(n_840),
.Y(n_3749)
);

OAI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3519),
.A2(n_844),
.B(n_842),
.Y(n_3750)
);

OAI21x1_ASAP7_75t_L g3751 ( 
.A1(n_3424),
.A2(n_845),
.B(n_844),
.Y(n_3751)
);

OAI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3537),
.A2(n_846),
.B(n_845),
.Y(n_3752)
);

AOI21xp5_ASAP7_75t_L g3753 ( 
.A1(n_3512),
.A2(n_847),
.B(n_846),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3237),
.Y(n_3754)
);

BUFx6f_ASAP7_75t_L g3755 ( 
.A(n_3238),
.Y(n_3755)
);

INVx1_ASAP7_75t_SL g3756 ( 
.A(n_3403),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3591),
.A2(n_848),
.B(n_847),
.Y(n_3757)
);

OAI21x1_ASAP7_75t_L g3758 ( 
.A1(n_3597),
.A2(n_849),
.B(n_848),
.Y(n_3758)
);

OR2x2_ASAP7_75t_L g3759 ( 
.A(n_3278),
.B(n_849),
.Y(n_3759)
);

BUFx6f_ASAP7_75t_L g3760 ( 
.A(n_3238),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3270),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_3437),
.A2(n_3489),
.B(n_3458),
.Y(n_3762)
);

AOI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3520),
.A2(n_850),
.B(n_849),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3239),
.Y(n_3764)
);

NAND2x1_ASAP7_75t_L g3765 ( 
.A(n_3296),
.B(n_851),
.Y(n_3765)
);

OAI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3384),
.A2(n_853),
.B1(n_854),
.B2(n_852),
.Y(n_3766)
);

OAI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3292),
.A2(n_3233),
.B(n_3596),
.Y(n_3767)
);

OAI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_3572),
.A2(n_854),
.B(n_853),
.Y(n_3768)
);

OAI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3380),
.A2(n_855),
.B(n_854),
.Y(n_3769)
);

AO31x2_ASAP7_75t_L g3770 ( 
.A1(n_3325),
.A2(n_856),
.A3(n_857),
.B(n_855),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_3536),
.A2(n_858),
.B(n_857),
.Y(n_3771)
);

O2A1O1Ixp5_ASAP7_75t_L g3772 ( 
.A1(n_3579),
.A2(n_858),
.B(n_859),
.C(n_857),
.Y(n_3772)
);

OAI22xp5_ASAP7_75t_L g3773 ( 
.A1(n_3324),
.A2(n_861),
.B1(n_862),
.B2(n_860),
.Y(n_3773)
);

AOI221xp5_ASAP7_75t_L g3774 ( 
.A1(n_3378),
.A2(n_862),
.B1(n_863),
.B2(n_861),
.C(n_860),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3552),
.B(n_860),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3417),
.Y(n_3776)
);

INVx3_ASAP7_75t_SL g3777 ( 
.A(n_3464),
.Y(n_3777)
);

AOI21x1_ASAP7_75t_L g3778 ( 
.A1(n_3526),
.A2(n_863),
.B(n_862),
.Y(n_3778)
);

OAI21x1_ASAP7_75t_L g3779 ( 
.A1(n_3311),
.A2(n_865),
.B(n_864),
.Y(n_3779)
);

OAI22xp5_ASAP7_75t_L g3780 ( 
.A1(n_3372),
.A2(n_866),
.B1(n_867),
.B2(n_865),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3331),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3266),
.B(n_865),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3341),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3362),
.Y(n_3784)
);

O2A1O1Ixp33_ASAP7_75t_SL g3785 ( 
.A1(n_3332),
.A2(n_868),
.B(n_869),
.C(n_867),
.Y(n_3785)
);

OAI21x1_ASAP7_75t_L g3786 ( 
.A1(n_3312),
.A2(n_868),
.B(n_867),
.Y(n_3786)
);

INVx1_ASAP7_75t_SL g3787 ( 
.A(n_3321),
.Y(n_3787)
);

NAND2xp33_ASAP7_75t_R g3788 ( 
.A(n_3370),
.B(n_1075),
.Y(n_3788)
);

OA21x2_ASAP7_75t_L g3789 ( 
.A1(n_3430),
.A2(n_3431),
.B(n_3229),
.Y(n_3789)
);

NAND3x1_ASAP7_75t_L g3790 ( 
.A(n_3303),
.B(n_869),
.C(n_868),
.Y(n_3790)
);

BUFx12f_ASAP7_75t_L g3791 ( 
.A(n_3409),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3262),
.B(n_875),
.Y(n_3792)
);

OAI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3551),
.A2(n_877),
.B(n_876),
.Y(n_3793)
);

OAI21x1_ASAP7_75t_SL g3794 ( 
.A1(n_3375),
.A2(n_878),
.B(n_877),
.Y(n_3794)
);

INVx3_ASAP7_75t_L g3795 ( 
.A(n_3503),
.Y(n_3795)
);

OR2x2_ASAP7_75t_L g3796 ( 
.A(n_3285),
.B(n_878),
.Y(n_3796)
);

AOI21xp5_ASAP7_75t_L g3797 ( 
.A1(n_3261),
.A2(n_880),
.B(n_879),
.Y(n_3797)
);

AO32x2_ASAP7_75t_L g3798 ( 
.A1(n_3388),
.A2(n_895),
.A3(n_903),
.B1(n_887),
.B2(n_880),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3421),
.B(n_879),
.Y(n_3799)
);

OA21x2_ASAP7_75t_L g3800 ( 
.A1(n_3514),
.A2(n_882),
.B(n_881),
.Y(n_3800)
);

NOR2xp33_ASAP7_75t_L g3801 ( 
.A(n_3244),
.B(n_882),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3294),
.Y(n_3802)
);

OA21x2_ASAP7_75t_L g3803 ( 
.A1(n_3565),
.A2(n_885),
.B(n_884),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3365),
.B(n_884),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3293),
.B(n_885),
.Y(n_3805)
);

OAI21x1_ASAP7_75t_L g3806 ( 
.A1(n_3344),
.A2(n_887),
.B(n_886),
.Y(n_3806)
);

NOR3xp33_ASAP7_75t_L g3807 ( 
.A(n_3425),
.B(n_897),
.C(n_889),
.Y(n_3807)
);

A2O1A1Ixp33_ASAP7_75t_L g3808 ( 
.A1(n_3351),
.A2(n_889),
.B(n_890),
.C(n_888),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3510),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3295),
.B(n_888),
.Y(n_3810)
);

AOI221x1_ASAP7_75t_L g3811 ( 
.A1(n_3515),
.A2(n_893),
.B1(n_894),
.B2(n_892),
.C(n_891),
.Y(n_3811)
);

AOI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_3589),
.A2(n_894),
.B(n_893),
.Y(n_3812)
);

BUFx6f_ASAP7_75t_L g3813 ( 
.A(n_3493),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_SL g3814 ( 
.A(n_3411),
.B(n_895),
.Y(n_3814)
);

OAI22xp5_ASAP7_75t_L g3815 ( 
.A1(n_3379),
.A2(n_898),
.B1(n_899),
.B2(n_897),
.Y(n_3815)
);

OAI21x1_ASAP7_75t_L g3816 ( 
.A1(n_3347),
.A2(n_901),
.B(n_900),
.Y(n_3816)
);

AO21x1_ASAP7_75t_L g3817 ( 
.A1(n_3419),
.A2(n_902),
.B(n_900),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_R g3818 ( 
.A(n_3585),
.B(n_902),
.Y(n_3818)
);

OAI21x1_ASAP7_75t_L g3819 ( 
.A1(n_3469),
.A2(n_905),
.B(n_904),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3301),
.B(n_904),
.Y(n_3820)
);

OAI21x1_ASAP7_75t_L g3821 ( 
.A1(n_3546),
.A2(n_3549),
.B(n_3547),
.Y(n_3821)
);

NAND3xp33_ASAP7_75t_L g3822 ( 
.A(n_3500),
.B(n_906),
.C(n_905),
.Y(n_3822)
);

OAI21x1_ASAP7_75t_SL g3823 ( 
.A1(n_3320),
.A2(n_906),
.B(n_905),
.Y(n_3823)
);

A2O1A1Ixp33_ASAP7_75t_L g3824 ( 
.A1(n_3491),
.A2(n_907),
.B(n_908),
.C(n_906),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3540),
.B(n_907),
.Y(n_3825)
);

OAI21x1_ASAP7_75t_SL g3826 ( 
.A1(n_3407),
.A2(n_909),
.B(n_908),
.Y(n_3826)
);

OAI21x1_ASAP7_75t_L g3827 ( 
.A1(n_3553),
.A2(n_3554),
.B(n_3281),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3589),
.A2(n_910),
.B(n_909),
.Y(n_3828)
);

AO31x2_ASAP7_75t_L g3829 ( 
.A1(n_3451),
.A2(n_911),
.A3(n_912),
.B(n_910),
.Y(n_3829)
);

AOI21xp5_ASAP7_75t_L g3830 ( 
.A1(n_3589),
.A2(n_911),
.B(n_910),
.Y(n_3830)
);

AO22x2_ASAP7_75t_L g3831 ( 
.A1(n_3414),
.A2(n_912),
.B1(n_913),
.B2(n_911),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3525),
.B(n_913),
.Y(n_3832)
);

INVx3_ASAP7_75t_L g3833 ( 
.A(n_3232),
.Y(n_3833)
);

A2O1A1Ixp33_ASAP7_75t_L g3834 ( 
.A1(n_3542),
.A2(n_914),
.B(n_915),
.C(n_913),
.Y(n_3834)
);

OAI21x1_ASAP7_75t_L g3835 ( 
.A1(n_3373),
.A2(n_916),
.B(n_915),
.Y(n_3835)
);

OAI22x1_ASAP7_75t_L g3836 ( 
.A1(n_3322),
.A2(n_916),
.B1(n_917),
.B2(n_915),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3294),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3392),
.A2(n_918),
.B(n_917),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3315),
.Y(n_3839)
);

A2O1A1Ixp33_ASAP7_75t_L g3840 ( 
.A1(n_3438),
.A2(n_919),
.B(n_920),
.C(n_918),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3602),
.Y(n_3841)
);

OAI21x1_ASAP7_75t_L g3842 ( 
.A1(n_3389),
.A2(n_920),
.B(n_919),
.Y(n_3842)
);

INVx2_ASAP7_75t_SL g3843 ( 
.A(n_3254),
.Y(n_3843)
);

OAI21x1_ASAP7_75t_L g3844 ( 
.A1(n_3398),
.A2(n_921),
.B(n_920),
.Y(n_3844)
);

NOR2xp33_ASAP7_75t_L g3845 ( 
.A(n_3288),
.B(n_921),
.Y(n_3845)
);

AND2x6_ASAP7_75t_L g3846 ( 
.A(n_3254),
.B(n_921),
.Y(n_3846)
);

NAND3xp33_ASAP7_75t_L g3847 ( 
.A(n_3501),
.B(n_3495),
.C(n_3487),
.Y(n_3847)
);

INVx3_ASAP7_75t_L g3848 ( 
.A(n_3296),
.Y(n_3848)
);

INVx4_ASAP7_75t_L g3849 ( 
.A(n_3296),
.Y(n_3849)
);

AOI21xp33_ASAP7_75t_L g3850 ( 
.A1(n_3272),
.A2(n_3279),
.B(n_3470),
.Y(n_3850)
);

NOR2xp33_ASAP7_75t_SL g3851 ( 
.A(n_3573),
.B(n_924),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3287),
.B(n_924),
.Y(n_3852)
);

O2A1O1Ixp33_ASAP7_75t_L g3853 ( 
.A1(n_3400),
.A2(n_926),
.B(n_927),
.C(n_925),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3530),
.B(n_925),
.Y(n_3854)
);

AOI21xp5_ASAP7_75t_L g3855 ( 
.A1(n_3371),
.A2(n_926),
.B(n_925),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3562),
.Y(n_3856)
);

BUFx6f_ASAP7_75t_L g3857 ( 
.A(n_3227),
.Y(n_3857)
);

OR2x6_ASAP7_75t_L g3858 ( 
.A(n_3433),
.B(n_926),
.Y(n_3858)
);

OA21x2_ASAP7_75t_L g3859 ( 
.A1(n_3436),
.A2(n_928),
.B(n_927),
.Y(n_3859)
);

INVx8_ASAP7_75t_L g3860 ( 
.A(n_3289),
.Y(n_3860)
);

INVx3_ASAP7_75t_L g3861 ( 
.A(n_3289),
.Y(n_3861)
);

INVx2_ASAP7_75t_SL g3862 ( 
.A(n_3227),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_SL g3863 ( 
.A1(n_3450),
.A2(n_3462),
.B(n_3449),
.Y(n_3863)
);

OAI21x1_ASAP7_75t_L g3864 ( 
.A1(n_3429),
.A2(n_928),
.B(n_927),
.Y(n_3864)
);

O2A1O1Ixp5_ASAP7_75t_L g3865 ( 
.A1(n_3524),
.A2(n_929),
.B(n_930),
.C(n_928),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3545),
.B(n_929),
.Y(n_3866)
);

BUFx6f_ASAP7_75t_L g3867 ( 
.A(n_3227),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_3371),
.Y(n_3868)
);

BUFx2_ASAP7_75t_L g3869 ( 
.A(n_3236),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3581),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3581),
.Y(n_3871)
);

INVx3_ASAP7_75t_SL g3872 ( 
.A(n_3371),
.Y(n_3872)
);

NOR2xp67_ASAP7_75t_L g3873 ( 
.A(n_3337),
.B(n_3313),
.Y(n_3873)
);

INVx1_ASAP7_75t_SL g3874 ( 
.A(n_3465),
.Y(n_3874)
);

NAND3xp33_ASAP7_75t_SL g3875 ( 
.A(n_3276),
.B(n_57),
.C(n_58),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3359),
.B(n_931),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3383),
.B(n_931),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_3453),
.B(n_932),
.Y(n_3878)
);

OAI22xp5_ASAP7_75t_L g3879 ( 
.A1(n_3490),
.A2(n_3483),
.B1(n_3448),
.B2(n_3488),
.Y(n_3879)
);

OAI21x1_ASAP7_75t_L g3880 ( 
.A1(n_3441),
.A2(n_934),
.B(n_933),
.Y(n_3880)
);

OAI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3578),
.A2(n_3576),
.B(n_3555),
.Y(n_3881)
);

OAI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3544),
.A2(n_936),
.B(n_935),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3393),
.B(n_936),
.Y(n_3883)
);

INVx2_ASAP7_75t_SL g3884 ( 
.A(n_3236),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3401),
.B(n_937),
.Y(n_3885)
);

AOI221xp5_ASAP7_75t_SL g3886 ( 
.A1(n_3369),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.C(n_61),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_3472),
.A2(n_938),
.B(n_937),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3444),
.B(n_3556),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3482),
.A2(n_940),
.B(n_939),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_3517),
.B(n_940),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3508),
.B(n_940),
.Y(n_3891)
);

AOI22xp33_ASAP7_75t_L g3892 ( 
.A1(n_3340),
.A2(n_942),
.B1(n_943),
.B2(n_941),
.Y(n_3892)
);

AOI31xp67_ASAP7_75t_L g3893 ( 
.A1(n_3604),
.A2(n_3382),
.A3(n_3405),
.B(n_3368),
.Y(n_3893)
);

CKINVDCx20_ASAP7_75t_R g3894 ( 
.A(n_3696),
.Y(n_3894)
);

AOI221xp5_ASAP7_75t_L g3895 ( 
.A1(n_3639),
.A2(n_3364),
.B1(n_3390),
.B2(n_3376),
.C(n_3456),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3847),
.A2(n_3563),
.B1(n_3366),
.B2(n_3559),
.Y(n_3896)
);

OAI21x1_ASAP7_75t_L g3897 ( 
.A1(n_3656),
.A2(n_3355),
.B(n_3443),
.Y(n_3897)
);

AOI222xp33_ASAP7_75t_SL g3898 ( 
.A1(n_3647),
.A2(n_3577),
.B1(n_3586),
.B2(n_3534),
.C1(n_3533),
.C2(n_3539),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3690),
.Y(n_3899)
);

BUFx6f_ASAP7_75t_L g3900 ( 
.A(n_3680),
.Y(n_3900)
);

OAI211xp5_ASAP7_75t_L g3901 ( 
.A1(n_3611),
.A2(n_3538),
.B(n_3504),
.C(n_3566),
.Y(n_3901)
);

O2A1O1Ixp33_ASAP7_75t_SL g3902 ( 
.A1(n_3657),
.A2(n_3592),
.B(n_3564),
.C(n_3571),
.Y(n_3902)
);

AO21x2_ASAP7_75t_L g3903 ( 
.A1(n_3797),
.A2(n_3452),
.B(n_3402),
.Y(n_3903)
);

OAI21x1_ASAP7_75t_L g3904 ( 
.A1(n_3619),
.A2(n_3509),
.B(n_3505),
.Y(n_3904)
);

OAI21x1_ASAP7_75t_L g3905 ( 
.A1(n_3675),
.A2(n_3494),
.B(n_3297),
.Y(n_3905)
);

AND2x2_ASAP7_75t_SL g3906 ( 
.A(n_3734),
.B(n_3236),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3873),
.A2(n_3879),
.B1(n_3807),
.B2(n_3851),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3614),
.Y(n_3908)
);

INVx6_ASAP7_75t_L g3909 ( 
.A(n_3709),
.Y(n_3909)
);

OR2x2_ASAP7_75t_L g3910 ( 
.A(n_3651),
.B(n_3496),
.Y(n_3910)
);

OAI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3748),
.A2(n_3588),
.B1(n_3511),
.B2(n_3590),
.Y(n_3911)
);

OAI22xp33_ASAP7_75t_L g3912 ( 
.A1(n_3788),
.A2(n_3570),
.B1(n_3574),
.B2(n_3568),
.Y(n_3912)
);

AO31x2_ASAP7_75t_L g3913 ( 
.A1(n_3640),
.A2(n_3316),
.A3(n_3477),
.B(n_3475),
.Y(n_3913)
);

AOI21x1_ASAP7_75t_L g3914 ( 
.A1(n_3686),
.A2(n_3484),
.B(n_3455),
.Y(n_3914)
);

O2A1O1Ixp33_ASAP7_75t_SL g3915 ( 
.A1(n_3607),
.A2(n_3580),
.B(n_3583),
.C(n_3557),
.Y(n_3915)
);

INVx3_ASAP7_75t_L g3916 ( 
.A(n_3681),
.Y(n_3916)
);

OAI21x1_ASAP7_75t_L g3917 ( 
.A1(n_3626),
.A2(n_3298),
.B(n_3291),
.Y(n_3917)
);

OAI21x1_ASAP7_75t_L g3918 ( 
.A1(n_3739),
.A2(n_3302),
.B(n_3600),
.Y(n_3918)
);

AOI221xp5_ASAP7_75t_L g3919 ( 
.A1(n_3643),
.A2(n_3446),
.B1(n_3434),
.B2(n_3439),
.C(n_3498),
.Y(n_3919)
);

INVx1_ASAP7_75t_SL g3920 ( 
.A(n_3777),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3754),
.B(n_3535),
.Y(n_3921)
);

NAND2x1p5_ASAP7_75t_L g3922 ( 
.A(n_3630),
.B(n_3486),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3856),
.B(n_3502),
.Y(n_3923)
);

OAI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3637),
.A2(n_3426),
.B(n_3593),
.Y(n_3924)
);

OAI21xp5_ASAP7_75t_L g3925 ( 
.A1(n_3762),
.A2(n_3532),
.B(n_3518),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3645),
.Y(n_3926)
);

AO31x2_ASAP7_75t_L g3927 ( 
.A1(n_3869),
.A2(n_3541),
.A3(n_3594),
.B(n_3582),
.Y(n_3927)
);

AO21x2_ASAP7_75t_L g3928 ( 
.A1(n_3716),
.A2(n_3548),
.B(n_3442),
.Y(n_3928)
);

OAI21x1_ASAP7_75t_L g3929 ( 
.A1(n_3692),
.A2(n_3397),
.B(n_3440),
.Y(n_3929)
);

NOR2x1_ASAP7_75t_R g3930 ( 
.A(n_3664),
.B(n_3243),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3606),
.B(n_3486),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3761),
.B(n_3486),
.Y(n_3932)
);

AOI221xp5_ASAP7_75t_L g3933 ( 
.A1(n_3801),
.A2(n_3499),
.B1(n_3308),
.B2(n_3243),
.C(n_3492),
.Y(n_3933)
);

AOI21x1_ASAP7_75t_L g3934 ( 
.A1(n_3763),
.A2(n_3308),
.B(n_3499),
.Y(n_3934)
);

OAI22xp5_ASAP7_75t_L g3935 ( 
.A1(n_3698),
.A2(n_3492),
.B1(n_3243),
.B2(n_942),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3625),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3648),
.Y(n_3937)
);

NAND2x1p5_ASAP7_75t_L g3938 ( 
.A(n_3699),
.B(n_3492),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3660),
.Y(n_3939)
);

AOI22xp33_ASAP7_75t_SL g3940 ( 
.A1(n_3818),
.A2(n_942),
.B1(n_943),
.B2(n_941),
.Y(n_3940)
);

OAI21x1_ASAP7_75t_L g3941 ( 
.A1(n_3659),
.A2(n_944),
.B(n_943),
.Y(n_3941)
);

BUFx8_ASAP7_75t_L g3942 ( 
.A(n_3670),
.Y(n_3942)
);

OA21x2_ASAP7_75t_L g3943 ( 
.A1(n_3767),
.A2(n_3850),
.B(n_3635),
.Y(n_3943)
);

CKINVDCx16_ASAP7_75t_R g3944 ( 
.A(n_3627),
.Y(n_3944)
);

INVx2_ASAP7_75t_SL g3945 ( 
.A(n_3663),
.Y(n_3945)
);

INVx3_ASAP7_75t_L g3946 ( 
.A(n_3655),
.Y(n_3946)
);

AO31x2_ASAP7_75t_L g3947 ( 
.A1(n_3802),
.A2(n_1089),
.A3(n_946),
.B(n_947),
.Y(n_3947)
);

OAI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_3822),
.A2(n_948),
.B(n_947),
.Y(n_3948)
);

OAI21x1_ASAP7_75t_L g3949 ( 
.A1(n_3605),
.A2(n_949),
.B(n_948),
.Y(n_3949)
);

OAI221xp5_ASAP7_75t_L g3950 ( 
.A1(n_3644),
.A2(n_951),
.B1(n_952),
.B2(n_950),
.C(n_949),
.Y(n_3950)
);

BUFx2_ASAP7_75t_L g3951 ( 
.A(n_3717),
.Y(n_3951)
);

AND2x4_ASAP7_75t_L g3952 ( 
.A(n_3755),
.B(n_3760),
.Y(n_3952)
);

OAI21xp5_ASAP7_75t_L g3953 ( 
.A1(n_3674),
.A2(n_953),
.B(n_952),
.Y(n_3953)
);

INVx8_ASAP7_75t_L g3954 ( 
.A(n_3860),
.Y(n_3954)
);

OAI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3641),
.A2(n_954),
.B(n_953),
.Y(n_3955)
);

INVx4_ASAP7_75t_L g3956 ( 
.A(n_3652),
.Y(n_3956)
);

AOI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3863),
.A2(n_954),
.B(n_953),
.Y(n_3957)
);

AO31x2_ASAP7_75t_L g3958 ( 
.A1(n_3837),
.A2(n_956),
.A3(n_957),
.B(n_955),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3704),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3705),
.Y(n_3960)
);

BUFx2_ASAP7_75t_L g3961 ( 
.A(n_3872),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3706),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3730),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3735),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3740),
.Y(n_3965)
);

OA21x2_ASAP7_75t_L g3966 ( 
.A1(n_3616),
.A2(n_3615),
.B(n_3733),
.Y(n_3966)
);

OA21x2_ASAP7_75t_L g3967 ( 
.A1(n_3725),
.A2(n_961),
.B(n_959),
.Y(n_3967)
);

INVxp33_ASAP7_75t_L g3968 ( 
.A(n_3813),
.Y(n_3968)
);

O2A1O1Ixp33_ASAP7_75t_SL g3969 ( 
.A1(n_3715),
.A2(n_3765),
.B(n_3629),
.C(n_3669),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3745),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3764),
.Y(n_3971)
);

INVx1_ASAP7_75t_SL g3972 ( 
.A(n_3756),
.Y(n_3972)
);

BUFx2_ASAP7_75t_L g3973 ( 
.A(n_3868),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3759),
.Y(n_3974)
);

OAI21x1_ASAP7_75t_L g3975 ( 
.A1(n_3646),
.A2(n_963),
.B(n_962),
.Y(n_3975)
);

OAI21x1_ASAP7_75t_L g3976 ( 
.A1(n_3688),
.A2(n_964),
.B(n_963),
.Y(n_3976)
);

BUFx2_ASAP7_75t_L g3977 ( 
.A(n_3870),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3871),
.Y(n_3978)
);

NOR2x1_ASAP7_75t_SL g3979 ( 
.A(n_3849),
.B(n_965),
.Y(n_3979)
);

AO21x2_ASAP7_75t_L g3980 ( 
.A1(n_3724),
.A2(n_967),
.B(n_966),
.Y(n_3980)
);

AO21x2_ASAP7_75t_L g3981 ( 
.A1(n_3771),
.A2(n_3778),
.B(n_3875),
.Y(n_3981)
);

OAI21x1_ASAP7_75t_L g3982 ( 
.A1(n_3827),
.A2(n_967),
.B(n_966),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3839),
.Y(n_3983)
);

NAND2xp33_ASAP7_75t_L g3984 ( 
.A(n_3846),
.B(n_968),
.Y(n_3984)
);

AOI22xp33_ASAP7_75t_L g3985 ( 
.A1(n_3672),
.A2(n_969),
.B1(n_970),
.B2(n_968),
.Y(n_3985)
);

OAI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3858),
.A2(n_972),
.B1(n_973),
.B2(n_971),
.Y(n_3986)
);

OA21x2_ASAP7_75t_L g3987 ( 
.A1(n_3701),
.A2(n_973),
.B(n_972),
.Y(n_3987)
);

NOR2xp67_ASAP7_75t_SL g3988 ( 
.A(n_3694),
.B(n_975),
.Y(n_3988)
);

INVx2_ASAP7_75t_SL g3989 ( 
.A(n_3791),
.Y(n_3989)
);

NOR2xp67_ASAP7_75t_L g3990 ( 
.A(n_3795),
.B(n_978),
.Y(n_3990)
);

AO32x2_ASAP7_75t_L g3991 ( 
.A1(n_3718),
.A2(n_980),
.A3(n_981),
.B1(n_979),
.B2(n_978),
.Y(n_3991)
);

AO32x2_ASAP7_75t_L g3992 ( 
.A1(n_3766),
.A2(n_980),
.A3(n_981),
.B1(n_979),
.B2(n_978),
.Y(n_3992)
);

CKINVDCx20_ASAP7_75t_R g3993 ( 
.A(n_3678),
.Y(n_3993)
);

AOI21xp5_ASAP7_75t_L g3994 ( 
.A1(n_3874),
.A2(n_983),
.B(n_982),
.Y(n_3994)
);

OAI21x1_ASAP7_75t_L g3995 ( 
.A1(n_3653),
.A2(n_983),
.B(n_982),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3776),
.Y(n_3996)
);

INVx2_ASAP7_75t_SL g3997 ( 
.A(n_3860),
.Y(n_3997)
);

AOI22xp33_ASAP7_75t_L g3998 ( 
.A1(n_3672),
.A2(n_985),
.B1(n_986),
.B2(n_984),
.Y(n_3998)
);

AO21x2_ASAP7_75t_L g3999 ( 
.A1(n_3633),
.A2(n_987),
.B(n_986),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3617),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3796),
.Y(n_4001)
);

NOR2xp67_ASAP7_75t_L g4002 ( 
.A(n_3610),
.B(n_988),
.Y(n_4002)
);

NAND3xp33_ASAP7_75t_L g4003 ( 
.A(n_3886),
.B(n_989),
.C(n_988),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3672),
.A2(n_991),
.B1(n_992),
.B2(n_990),
.Y(n_4004)
);

O2A1O1Ixp33_ASAP7_75t_SL g4005 ( 
.A1(n_3834),
.A2(n_991),
.B(n_992),
.C(n_990),
.Y(n_4005)
);

OAI21x1_ASAP7_75t_L g4006 ( 
.A1(n_3751),
.A2(n_3697),
.B(n_3693),
.Y(n_4006)
);

INVx4_ASAP7_75t_L g4007 ( 
.A(n_3649),
.Y(n_4007)
);

NOR2x1_ASAP7_75t_SL g4008 ( 
.A(n_3628),
.B(n_994),
.Y(n_4008)
);

AO21x2_ASAP7_75t_L g4009 ( 
.A1(n_3702),
.A2(n_996),
.B(n_995),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3617),
.Y(n_4010)
);

OAI21x1_ASAP7_75t_L g4011 ( 
.A1(n_3821),
.A2(n_998),
.B(n_997),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3621),
.Y(n_4012)
);

BUFx6f_ASAP7_75t_L g4013 ( 
.A(n_3857),
.Y(n_4013)
);

OAI21x1_ASAP7_75t_L g4014 ( 
.A1(n_3731),
.A2(n_999),
.B(n_998),
.Y(n_4014)
);

OAI21x1_ASAP7_75t_L g4015 ( 
.A1(n_3708),
.A2(n_1002),
.B(n_1001),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_3809),
.Y(n_4016)
);

OAI21x1_ASAP7_75t_L g4017 ( 
.A1(n_3711),
.A2(n_1003),
.B(n_1002),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3621),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3841),
.B(n_1004),
.Y(n_4019)
);

AO32x2_ASAP7_75t_L g4020 ( 
.A1(n_3843),
.A2(n_1006),
.A3(n_1007),
.B1(n_1005),
.B2(n_1004),
.Y(n_4020)
);

INVx1_ASAP7_75t_SL g4021 ( 
.A(n_3787),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3621),
.Y(n_4022)
);

OAI21x1_ASAP7_75t_L g4023 ( 
.A1(n_3835),
.A2(n_1008),
.B(n_1007),
.Y(n_4023)
);

CKINVDCx6p67_ASAP7_75t_R g4024 ( 
.A(n_3846),
.Y(n_4024)
);

AO31x2_ASAP7_75t_L g4025 ( 
.A1(n_3817),
.A2(n_1084),
.A3(n_1008),
.B(n_1009),
.Y(n_4025)
);

INVx8_ASAP7_75t_L g4026 ( 
.A(n_3846),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3631),
.Y(n_4027)
);

OAI21x1_ASAP7_75t_L g4028 ( 
.A1(n_3842),
.A2(n_1011),
.B(n_1010),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3631),
.Y(n_4029)
);

AO32x2_ASAP7_75t_L g4030 ( 
.A1(n_3773),
.A2(n_1013),
.A3(n_1014),
.B1(n_1012),
.B2(n_1011),
.Y(n_4030)
);

OAI21x1_ASAP7_75t_L g4031 ( 
.A1(n_3844),
.A2(n_1013),
.B(n_1012),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3781),
.B(n_1083),
.Y(n_4032)
);

OAI21x1_ASAP7_75t_L g4033 ( 
.A1(n_3848),
.A2(n_1013),
.B(n_1012),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3833),
.Y(n_4034)
);

NOR2x1_ASAP7_75t_R g4035 ( 
.A(n_3612),
.B(n_3695),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3784),
.Y(n_4036)
);

AO31x2_ASAP7_75t_L g4037 ( 
.A1(n_3811),
.A2(n_1083),
.A3(n_1017),
.B(n_1018),
.Y(n_4037)
);

AO31x2_ASAP7_75t_L g4038 ( 
.A1(n_3671),
.A2(n_1020),
.A3(n_1021),
.B(n_1019),
.Y(n_4038)
);

AO21x2_ASAP7_75t_L g4039 ( 
.A1(n_3613),
.A2(n_1021),
.B(n_1020),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3783),
.B(n_3888),
.Y(n_4040)
);

OAI21x1_ASAP7_75t_SL g4041 ( 
.A1(n_3826),
.A2(n_1021),
.B(n_1020),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3679),
.B(n_1083),
.Y(n_4042)
);

AOI22xp33_ASAP7_75t_L g4043 ( 
.A1(n_3831),
.A2(n_3729),
.B1(n_3845),
.B2(n_3752),
.Y(n_4043)
);

OA21x2_ASAP7_75t_L g4044 ( 
.A1(n_3603),
.A2(n_1023),
.B(n_1022),
.Y(n_4044)
);

BUFx3_ASAP7_75t_L g4045 ( 
.A(n_3742),
.Y(n_4045)
);

NOR2xp33_ASAP7_75t_L g4046 ( 
.A(n_3632),
.B(n_62),
.Y(n_4046)
);

INVx2_ASAP7_75t_L g4047 ( 
.A(n_3862),
.Y(n_4047)
);

AND2x4_ASAP7_75t_L g4048 ( 
.A(n_3861),
.B(n_1022),
.Y(n_4048)
);

CKINVDCx5p33_ASAP7_75t_R g4049 ( 
.A(n_3687),
.Y(n_4049)
);

OA21x2_ASAP7_75t_L g4050 ( 
.A1(n_3623),
.A2(n_1025),
.B(n_1024),
.Y(n_4050)
);

BUFx6f_ASAP7_75t_L g4051 ( 
.A(n_3867),
.Y(n_4051)
);

OAI21x1_ASAP7_75t_L g4052 ( 
.A1(n_3741),
.A2(n_1025),
.B(n_1024),
.Y(n_4052)
);

OA21x2_ASAP7_75t_L g4053 ( 
.A1(n_3753),
.A2(n_3828),
.B(n_3812),
.Y(n_4053)
);

OAI21xp5_ASAP7_75t_L g4054 ( 
.A1(n_3865),
.A2(n_1028),
.B(n_1027),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3831),
.A2(n_1028),
.B1(n_1029),
.B2(n_1027),
.Y(n_4055)
);

BUFx6f_ASAP7_75t_L g4056 ( 
.A(n_3867),
.Y(n_4056)
);

BUFx3_ASAP7_75t_L g4057 ( 
.A(n_3742),
.Y(n_4057)
);

OAI21x1_ASAP7_75t_L g4058 ( 
.A1(n_3769),
.A2(n_1030),
.B(n_1029),
.Y(n_4058)
);

OAI21x1_ASAP7_75t_L g4059 ( 
.A1(n_3819),
.A2(n_1032),
.B(n_1031),
.Y(n_4059)
);

OA21x2_ASAP7_75t_L g4060 ( 
.A1(n_3830),
.A2(n_1033),
.B(n_1032),
.Y(n_4060)
);

BUFx2_ASAP7_75t_L g4061 ( 
.A(n_3956),
.Y(n_4061)
);

OA21x2_ASAP7_75t_L g4062 ( 
.A1(n_4012),
.A2(n_3622),
.B(n_3799),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3908),
.Y(n_4063)
);

AND2x4_ASAP7_75t_L g4064 ( 
.A(n_4045),
.B(n_3884),
.Y(n_4064)
);

INVx3_ASAP7_75t_L g4065 ( 
.A(n_3954),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_L g4066 ( 
.A1(n_4017),
.A2(n_3634),
.B(n_3722),
.Y(n_4066)
);

OAI21x1_ASAP7_75t_SL g4067 ( 
.A1(n_3979),
.A2(n_3793),
.B(n_3794),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3926),
.Y(n_4068)
);

NOR2xp33_ASAP7_75t_L g4069 ( 
.A(n_3968),
.B(n_3668),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3931),
.B(n_3638),
.Y(n_4070)
);

OA21x2_ASAP7_75t_L g4071 ( 
.A1(n_4018),
.A2(n_3691),
.B(n_3684),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3899),
.Y(n_4072)
);

A2O1A1Ixp33_ASAP7_75t_L g4073 ( 
.A1(n_3906),
.A2(n_4002),
.B(n_3984),
.C(n_3988),
.Y(n_4073)
);

AND2x2_ASAP7_75t_L g4074 ( 
.A(n_3951),
.B(n_3676),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_3907),
.A2(n_3790),
.B1(n_3667),
.B2(n_3666),
.Y(n_4075)
);

AO21x2_ASAP7_75t_L g4076 ( 
.A1(n_4022),
.A2(n_3723),
.B(n_3703),
.Y(n_4076)
);

OAI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_4024),
.A2(n_3609),
.B1(n_3840),
.B2(n_3814),
.Y(n_4077)
);

OAI21xp5_ASAP7_75t_L g4078 ( 
.A1(n_3940),
.A2(n_3878),
.B(n_3642),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3951),
.B(n_3852),
.Y(n_4079)
);

CKINVDCx20_ASAP7_75t_R g4080 ( 
.A(n_3894),
.Y(n_4080)
);

OAI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_3957),
.A2(n_3853),
.B(n_3772),
.Y(n_4081)
);

OR2x2_ASAP7_75t_L g4082 ( 
.A(n_3977),
.B(n_3936),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3939),
.B(n_4036),
.Y(n_4083)
);

AND2x4_ASAP7_75t_L g4084 ( 
.A(n_4057),
.B(n_3728),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_3961),
.B(n_3728),
.Y(n_4085)
);

AOI22x1_ASAP7_75t_L g4086 ( 
.A1(n_3944),
.A2(n_3836),
.B1(n_3747),
.B2(n_3804),
.Y(n_4086)
);

AOI21xp5_ASAP7_75t_L g4087 ( 
.A1(n_3915),
.A2(n_3785),
.B(n_3789),
.Y(n_4087)
);

AOI21x1_ASAP7_75t_L g4088 ( 
.A1(n_3990),
.A2(n_3743),
.B(n_3650),
.Y(n_4088)
);

AOI221x1_ASAP7_75t_SL g4089 ( 
.A1(n_3912),
.A2(n_3866),
.B1(n_3854),
.B2(n_3832),
.C(n_3877),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_4043),
.A2(n_3803),
.B1(n_3750),
.B2(n_3881),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3971),
.Y(n_4091)
);

AO31x2_ASAP7_75t_L g4092 ( 
.A1(n_4027),
.A2(n_3608),
.A3(n_3618),
.B(n_3838),
.Y(n_4092)
);

INVx4_ASAP7_75t_SL g4093 ( 
.A(n_3909),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3974),
.B(n_3719),
.Y(n_4094)
);

OA21x2_ASAP7_75t_L g4095 ( 
.A1(n_4029),
.A2(n_3683),
.B(n_3682),
.Y(n_4095)
);

OA21x2_ASAP7_75t_L g4096 ( 
.A1(n_4000),
.A2(n_3658),
.B(n_3654),
.Y(n_4096)
);

INVx2_ASAP7_75t_L g4097 ( 
.A(n_3937),
.Y(n_4097)
);

OA21x2_ASAP7_75t_L g4098 ( 
.A1(n_4010),
.A2(n_3661),
.B(n_3685),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3960),
.Y(n_4099)
);

AOI21x1_ASAP7_75t_L g4100 ( 
.A1(n_3914),
.A2(n_3689),
.B(n_3859),
.Y(n_4100)
);

BUFx8_ASAP7_75t_L g4101 ( 
.A(n_3989),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_SL g4102 ( 
.A1(n_4026),
.A2(n_3803),
.B1(n_3859),
.B2(n_3823),
.Y(n_4102)
);

AOI22xp33_ASAP7_75t_SL g4103 ( 
.A1(n_4026),
.A2(n_3768),
.B1(n_3732),
.B2(n_3882),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3964),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3965),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3959),
.Y(n_4106)
);

OA21x2_ASAP7_75t_L g4107 ( 
.A1(n_3970),
.A2(n_3673),
.B(n_3662),
.Y(n_4107)
);

AO31x2_ASAP7_75t_L g4108 ( 
.A1(n_3973),
.A2(n_3712),
.A3(n_3713),
.B(n_3700),
.Y(n_4108)
);

HB1xp67_ASAP7_75t_L g4109 ( 
.A(n_4021),
.Y(n_4109)
);

AO21x2_ASAP7_75t_L g4110 ( 
.A1(n_3955),
.A2(n_3721),
.B(n_3714),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3962),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3963),
.Y(n_4112)
);

OAI21x1_ASAP7_75t_L g4113 ( 
.A1(n_4006),
.A2(n_3786),
.B(n_3779),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_4001),
.B(n_3727),
.Y(n_4114)
);

AO31x2_ASAP7_75t_L g4115 ( 
.A1(n_3973),
.A2(n_3736),
.A3(n_3738),
.B(n_3737),
.Y(n_4115)
);

BUFx4f_ASAP7_75t_SL g4116 ( 
.A(n_3993),
.Y(n_4116)
);

OAI21x1_ASAP7_75t_L g4117 ( 
.A1(n_3918),
.A2(n_3880),
.B(n_3864),
.Y(n_4117)
);

AO21x2_ASAP7_75t_L g4118 ( 
.A1(n_3948),
.A2(n_3775),
.B(n_3624),
.Y(n_4118)
);

AO21x2_ASAP7_75t_L g4119 ( 
.A1(n_3953),
.A2(n_3782),
.B(n_3620),
.Y(n_4119)
);

INVx3_ASAP7_75t_L g4120 ( 
.A(n_3916),
.Y(n_4120)
);

OA21x2_ASAP7_75t_L g4121 ( 
.A1(n_3897),
.A2(n_3810),
.B(n_3805),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_3978),
.Y(n_4122)
);

OAI21x1_ASAP7_75t_L g4123 ( 
.A1(n_3982),
.A2(n_3904),
.B(n_3929),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_4016),
.Y(n_4124)
);

AOI21xp5_ASAP7_75t_L g4125 ( 
.A1(n_4035),
.A2(n_3707),
.B(n_3749),
.Y(n_4125)
);

OAI21x1_ASAP7_75t_L g4126 ( 
.A1(n_3905),
.A2(n_3816),
.B(n_3806),
.Y(n_4126)
);

HB1xp67_ASAP7_75t_L g4127 ( 
.A(n_3945),
.Y(n_4127)
);

AO31x2_ASAP7_75t_L g4128 ( 
.A1(n_4047),
.A2(n_3820),
.A3(n_3891),
.B(n_3876),
.Y(n_4128)
);

INVx6_ASAP7_75t_L g4129 ( 
.A(n_3900),
.Y(n_4129)
);

OR2x2_ASAP7_75t_L g4130 ( 
.A(n_3910),
.B(n_3726),
.Y(n_4130)
);

A2O1A1Ixp33_ASAP7_75t_L g4131 ( 
.A1(n_3946),
.A2(n_3774),
.B(n_3746),
.C(n_3744),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3996),
.Y(n_4132)
);

OAI21x1_ASAP7_75t_L g4133 ( 
.A1(n_4011),
.A2(n_3758),
.B(n_3757),
.Y(n_4133)
);

OAI21xp5_ASAP7_75t_L g4134 ( 
.A1(n_4003),
.A2(n_3808),
.B(n_3824),
.Y(n_4134)
);

OAI21x1_ASAP7_75t_L g4135 ( 
.A1(n_3941),
.A2(n_3800),
.B(n_3855),
.Y(n_4135)
);

NAND3xp33_ASAP7_75t_L g4136 ( 
.A(n_3943),
.B(n_3885),
.C(n_3883),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4034),
.B(n_3665),
.Y(n_4137)
);

AO31x2_ASAP7_75t_L g4138 ( 
.A1(n_3983),
.A2(n_3720),
.A3(n_3677),
.B(n_3792),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4040),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3932),
.Y(n_4140)
);

OAI21x1_ASAP7_75t_L g4141 ( 
.A1(n_3934),
.A2(n_3889),
.B(n_3887),
.Y(n_4141)
);

OAI22xp5_ASAP7_75t_L g4142 ( 
.A1(n_3896),
.A2(n_3892),
.B1(n_3890),
.B2(n_3825),
.Y(n_4142)
);

OA21x2_ASAP7_75t_L g4143 ( 
.A1(n_3925),
.A2(n_3815),
.B(n_3780),
.Y(n_4143)
);

AO31x2_ASAP7_75t_L g4144 ( 
.A1(n_4008),
.A2(n_3665),
.A3(n_3710),
.B(n_3798),
.Y(n_4144)
);

INVx2_ASAP7_75t_L g4145 ( 
.A(n_3938),
.Y(n_4145)
);

OAI21x1_ASAP7_75t_L g4146 ( 
.A1(n_3976),
.A2(n_3636),
.B(n_3726),
.Y(n_4146)
);

HB1xp67_ASAP7_75t_L g4147 ( 
.A(n_3972),
.Y(n_4147)
);

AO31x2_ASAP7_75t_L g4148 ( 
.A1(n_3935),
.A2(n_3710),
.A3(n_3798),
.B(n_3636),
.Y(n_4148)
);

OAI21x1_ASAP7_75t_L g4149 ( 
.A1(n_3995),
.A2(n_3770),
.B(n_3829),
.Y(n_4149)
);

AOI21xp5_ASAP7_75t_L g4150 ( 
.A1(n_3969),
.A2(n_3798),
.B(n_3770),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3902),
.A2(n_4005),
.B(n_3981),
.Y(n_4151)
);

AO21x2_ASAP7_75t_L g4152 ( 
.A1(n_4019),
.A2(n_3829),
.B(n_3770),
.Y(n_4152)
);

BUFx3_ASAP7_75t_L g4153 ( 
.A(n_3942),
.Y(n_4153)
);

OAI21x1_ASAP7_75t_L g4154 ( 
.A1(n_3975),
.A2(n_3922),
.B(n_3924),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4082),
.Y(n_4155)
);

INVxp67_ASAP7_75t_L g4156 ( 
.A(n_4061),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_4072),
.Y(n_4157)
);

BUFx2_ASAP7_75t_L g4158 ( 
.A(n_4093),
.Y(n_4158)
);

CKINVDCx6p67_ASAP7_75t_R g4159 ( 
.A(n_4153),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_4079),
.B(n_3920),
.Y(n_4160)
);

HB1xp67_ASAP7_75t_L g4161 ( 
.A(n_4147),
.Y(n_4161)
);

HB1xp67_ASAP7_75t_L g4162 ( 
.A(n_4127),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4063),
.Y(n_4163)
);

BUFx2_ASAP7_75t_SL g4164 ( 
.A(n_4065),
.Y(n_4164)
);

AO21x1_ASAP7_75t_SL g4165 ( 
.A1(n_4109),
.A2(n_3930),
.B(n_3985),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_4097),
.Y(n_4166)
);

INVx4_ASAP7_75t_L g4167 ( 
.A(n_4093),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4068),
.Y(n_4168)
);

HB1xp67_ASAP7_75t_L g4169 ( 
.A(n_4111),
.Y(n_4169)
);

BUFx2_ASAP7_75t_L g4170 ( 
.A(n_4101),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_L g4171 ( 
.A1(n_4086),
.A2(n_3911),
.B1(n_3950),
.B2(n_3903),
.Y(n_4171)
);

AO21x2_ASAP7_75t_L g4172 ( 
.A1(n_4151),
.A2(n_4032),
.B(n_3928),
.Y(n_4172)
);

OA21x2_ASAP7_75t_L g4173 ( 
.A1(n_4150),
.A2(n_3921),
.B(n_3923),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4099),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4104),
.Y(n_4175)
);

OR2x2_ASAP7_75t_L g4176 ( 
.A(n_4139),
.B(n_4083),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_4124),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4105),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_4091),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_4070),
.B(n_3952),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4106),
.Y(n_4181)
);

INVx3_ASAP7_75t_L g4182 ( 
.A(n_4085),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4122),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4132),
.Y(n_4184)
);

INVx3_ASAP7_75t_L g4185 ( 
.A(n_4120),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_4074),
.B(n_4007),
.Y(n_4186)
);

AND2x4_ASAP7_75t_L g4187 ( 
.A(n_4084),
.B(n_4140),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4112),
.Y(n_4188)
);

INVx3_ASAP7_75t_L g4189 ( 
.A(n_4064),
.Y(n_4189)
);

AOI21x1_ASAP7_75t_L g4190 ( 
.A1(n_4100),
.A2(n_3966),
.B(n_4050),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4130),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_4137),
.Y(n_4192)
);

OAI21x1_ASAP7_75t_L g4193 ( 
.A1(n_4123),
.A2(n_4033),
.B(n_4041),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4114),
.Y(n_4194)
);

OA21x2_ASAP7_75t_L g4195 ( 
.A1(n_4136),
.A2(n_3933),
.B(n_4042),
.Y(n_4195)
);

AND2x4_ASAP7_75t_L g4196 ( 
.A(n_4145),
.B(n_3997),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4071),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4071),
.Y(n_4198)
);

AND2x4_ASAP7_75t_L g4199 ( 
.A(n_4094),
.B(n_4013),
.Y(n_4199)
);

AOI21x1_ASAP7_75t_L g4200 ( 
.A1(n_4087),
.A2(n_4050),
.B(n_3967),
.Y(n_4200)
);

BUFx3_ASAP7_75t_L g4201 ( 
.A(n_4116),
.Y(n_4201)
);

INVx3_ASAP7_75t_L g4202 ( 
.A(n_4129),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4121),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4128),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4108),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4115),
.Y(n_4206)
);

CKINVDCx20_ASAP7_75t_R g4207 ( 
.A(n_4080),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4062),
.Y(n_4208)
);

INVxp67_ASAP7_75t_L g4209 ( 
.A(n_4069),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_4152),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_4062),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4149),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_4113),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4146),
.Y(n_4214)
);

INVx3_ASAP7_75t_L g4215 ( 
.A(n_4088),
.Y(n_4215)
);

NOR2xp33_ASAP7_75t_L g4216 ( 
.A(n_4159),
.B(n_4049),
.Y(n_4216)
);

AOI221xp5_ASAP7_75t_L g4217 ( 
.A1(n_4171),
.A2(n_4089),
.B1(n_4075),
.B2(n_4090),
.C(n_4046),
.Y(n_4217)
);

CKINVDCx5p33_ASAP7_75t_R g4218 ( 
.A(n_4207),
.Y(n_4218)
);

OAI22xp5_ASAP7_75t_L g4219 ( 
.A1(n_4164),
.A2(n_4073),
.B1(n_4102),
.B2(n_4103),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4188),
.Y(n_4220)
);

OAI221xp5_ASAP7_75t_L g4221 ( 
.A1(n_4195),
.A2(n_4078),
.B1(n_4134),
.B2(n_4125),
.C(n_4081),
.Y(n_4221)
);

AND2x4_ASAP7_75t_L g4222 ( 
.A(n_4182),
.B(n_4154),
.Y(n_4222)
);

BUFx2_ASAP7_75t_L g4223 ( 
.A(n_4167),
.Y(n_4223)
);

HB1xp67_ASAP7_75t_L g4224 ( 
.A(n_4169),
.Y(n_4224)
);

AOI22xp33_ASAP7_75t_L g4225 ( 
.A1(n_4165),
.A2(n_4143),
.B1(n_4067),
.B2(n_4077),
.Y(n_4225)
);

INVx2_ASAP7_75t_L g4226 ( 
.A(n_4203),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_4189),
.B(n_4076),
.Y(n_4227)
);

HB1xp67_ASAP7_75t_L g4228 ( 
.A(n_4161),
.Y(n_4228)
);

BUFx3_ASAP7_75t_L g4229 ( 
.A(n_4170),
.Y(n_4229)
);

OAI21xp5_ASAP7_75t_L g4230 ( 
.A1(n_4158),
.A2(n_3986),
.B(n_4131),
.Y(n_4230)
);

INVx2_ASAP7_75t_L g4231 ( 
.A(n_4197),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4188),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4180),
.B(n_4092),
.Y(n_4233)
);

INVx4_ASAP7_75t_L g4234 ( 
.A(n_4201),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_4156),
.A2(n_4004),
.B1(n_3998),
.B2(n_4055),
.Y(n_4235)
);

AO21x2_ASAP7_75t_L g4236 ( 
.A1(n_4205),
.A2(n_4066),
.B(n_4126),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4162),
.B(n_4098),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4163),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_4198),
.Y(n_4239)
);

OAI22xp33_ASAP7_75t_L g4240 ( 
.A1(n_4185),
.A2(n_4095),
.B1(n_4107),
.B2(n_3967),
.Y(n_4240)
);

OAI221xp5_ASAP7_75t_L g4241 ( 
.A1(n_4206),
.A2(n_3901),
.B1(n_4142),
.B2(n_3895),
.C(n_4054),
.Y(n_4241)
);

AOI21xp33_ASAP7_75t_L g4242 ( 
.A1(n_4172),
.A2(n_4110),
.B(n_4119),
.Y(n_4242)
);

NAND3xp33_ASAP7_75t_L g4243 ( 
.A(n_4208),
.B(n_3898),
.C(n_3919),
.Y(n_4243)
);

AOI22xp33_ASAP7_75t_L g4244 ( 
.A1(n_4209),
.A2(n_4118),
.B1(n_4053),
.B2(n_4009),
.Y(n_4244)
);

OR2x6_ASAP7_75t_L g4245 ( 
.A(n_4196),
.B(n_4048),
.Y(n_4245)
);

AOI22xp33_ASAP7_75t_L g4246 ( 
.A1(n_4187),
.A2(n_4053),
.B1(n_4060),
.B2(n_3980),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_4173),
.A2(n_4211),
.B(n_4193),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4163),
.Y(n_4248)
);

OAI21x1_ASAP7_75t_L g4249 ( 
.A1(n_4215),
.A2(n_4117),
.B(n_4141),
.Y(n_4249)
);

NAND3xp33_ASAP7_75t_L g4250 ( 
.A(n_4211),
.B(n_4096),
.C(n_3994),
.Y(n_4250)
);

AOI221xp5_ASAP7_75t_L g4251 ( 
.A1(n_4204),
.A2(n_4039),
.B1(n_3999),
.B2(n_4056),
.C(n_4051),
.Y(n_4251)
);

AOI221xp5_ASAP7_75t_L g4252 ( 
.A1(n_4194),
.A2(n_3991),
.B1(n_3992),
.B2(n_4020),
.C(n_4030),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_4186),
.Y(n_4253)
);

OR2x2_ASAP7_75t_L g4254 ( 
.A(n_4191),
.B(n_4148),
.Y(n_4254)
);

CKINVDCx14_ASAP7_75t_R g4255 ( 
.A(n_4160),
.Y(n_4255)
);

NAND3xp33_ASAP7_75t_L g4256 ( 
.A(n_4210),
.B(n_4044),
.C(n_3987),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4155),
.B(n_4148),
.Y(n_4257)
);

AOI22xp33_ASAP7_75t_L g4258 ( 
.A1(n_4199),
.A2(n_4135),
.B1(n_4133),
.B2(n_3917),
.Y(n_4258)
);

OAI33xp33_ASAP7_75t_L g4259 ( 
.A1(n_4176),
.A2(n_3992),
.A3(n_4030),
.B1(n_4144),
.B2(n_66),
.B3(n_68),
.Y(n_4259)
);

AO31x2_ASAP7_75t_L g4260 ( 
.A1(n_4212),
.A2(n_3893),
.A3(n_3927),
.B(n_4138),
.Y(n_4260)
);

BUFx2_ASAP7_75t_L g4261 ( 
.A(n_4196),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4183),
.Y(n_4262)
);

OR2x2_ASAP7_75t_L g4263 ( 
.A(n_4192),
.B(n_3947),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4157),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4183),
.Y(n_4265)
);

OAI22xp33_ASAP7_75t_L g4266 ( 
.A1(n_4200),
.A2(n_4038),
.B1(n_4037),
.B2(n_4025),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4224),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4220),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_4261),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4232),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4228),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4257),
.B(n_4184),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4226),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4238),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4233),
.B(n_4202),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4248),
.Y(n_4276)
);

INVxp67_ASAP7_75t_L g4277 ( 
.A(n_4229),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4231),
.Y(n_4278)
);

NAND2x1_ASAP7_75t_SL g4279 ( 
.A(n_4234),
.B(n_4200),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4239),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4262),
.Y(n_4281)
);

NOR2xp67_ASAP7_75t_L g4282 ( 
.A(n_4219),
.B(n_4213),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_4264),
.Y(n_4283)
);

HB1xp67_ASAP7_75t_L g4284 ( 
.A(n_4255),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_4223),
.B(n_4214),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_SL g4286 ( 
.A(n_4225),
.B(n_4181),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4265),
.B(n_4168),
.Y(n_4287)
);

BUFx3_ASAP7_75t_L g4288 ( 
.A(n_4218),
.Y(n_4288)
);

OR2x2_ASAP7_75t_L g4289 ( 
.A(n_4254),
.B(n_4177),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_4236),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_4263),
.B(n_4166),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4237),
.Y(n_4292)
);

AOI22xp5_ASAP7_75t_L g4293 ( 
.A1(n_4217),
.A2(n_4175),
.B1(n_4178),
.B2(n_4174),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4227),
.Y(n_4294)
);

INVx4_ASAP7_75t_L g4295 ( 
.A(n_4245),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4243),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4244),
.B(n_4179),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4247),
.Y(n_4298)
);

BUFx2_ASAP7_75t_L g4299 ( 
.A(n_4253),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4249),
.Y(n_4300)
);

AOI22xp33_ASAP7_75t_L g4301 ( 
.A1(n_4221),
.A2(n_4014),
.B1(n_3949),
.B2(n_4015),
.Y(n_4301)
);

INVxp67_ASAP7_75t_SL g4302 ( 
.A(n_4230),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4222),
.B(n_4190),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4256),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4287),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4291),
.Y(n_4306)
);

HB1xp67_ASAP7_75t_L g4307 ( 
.A(n_4284),
.Y(n_4307)
);

BUFx3_ASAP7_75t_L g4308 ( 
.A(n_4288),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4287),
.Y(n_4309)
);

AND2x4_ASAP7_75t_L g4310 ( 
.A(n_4295),
.B(n_4258),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4293),
.B(n_4302),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4293),
.B(n_4251),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4289),
.Y(n_4313)
);

AND2x2_ASAP7_75t_L g4314 ( 
.A(n_4295),
.B(n_4242),
.Y(n_4314)
);

HB1xp67_ASAP7_75t_L g4315 ( 
.A(n_4267),
.Y(n_4315)
);

NOR2xp67_ASAP7_75t_L g4316 ( 
.A(n_4282),
.B(n_4298),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_4273),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4304),
.B(n_4252),
.Y(n_4318)
);

AOI221x1_ASAP7_75t_SL g4319 ( 
.A1(n_4296),
.A2(n_4216),
.B1(n_4235),
.B2(n_4240),
.C(n_4266),
.Y(n_4319)
);

AND2x2_ASAP7_75t_L g4320 ( 
.A(n_4275),
.B(n_4246),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4271),
.B(n_4297),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4268),
.Y(n_4322)
);

AND2x4_ASAP7_75t_L g4323 ( 
.A(n_4277),
.B(n_4250),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4278),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_4269),
.B(n_4292),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4270),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4274),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4280),
.Y(n_4328)
);

INVx1_ASAP7_75t_SL g4329 ( 
.A(n_4299),
.Y(n_4329)
);

OR2x2_ASAP7_75t_L g4330 ( 
.A(n_4272),
.B(n_4260),
.Y(n_4330)
);

INVx2_ASAP7_75t_L g4331 ( 
.A(n_4283),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4276),
.Y(n_4332)
);

OR2x2_ASAP7_75t_L g4333 ( 
.A(n_4272),
.B(n_4241),
.Y(n_4333)
);

AND2x4_ASAP7_75t_L g4334 ( 
.A(n_4285),
.B(n_3913),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4281),
.Y(n_4335)
);

NAND2x1_ASAP7_75t_SL g4336 ( 
.A(n_4303),
.B(n_4259),
.Y(n_4336)
);

OR2x2_ASAP7_75t_L g4337 ( 
.A(n_4286),
.B(n_4294),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4290),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4300),
.B(n_3958),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4279),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4307),
.B(n_4301),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_4329),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4315),
.Y(n_4343)
);

AND2x4_ASAP7_75t_L g4344 ( 
.A(n_4308),
.B(n_4059),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4335),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_4319),
.B(n_4058),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4325),
.Y(n_4347)
);

INVx3_ASAP7_75t_L g4348 ( 
.A(n_4310),
.Y(n_4348)
);

OR2x2_ASAP7_75t_SL g4349 ( 
.A(n_4318),
.B(n_4023),
.Y(n_4349)
);

NAND2x1_ASAP7_75t_L g4350 ( 
.A(n_4316),
.B(n_4323),
.Y(n_4350)
);

OR2x2_ASAP7_75t_L g4351 ( 
.A(n_4333),
.B(n_64),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4305),
.Y(n_4352)
);

INVx4_ASAP7_75t_L g4353 ( 
.A(n_4323),
.Y(n_4353)
);

NOR2xp67_ASAP7_75t_L g4354 ( 
.A(n_4340),
.B(n_64),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4313),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4322),
.Y(n_4356)
);

OAI221xp5_ASAP7_75t_L g4357 ( 
.A1(n_4336),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.C(n_69),
.Y(n_4357)
);

OAI322xp33_ASAP7_75t_SL g4358 ( 
.A1(n_4311),
.A2(n_1073),
.A3(n_1072),
.B1(n_1070),
.B2(n_1069),
.C1(n_1068),
.C2(n_1067),
.Y(n_4358)
);

OAI22xp5_ASAP7_75t_SL g4359 ( 
.A1(n_4312),
.A2(n_4031),
.B1(n_4028),
.B2(n_4052),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4326),
.Y(n_4360)
);

OR2x2_ASAP7_75t_L g4361 ( 
.A(n_4321),
.B(n_66),
.Y(n_4361)
);

HB1xp67_ASAP7_75t_L g4362 ( 
.A(n_4339),
.Y(n_4362)
);

INVx1_ASAP7_75t_SL g4363 ( 
.A(n_4314),
.Y(n_4363)
);

NAND2x1p5_ASAP7_75t_L g4364 ( 
.A(n_4354),
.B(n_4340),
.Y(n_4364)
);

BUFx2_ASAP7_75t_L g4365 ( 
.A(n_4353),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4342),
.B(n_4309),
.Y(n_4366)
);

AND2x4_ASAP7_75t_L g4367 ( 
.A(n_4343),
.B(n_4353),
.Y(n_4367)
);

OR2x2_ASAP7_75t_L g4368 ( 
.A(n_4351),
.B(n_4337),
.Y(n_4368)
);

INVxp67_ASAP7_75t_SL g4369 ( 
.A(n_4361),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4355),
.Y(n_4370)
);

AND2x2_ASAP7_75t_L g4371 ( 
.A(n_4348),
.B(n_4320),
.Y(n_4371)
);

INVx3_ASAP7_75t_L g4372 ( 
.A(n_4350),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4352),
.B(n_4327),
.Y(n_4373)
);

NAND4xp25_ASAP7_75t_SL g4374 ( 
.A(n_4363),
.B(n_4357),
.C(n_4346),
.D(n_4341),
.Y(n_4374)
);

INVx1_ASAP7_75t_SL g4375 ( 
.A(n_4344),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4347),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4362),
.B(n_4306),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_4356),
.B(n_4332),
.Y(n_4378)
);

BUFx2_ASAP7_75t_L g4379 ( 
.A(n_4349),
.Y(n_4379)
);

INVx1_ASAP7_75t_SL g4380 ( 
.A(n_4365),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_4371),
.B(n_4360),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4366),
.Y(n_4382)
);

AND2x2_ASAP7_75t_L g4383 ( 
.A(n_4367),
.B(n_4345),
.Y(n_4383)
);

OR2x2_ASAP7_75t_L g4384 ( 
.A(n_4370),
.B(n_4330),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4367),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_4377),
.B(n_4317),
.Y(n_4386)
);

INVx1_ASAP7_75t_SL g4387 ( 
.A(n_4372),
.Y(n_4387)
);

OR2x2_ASAP7_75t_L g4388 ( 
.A(n_4369),
.B(n_4324),
.Y(n_4388)
);

NAND2x1p5_ASAP7_75t_L g4389 ( 
.A(n_4372),
.B(n_4358),
.Y(n_4389)
);

OR2x2_ASAP7_75t_L g4390 ( 
.A(n_4368),
.B(n_4328),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4376),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4378),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4364),
.B(n_4331),
.Y(n_4393)
);

AOI221xp5_ASAP7_75t_L g4394 ( 
.A1(n_4374),
.A2(n_4359),
.B1(n_4338),
.B2(n_4334),
.C(n_69),
.Y(n_4394)
);

OR2x2_ASAP7_75t_L g4395 ( 
.A(n_4375),
.B(n_68),
.Y(n_4395)
);

OR2x2_ASAP7_75t_L g4396 ( 
.A(n_4375),
.B(n_70),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4373),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4379),
.B(n_70),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_SL g4399 ( 
.A1(n_4380),
.A2(n_4387),
.B1(n_4385),
.B2(n_4389),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4396),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4388),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4390),
.Y(n_4402)
);

OR2x2_ASAP7_75t_L g4403 ( 
.A(n_4398),
.B(n_72),
.Y(n_4403)
);

AOI22xp33_ASAP7_75t_L g4404 ( 
.A1(n_4393),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_4404)
);

AND2x2_ASAP7_75t_L g4405 ( 
.A(n_4386),
.B(n_74),
.Y(n_4405)
);

HB1xp67_ASAP7_75t_L g4406 ( 
.A(n_4391),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4384),
.Y(n_4407)
);

AOI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_4381),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_4408)
);

INVxp33_ASAP7_75t_L g4409 ( 
.A(n_4383),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4382),
.Y(n_4410)
);

OR2x2_ASAP7_75t_L g4411 ( 
.A(n_4392),
.B(n_76),
.Y(n_4411)
);

OAI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_4397),
.A2(n_77),
.B(n_78),
.Y(n_4412)
);

O2A1O1Ixp33_ASAP7_75t_L g4413 ( 
.A1(n_4380),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_4413)
);

INVxp67_ASAP7_75t_SL g4414 ( 
.A(n_4395),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4395),
.Y(n_4415)
);

NAND4xp25_ASAP7_75t_L g4416 ( 
.A(n_4394),
.B(n_83),
.C(n_81),
.D(n_82),
.Y(n_4416)
);

AOI22xp5_ASAP7_75t_L g4417 ( 
.A1(n_4380),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_L g4418 ( 
.A(n_4405),
.B(n_82),
.Y(n_4418)
);

OAI221xp5_ASAP7_75t_L g4419 ( 
.A1(n_4399),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.C(n_86),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_SL g4420 ( 
.A1(n_4401),
.A2(n_4402),
.B1(n_4414),
.B2(n_4407),
.Y(n_4420)
);

AND2x2_ASAP7_75t_L g4421 ( 
.A(n_4409),
.B(n_85),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4404),
.B(n_86),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4406),
.Y(n_4423)
);

OR2x2_ASAP7_75t_L g4424 ( 
.A(n_4411),
.B(n_89),
.Y(n_4424)
);

OR2x2_ASAP7_75t_L g4425 ( 
.A(n_4403),
.B(n_89),
.Y(n_4425)
);

AND2x4_ASAP7_75t_L g4426 ( 
.A(n_4400),
.B(n_90),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4417),
.Y(n_4427)
);

AOI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4413),
.A2(n_91),
.B(n_93),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4415),
.B(n_4408),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_4412),
.B(n_93),
.Y(n_4430)
);

OAI21xp33_ASAP7_75t_L g4431 ( 
.A1(n_4410),
.A2(n_95),
.B(n_96),
.Y(n_4431)
);

OAI211xp5_ASAP7_75t_L g4432 ( 
.A1(n_4399),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_4432)
);

OAI22xp33_ASAP7_75t_L g4433 ( 
.A1(n_4416),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4405),
.B(n_100),
.Y(n_4434)
);

OAI22xp5_ASAP7_75t_L g4435 ( 
.A1(n_4399),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_4416),
.B(n_102),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4405),
.B(n_103),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4405),
.B(n_103),
.Y(n_4438)
);

OAI221xp5_ASAP7_75t_L g4439 ( 
.A1(n_4399),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.C(n_107),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4406),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_4406),
.Y(n_4441)
);

AOI21xp5_ASAP7_75t_L g4442 ( 
.A1(n_4435),
.A2(n_107),
.B(n_108),
.Y(n_4442)
);

AOI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_4432),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_4443)
);

O2A1O1Ixp33_ASAP7_75t_L g4444 ( 
.A1(n_4419),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4437),
.B(n_111),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_SL g4446 ( 
.A(n_4433),
.B(n_111),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4421),
.Y(n_4447)
);

OAI221xp5_ASAP7_75t_L g4448 ( 
.A1(n_4439),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.C(n_117),
.Y(n_4448)
);

AOI322xp5_ASAP7_75t_L g4449 ( 
.A1(n_4427),
.A2(n_113),
.A3(n_114),
.B1(n_116),
.B2(n_118),
.C1(n_119),
.C2(n_120),
.Y(n_4449)
);

OR2x2_ASAP7_75t_L g4450 ( 
.A(n_4424),
.B(n_116),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4425),
.Y(n_4451)
);

AOI221xp5_ASAP7_75t_L g4452 ( 
.A1(n_4423),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.C(n_123),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4440),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4436),
.B(n_120),
.Y(n_4454)
);

OAI21xp33_ASAP7_75t_L g4455 ( 
.A1(n_4420),
.A2(n_121),
.B(n_122),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4441),
.Y(n_4456)
);

AOI21xp5_ASAP7_75t_L g4457 ( 
.A1(n_4428),
.A2(n_121),
.B(n_122),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4426),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4426),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4418),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_4430),
.B(n_123),
.Y(n_4461)
);

INVx1_ASAP7_75t_SL g4462 ( 
.A(n_4434),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4438),
.Y(n_4463)
);

INVxp67_ASAP7_75t_SL g4464 ( 
.A(n_4422),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4431),
.Y(n_4465)
);

NOR3xp33_ASAP7_75t_L g4466 ( 
.A(n_4446),
.B(n_4429),
.C(n_124),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4450),
.Y(n_4467)
);

AOI211xp5_ASAP7_75t_L g4468 ( 
.A1(n_4448),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_4468)
);

AOI222xp33_ASAP7_75t_L g4469 ( 
.A1(n_4465),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.C1(n_129),
.C2(n_130),
.Y(n_4469)
);

NOR2xp67_ASAP7_75t_SL g4470 ( 
.A(n_4453),
.B(n_4456),
.Y(n_4470)
);

AOI221xp5_ASAP7_75t_L g4471 ( 
.A1(n_4444),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.C(n_129),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4449),
.B(n_126),
.Y(n_4472)
);

NAND3xp33_ASAP7_75t_L g4473 ( 
.A(n_4452),
.B(n_129),
.C(n_130),
.Y(n_4473)
);

OAI221xp5_ASAP7_75t_L g4474 ( 
.A1(n_4443),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_135),
.Y(n_4474)
);

AOI221xp5_ASAP7_75t_L g4475 ( 
.A1(n_4457),
.A2(n_135),
.B1(n_132),
.B2(n_134),
.C(n_136),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4445),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_SL g4477 ( 
.A(n_4443),
.B(n_135),
.Y(n_4477)
);

INVx1_ASAP7_75t_SL g4478 ( 
.A(n_4458),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4459),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4454),
.B(n_137),
.Y(n_4480)
);

AOI222xp33_ASAP7_75t_L g4481 ( 
.A1(n_4447),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.C1(n_142),
.C2(n_143),
.Y(n_4481)
);

AOI221xp5_ASAP7_75t_L g4482 ( 
.A1(n_4442),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.C(n_142),
.Y(n_4482)
);

OAI21xp5_ASAP7_75t_SL g4483 ( 
.A1(n_4462),
.A2(n_4451),
.B(n_4460),
.Y(n_4483)
);

AOI22xp5_ASAP7_75t_L g4484 ( 
.A1(n_4464),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_4484)
);

AOI211x1_ASAP7_75t_L g4485 ( 
.A1(n_4463),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_4485)
);

AOI211xp5_ASAP7_75t_SL g4486 ( 
.A1(n_4455),
.A2(n_150),
.B(n_147),
.C(n_148),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4461),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4480),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_4477),
.Y(n_4489)
);

OAI32xp33_ASAP7_75t_L g4490 ( 
.A1(n_4478),
.A2(n_152),
.A3(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_4479),
.Y(n_4491)
);

INVxp67_ASAP7_75t_L g4492 ( 
.A(n_4470),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4469),
.B(n_158),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_4486),
.B(n_160),
.Y(n_4494)
);

OAI221xp5_ASAP7_75t_L g4495 ( 
.A1(n_4471),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.C(n_163),
.Y(n_4495)
);

OAI221xp5_ASAP7_75t_L g4496 ( 
.A1(n_4482),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.C(n_163),
.Y(n_4496)
);

OAI211xp5_ASAP7_75t_L g4497 ( 
.A1(n_4468),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4484),
.Y(n_4498)
);

INVxp33_ASAP7_75t_L g4499 ( 
.A(n_4466),
.Y(n_4499)
);

OAI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4472),
.A2(n_164),
.B1(n_161),
.B2(n_162),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4485),
.Y(n_4501)
);

OR2x2_ASAP7_75t_L g4502 ( 
.A(n_4476),
.B(n_166),
.Y(n_4502)
);

OAI22xp33_ASAP7_75t_L g4503 ( 
.A1(n_4473),
.A2(n_4474),
.B1(n_4467),
.B2(n_4483),
.Y(n_4503)
);

OAI211xp5_ASAP7_75t_L g4504 ( 
.A1(n_4481),
.A2(n_170),
.B(n_167),
.C(n_169),
.Y(n_4504)
);

AOI211xp5_ASAP7_75t_L g4505 ( 
.A1(n_4475),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4487),
.Y(n_4506)
);

AOI21xp33_ASAP7_75t_SL g4507 ( 
.A1(n_4503),
.A2(n_171),
.B(n_172),
.Y(n_4507)
);

AOI211xp5_ASAP7_75t_SL g4508 ( 
.A1(n_4497),
.A2(n_174),
.B(n_171),
.C(n_173),
.Y(n_4508)
);

AOI22xp5_ASAP7_75t_L g4509 ( 
.A1(n_4492),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_4509)
);

AOI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_4500),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_4510)
);

AOI221xp5_ASAP7_75t_L g4511 ( 
.A1(n_4490),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.C(n_179),
.Y(n_4511)
);

OAI22xp5_ASAP7_75t_L g4512 ( 
.A1(n_4494),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_4512)
);

INVx1_ASAP7_75t_SL g4513 ( 
.A(n_4491),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4489),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4502),
.Y(n_4515)
);

OAI22xp5_ASAP7_75t_L g4516 ( 
.A1(n_4493),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4501),
.B(n_180),
.Y(n_4517)
);

OAI22xp33_ASAP7_75t_L g4518 ( 
.A1(n_4499),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4498),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4495),
.Y(n_4520)
);

AOI22xp5_ASAP7_75t_L g4521 ( 
.A1(n_4504),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_4521)
);

AO221x1_ASAP7_75t_L g4522 ( 
.A1(n_4488),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.C(n_188),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4496),
.Y(n_4523)
);

AOI22xp5_ASAP7_75t_L g4524 ( 
.A1(n_4506),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_4524)
);

AND2x4_ASAP7_75t_L g4525 ( 
.A(n_4514),
.B(n_4505),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4522),
.Y(n_4526)
);

AOI221x1_ASAP7_75t_L g4527 ( 
.A1(n_4507),
.A2(n_4519),
.B1(n_4516),
.B2(n_4512),
.C(n_4520),
.Y(n_4527)
);

NAND3xp33_ASAP7_75t_L g4528 ( 
.A(n_4511),
.B(n_189),
.C(n_190),
.Y(n_4528)
);

OAI211xp5_ASAP7_75t_L g4529 ( 
.A1(n_4521),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_4529)
);

OAI22xp33_ASAP7_75t_SL g4530 ( 
.A1(n_4517),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_4530)
);

NAND3xp33_ASAP7_75t_SL g4531 ( 
.A(n_4513),
.B(n_192),
.C(n_193),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4509),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4508),
.B(n_193),
.Y(n_4533)
);

OR3x1_ASAP7_75t_L g4534 ( 
.A(n_4523),
.B(n_194),
.C(n_195),
.Y(n_4534)
);

OA22x2_ASAP7_75t_SL g4535 ( 
.A1(n_4515),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_4535)
);

AOI21xp5_ASAP7_75t_L g4536 ( 
.A1(n_4518),
.A2(n_198),
.B(n_199),
.Y(n_4536)
);

NOR2x1_ASAP7_75t_L g4537 ( 
.A(n_4534),
.B(n_4524),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4526),
.Y(n_4538)
);

NOR2x1_ASAP7_75t_L g4539 ( 
.A(n_4528),
.B(n_4510),
.Y(n_4539)
);

NOR2x1_ASAP7_75t_L g4540 ( 
.A(n_4533),
.B(n_199),
.Y(n_4540)
);

AO22x1_ASAP7_75t_L g4541 ( 
.A1(n_4525),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_4541)
);

NOR2x1_ASAP7_75t_L g4542 ( 
.A(n_4531),
.B(n_200),
.Y(n_4542)
);

AOI221xp5_ASAP7_75t_L g4543 ( 
.A1(n_4530),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_4543)
);

OR2x2_ASAP7_75t_L g4544 ( 
.A(n_4532),
.B(n_205),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4536),
.B(n_205),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4535),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4529),
.Y(n_4547)
);

NOR2x1p5_ASAP7_75t_L g4548 ( 
.A(n_4538),
.B(n_4527),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4544),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4542),
.Y(n_4550)
);

NAND4xp75_ASAP7_75t_L g4551 ( 
.A(n_4540),
.B(n_205),
.C(n_206),
.D(n_207),
.Y(n_4551)
);

XOR2x2_ASAP7_75t_L g4552 ( 
.A(n_4537),
.B(n_206),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_4546),
.B(n_4547),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4545),
.Y(n_4554)
);

XNOR2xp5_ASAP7_75t_L g4555 ( 
.A(n_4539),
.B(n_208),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4541),
.B(n_208),
.Y(n_4556)
);

NAND3xp33_ASAP7_75t_L g4557 ( 
.A(n_4543),
.B(n_208),
.C(n_209),
.Y(n_4557)
);

AOI32xp33_ASAP7_75t_L g4558 ( 
.A1(n_4553),
.A2(n_210),
.A3(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_4558)
);

AOI221xp5_ASAP7_75t_L g4559 ( 
.A1(n_4556),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.C(n_213),
.Y(n_4559)
);

AOI22xp5_ASAP7_75t_L g4560 ( 
.A1(n_4548),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_4560)
);

AOI211xp5_ASAP7_75t_L g4561 ( 
.A1(n_4557),
.A2(n_214),
.B(n_215),
.C(n_216),
.Y(n_4561)
);

AOI22xp5_ASAP7_75t_L g4562 ( 
.A1(n_4555),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_4562)
);

OR5x1_ASAP7_75t_L g4563 ( 
.A(n_4552),
.B(n_217),
.C(n_218),
.D(n_219),
.E(n_220),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4562),
.B(n_4549),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4563),
.Y(n_4565)
);

XNOR2x1_ASAP7_75t_L g4566 ( 
.A(n_4560),
.B(n_4551),
.Y(n_4566)
);

AND2x2_ASAP7_75t_SL g4567 ( 
.A(n_4559),
.B(n_4554),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4558),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4561),
.Y(n_4569)
);

NOR2xp33_ASAP7_75t_L g4570 ( 
.A(n_4568),
.B(n_4550),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4565),
.Y(n_4571)
);

BUFx3_ASAP7_75t_L g4572 ( 
.A(n_4564),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4567),
.Y(n_4573)
);

INVx3_ASAP7_75t_L g4574 ( 
.A(n_4566),
.Y(n_4574)
);

AOI22xp5_ASAP7_75t_L g4575 ( 
.A1(n_4569),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_4575)
);

NOR2x1_ASAP7_75t_L g4576 ( 
.A(n_4572),
.B(n_4573),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_4576),
.Y(n_4577)
);

CKINVDCx20_ASAP7_75t_R g4578 ( 
.A(n_4577),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4577),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_4578),
.A2(n_4570),
.B1(n_4571),
.B2(n_4574),
.Y(n_4580)
);

INVx2_ASAP7_75t_L g4581 ( 
.A(n_4579),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4581),
.Y(n_4582)
);

AOI22xp5_ASAP7_75t_L g4583 ( 
.A1(n_4580),
.A2(n_4575),
.B1(n_222),
.B2(n_223),
.Y(n_4583)
);

OAI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_4582),
.A2(n_221),
.B(n_222),
.Y(n_4584)
);

OAI22xp5_ASAP7_75t_SL g4585 ( 
.A1(n_4583),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_4585)
);

AOI222xp33_ASAP7_75t_SL g4586 ( 
.A1(n_4582),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.C1(n_228),
.C2(n_229),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4582),
.Y(n_4587)
);

AOI22xp5_ASAP7_75t_L g4588 ( 
.A1(n_4587),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_4588)
);

AOI22xp5_ASAP7_75t_SL g4589 ( 
.A1(n_4584),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_4589)
);

AOI22xp5_ASAP7_75t_L g4590 ( 
.A1(n_4586),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_4590)
);

OR2x2_ASAP7_75t_L g4591 ( 
.A(n_4588),
.B(n_4585),
.Y(n_4591)
);

OR2x6_ASAP7_75t_L g4592 ( 
.A(n_4590),
.B(n_1032),
.Y(n_4592)
);

AOI22x1_ASAP7_75t_L g4593 ( 
.A1(n_4589),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_4593)
);

AOI21xp5_ASAP7_75t_L g4594 ( 
.A1(n_4591),
.A2(n_230),
.B(n_231),
.Y(n_4594)
);

AOI211xp5_ASAP7_75t_L g4595 ( 
.A1(n_4594),
.A2(n_4592),
.B(n_4593),
.C(n_232),
.Y(n_4595)
);


endmodule