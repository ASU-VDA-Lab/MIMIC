module fake_jpeg_2756_n_185 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_24),
.Y(n_58)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_3),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_58),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_31),
.B1(n_19),
.B2(n_25),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_35),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_69),
.B1(n_76),
.B2(n_3),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_24),
.B1(n_17),
.B2(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_40),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_38),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_91),
.B1(n_94),
.B2(n_66),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_38),
.B1(n_40),
.B2(n_5),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_40),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_65),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_73),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_69),
.C(n_68),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_116),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_69),
.CI(n_76),
.CON(n_103),
.SN(n_103)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_112),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_97),
.A3(n_86),
.B1(n_69),
.B2(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_77),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_65),
.C(n_61),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_75),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_71),
.B(n_73),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_88),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_98),
.B1(n_89),
.B2(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_129),
.B1(n_134),
.B2(n_137),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_98),
.B1(n_80),
.B2(n_93),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_73),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_135),
.C(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_52),
.B1(n_101),
.B2(n_8),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_6),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_52),
.B1(n_7),
.B2(n_8),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_103),
.B1(n_117),
.B2(n_111),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_106),
.B(n_120),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_145),
.B(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_148),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_119),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_109),
.B1(n_115),
.B2(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_104),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_122),
.B1(n_127),
.B2(n_129),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_126),
.C(n_130),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_161),
.C(n_146),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_136),
.B(n_138),
.C(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_160),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_142),
.B1(n_140),
.B2(n_147),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_122),
.CI(n_113),
.CON(n_155),
.SN(n_155)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_105),
.B(n_108),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_105),
.A3(n_113),
.B1(n_104),
.B2(n_108),
.C1(n_7),
.C2(n_12),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_113),
.C(n_105),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_150),
.B1(n_143),
.B2(n_139),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_164),
.B1(n_168),
.B2(n_153),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_105),
.C(n_108),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_159),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_168)
);

OAI31xp33_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_170),
.A3(n_172),
.B(n_159),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_158),
.B(n_161),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_158),
.B(n_153),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_159),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_159),
.B1(n_167),
.B2(n_160),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_177),
.B1(n_155),
.B2(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_175),
.B(n_176),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_156),
.C(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_180),
.B(n_10),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_179),
.B(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_180),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_13),
.Y(n_185)
);


endmodule