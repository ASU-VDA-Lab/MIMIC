module fake_jpeg_27206_n_80 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_35),
.B1(n_29),
.B2(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_3),
.B(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_35),
.B1(n_30),
.B2(n_34),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_50),
.B(n_5),
.C(n_7),
.Y(n_64)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

OR2x2_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_57),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_15),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_60),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_16),
.A3(n_23),
.B1(n_22),
.B2(n_6),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_3),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_71),
.B1(n_68),
.B2(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_75),
.B(n_64),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_59),
.B(n_65),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_69),
.B1(n_72),
.B2(n_58),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_72),
.C(n_63),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_18),
.C2(n_19),
.Y(n_80)
);


endmodule