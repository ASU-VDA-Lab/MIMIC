module fake_aes_10633_n_803 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_191, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_803);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_803;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_698;
wire n_555;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g200 ( .A(n_120), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_28), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_181), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_153), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_143), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_95), .Y(n_205) );
INVx1_ASAP7_75t_SL g206 ( .A(n_150), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_59), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_32), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_82), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_97), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_13), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_115), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_8), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_84), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_27), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_58), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_190), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_85), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_112), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
BUFx10_ASAP7_75t_L g223 ( .A(n_16), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_121), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_99), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_68), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_47), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_90), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_173), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_137), .Y(n_230) );
CKINVDCx14_ASAP7_75t_R g231 ( .A(n_45), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_91), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_21), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_134), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_74), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_140), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_4), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_177), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_179), .Y(n_239) );
BUFx5_ASAP7_75t_L g240 ( .A(n_193), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_25), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_101), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_88), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_40), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_160), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_39), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_77), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_98), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_135), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_118), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_20), .Y(n_251) );
CKINVDCx14_ASAP7_75t_R g252 ( .A(n_195), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_96), .Y(n_253) );
NOR2xp67_ASAP7_75t_L g254 ( .A(n_2), .B(n_5), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_119), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_81), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_0), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_162), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_107), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_125), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_130), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_185), .Y(n_262) );
NOR2xp67_ASAP7_75t_L g263 ( .A(n_171), .B(n_42), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_53), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_172), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_111), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_198), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_22), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_41), .Y(n_269) );
INVx2_ASAP7_75t_SL g270 ( .A(n_133), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_75), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_67), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_164), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_16), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_127), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_102), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_155), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_65), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_106), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_136), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_78), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_188), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_69), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_167), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_138), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_174), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_83), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_182), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_12), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_100), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_76), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_31), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_49), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_129), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_176), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_54), .Y(n_296) );
CKINVDCx14_ASAP7_75t_R g297 ( .A(n_180), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_8), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_5), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_165), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_29), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_80), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_240), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_284), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_209), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_249), .B(n_0), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_209), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_251), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_240), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_204), .B(n_1), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_223), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_270), .B(n_1), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_240), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_240), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_211), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_214), .B(n_3), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_218), .A2(n_24), .B(n_23), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_213), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_237), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_265), .B(n_4), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_229), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_209), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_257), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_289), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_309), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_311), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_311), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_311), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_314), .B(n_238), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_305), .B(n_265), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_314), .B(n_245), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_304), .B(n_203), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_314), .B(n_254), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_303), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_313), .B(n_327), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_312), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_313), .B(n_298), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_307), .B(n_231), .Y(n_343) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_322), .B(n_200), .Y(n_344) );
AND3x2_ASAP7_75t_L g345 ( .A(n_322), .B(n_299), .C(n_205), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_317), .A2(n_262), .B1(n_272), .B2(n_202), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_312), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_320), .B(n_206), .Y(n_350) );
INVx8_ASAP7_75t_L g351 ( .A(n_336), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_335), .B(n_321), .Y(n_352) );
BUFx5_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_SL g354 ( .A1(n_333), .A2(n_297), .B(n_252), .C(n_325), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_338), .B(n_326), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_328), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_350), .B(n_223), .Y(n_359) );
INVx4_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_343), .B(n_318), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_341), .A2(n_319), .B(n_316), .Y(n_362) );
INVxp67_ASAP7_75t_R g363 ( .A(n_346), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_331), .Y(n_364) );
OA22x2_ASAP7_75t_L g365 ( .A1(n_345), .A2(n_323), .B1(n_319), .B2(n_316), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_330), .Y(n_366) );
OAI22xp33_ASAP7_75t_L g367 ( .A1(n_342), .A2(n_292), .B1(n_293), .B2(n_286), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_336), .B(n_323), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_336), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_332), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_332), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_344), .B(n_206), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_334), .B(n_219), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_334), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_366), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g378 ( .A1(n_352), .A2(n_344), .B(n_348), .C(n_349), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_361), .B(n_348), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_356), .B(n_348), .Y(n_380) );
OAI21xp33_ASAP7_75t_L g381 ( .A1(n_359), .A2(n_340), .B(n_339), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_362), .A2(n_355), .B(n_358), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_364), .A2(n_208), .B(n_207), .Y(n_383) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_357), .B(n_26), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_371), .A2(n_215), .B(n_212), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_374), .A2(n_220), .B1(n_221), .B2(n_217), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_374), .B(n_219), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_357), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_351), .B(n_247), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_373), .A2(n_224), .B(n_222), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_376), .A2(n_226), .B(n_225), .Y(n_391) );
NOR2x1_ASAP7_75t_R g392 ( .A(n_367), .B(n_216), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_369), .B(n_247), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_375), .A2(n_264), .B1(n_244), .B2(n_246), .Y(n_394) );
INVx5_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
OA22x2_ASAP7_75t_L g396 ( .A1(n_363), .A2(n_232), .B1(n_233), .B2(n_234), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_365), .A2(n_235), .B(n_227), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_360), .B(n_253), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_353), .B(n_236), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_372), .A2(n_258), .B(n_255), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_395), .B(n_360), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_377), .B(n_368), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_382), .A2(n_354), .B(n_370), .Y(n_403) );
OAI22x1_ASAP7_75t_L g404 ( .A1(n_392), .A2(n_280), .B1(n_273), .B2(n_268), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_378), .B(n_370), .C(n_271), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_379), .A2(n_353), .B1(n_277), .B2(n_248), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_395), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_399), .A2(n_278), .B(n_267), .Y(n_408) );
AO31x2_ASAP7_75t_L g409 ( .A1(n_385), .A2(n_288), .A3(n_279), .B(n_281), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_386), .B(n_353), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_397), .B(n_271), .C(n_228), .Y(n_411) );
AOI221x1_ASAP7_75t_L g412 ( .A1(n_381), .A2(n_291), .B1(n_283), .B2(n_285), .C(n_290), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_396), .A2(n_353), .B1(n_294), .B2(n_295), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_389), .B(n_271), .C(n_228), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_387), .A2(n_300), .B(n_296), .Y(n_415) );
INVx3_ASAP7_75t_SL g416 ( .A(n_395), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_398), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_393), .A2(n_302), .B(n_263), .Y(n_418) );
OAI21x1_ASAP7_75t_L g419 ( .A1(n_384), .A2(n_276), .B(n_228), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_390), .A2(n_241), .B(n_239), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_398), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_383), .A2(n_243), .B(n_242), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_391), .A2(n_256), .B(n_250), .Y(n_425) );
AO21x1_ASAP7_75t_L g426 ( .A1(n_394), .A2(n_308), .B(n_306), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_380), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_395), .B(n_201), .Y(n_428) );
AO21x2_ASAP7_75t_L g429 ( .A1(n_382), .A2(n_301), .B(n_276), .Y(n_429) );
AO21x2_ASAP7_75t_L g430 ( .A1(n_382), .A2(n_301), .B(n_306), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_416), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_430), .A2(n_308), .B(n_306), .Y(n_432) );
BUFx12f_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_421), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_405), .A2(n_324), .B(n_275), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_403), .A2(n_324), .B(n_210), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_423), .A2(n_6), .B(n_7), .C(n_9), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_407), .B(n_6), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_427), .B(n_7), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_422), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_412), .A2(n_426), .B(n_418), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
OAI21x1_ASAP7_75t_L g444 ( .A1(n_408), .A2(n_33), .B(n_30), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_415), .A2(n_287), .B(n_282), .C(n_269), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_402), .B(n_9), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_407), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_409), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_411), .A2(n_266), .B(n_261), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_429), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_401), .Y(n_451) );
OAI21x1_ASAP7_75t_SL g452 ( .A1(n_413), .A2(n_10), .B(n_11), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_410), .A2(n_260), .B(n_259), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_414), .A2(n_420), .B(n_406), .C(n_401), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_428), .B(n_10), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_404), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_424), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_458) );
OAI21x1_ASAP7_75t_L g459 ( .A1(n_425), .A2(n_117), .B(n_197), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
AO31x2_ASAP7_75t_L g463 ( .A1(n_426), .A2(n_14), .A3(n_15), .B(n_17), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_404), .B(n_14), .Y(n_464) );
OAI21x1_ASAP7_75t_L g465 ( .A1(n_419), .A2(n_116), .B(n_196), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_416), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_417), .B(n_15), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_417), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_407), .Y(n_471) );
AO31x2_ASAP7_75t_L g472 ( .A1(n_426), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_423), .B(n_18), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_423), .A2(n_19), .B(n_20), .C(n_34), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_423), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_417), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_404), .B(n_38), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_433), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_461), .Y(n_481) );
CKINVDCx14_ASAP7_75t_R g482 ( .A(n_466), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_441), .B(n_43), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_462), .Y(n_484) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_436), .A2(n_44), .B(n_46), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_460), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_460), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_447), .B(n_48), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_448), .B(n_50), .Y(n_489) );
OR2x6_ASAP7_75t_L g490 ( .A(n_438), .B(n_51), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_464), .B(n_52), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_439), .B(n_55), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_471), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_446), .B(n_199), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_457), .A2(n_56), .B1(n_57), .B2(n_60), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_473), .A2(n_61), .B(n_62), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_468), .A2(n_63), .B1(n_64), .B2(n_66), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_467), .Y(n_500) );
CKINVDCx6p67_ASAP7_75t_R g501 ( .A(n_474), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_469), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_470), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_477), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_473), .B(n_70), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_456), .B(n_71), .Y(n_506) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_475), .B(n_72), .C(n_73), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_471), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_451), .B(n_79), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_460), .B(n_86), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_479), .Y(n_511) );
INVx6_ASAP7_75t_L g512 ( .A(n_478), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_475), .B(n_437), .C(n_454), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_443), .B(n_87), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_446), .Y(n_515) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_436), .A2(n_89), .B(n_92), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_438), .Y(n_517) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_455), .Y(n_518) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_450), .A2(n_93), .B(n_94), .Y(n_519) );
BUFx3_ASAP7_75t_L g520 ( .A(n_452), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_472), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_454), .A2(n_103), .B(n_104), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_468), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_444), .Y(n_525) );
INVx4_ASAP7_75t_L g526 ( .A(n_432), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_463), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_442), .B(n_105), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_458), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_437), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_459), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_445), .B(n_108), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_445), .B(n_109), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_442), .B(n_110), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_463), .B(n_113), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_463), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_453), .B(n_114), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_465), .Y(n_539) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_476), .A2(n_449), .B(n_453), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_476), .B(n_122), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_435), .B(n_123), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_432), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_435), .Y(n_544) );
INVxp67_ASAP7_75t_SL g545 ( .A(n_449), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_447), .B(n_124), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_441), .B(n_126), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_471), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_457), .B(n_128), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_440), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_440), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_441), .B(n_131), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_493), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_481), .B(n_132), .Y(n_555) );
BUFx3_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_490), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_543), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_521), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_490), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_490), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_500), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_548), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_502), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_523), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_503), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_484), .B(n_139), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_515), .B(n_141), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_511), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_480), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_548), .B(n_142), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_550), .B(n_144), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_508), .B(n_145), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_551), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_488), .B(n_148), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_546), .B(n_151), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_536), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_508), .B(n_152), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_530), .B(n_154), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_499), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_480), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_526), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_487), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_504), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_524), .B(n_491), .Y(n_586) );
NOR2xp67_ASAP7_75t_L g587 ( .A(n_513), .B(n_156), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_486), .B(n_157), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_529), .B(n_158), .Y(n_589) );
INVx2_ASAP7_75t_SL g590 ( .A(n_501), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_492), .B(n_159), .Y(n_591) );
BUFx3_ASAP7_75t_L g592 ( .A(n_487), .Y(n_592) );
AO21x2_ASAP7_75t_L g593 ( .A1(n_528), .A2(n_534), .B(n_522), .Y(n_593) );
NOR2x1_ASAP7_75t_SL g594 ( .A(n_520), .B(n_161), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_163), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_512), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_512), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_526), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_512), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_518), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_539), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_518), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_527), .B(n_166), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_486), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_506), .B(n_168), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_513), .B(n_169), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_537), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_510), .Y(n_609) );
INVx4_ASAP7_75t_R g610 ( .A(n_482), .Y(n_610) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_541), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_510), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_517), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_483), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_541), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_549), .B(n_170), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g617 ( .A1(n_522), .A2(n_175), .B1(n_178), .B2(n_183), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_483), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_494), .B(n_194), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_489), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_545), .B(n_184), .Y(n_621) );
AND2x4_ASAP7_75t_L g622 ( .A(n_509), .B(n_186), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_532), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_544), .Y(n_624) );
NOR2x1_ASAP7_75t_SL g625 ( .A(n_538), .B(n_187), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_489), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_549), .B(n_189), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_533), .B(n_191), .Y(n_628) );
NAND2x1_ASAP7_75t_L g629 ( .A(n_535), .B(n_192), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_564), .B(n_554), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_586), .B(n_545), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_553), .Y(n_632) );
NAND3x1_ASAP7_75t_L g633 ( .A(n_557), .B(n_497), .C(n_534), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_581), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_563), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_565), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_567), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_570), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_585), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_575), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_564), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_554), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_561), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_558), .Y(n_644) );
AND2x2_ASAP7_75t_SL g645 ( .A(n_615), .B(n_525), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_561), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_611), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_613), .Y(n_648) );
XOR2xp5_ASAP7_75t_L g649 ( .A(n_590), .B(n_496), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_557), .Y(n_650) );
INVx3_ASAP7_75t_L g651 ( .A(n_560), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_556), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_611), .B(n_547), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_560), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_562), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_583), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_596), .B(n_547), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_562), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_604), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_597), .B(n_552), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_599), .B(n_531), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_582), .B(n_514), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_601), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_582), .B(n_505), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_571), .B(n_505), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_618), .B(n_620), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_605), .B(n_497), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_600), .B(n_540), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_602), .B(n_540), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_626), .B(n_542), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_601), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_614), .B(n_542), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_614), .B(n_623), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_572), .B(n_516), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_572), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_623), .B(n_519), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_598), .B(n_507), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_612), .B(n_485), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_603), .B(n_507), .Y(n_679) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_559), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_584), .B(n_498), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_589), .B(n_496), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_580), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_566), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_580), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_632), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_631), .B(n_566), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_641), .B(n_593), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_630), .B(n_578), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_645), .B(n_579), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_635), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_636), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_637), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_638), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_641), .B(n_593), .Y(n_695) );
OR2x2_ASAP7_75t_L g696 ( .A(n_630), .B(n_578), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_649), .B(n_595), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_639), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_643), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_643), .Y(n_700) );
INVx2_ASAP7_75t_SL g701 ( .A(n_634), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_640), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_650), .B(n_608), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_654), .B(n_608), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g705 ( .A(n_652), .B(n_610), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_642), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_646), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_655), .B(n_609), .Y(n_708) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_680), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_659), .B(n_624), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_648), .Y(n_711) );
BUFx3_ASAP7_75t_L g712 ( .A(n_651), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_666), .B(n_624), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_673), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_658), .B(n_609), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_673), .B(n_574), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_651), .B(n_574), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_680), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_663), .Y(n_719) );
INVx3_ASAP7_75t_SL g720 ( .A(n_645), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_675), .B(n_579), .Y(n_721) );
INVxp67_ASAP7_75t_L g722 ( .A(n_656), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_662), .B(n_592), .Y(n_723) );
NAND3xp33_ASAP7_75t_SL g724 ( .A(n_682), .B(n_617), .C(n_616), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_667), .B(n_616), .C(n_587), .D(n_607), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_653), .B(n_592), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_671), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_686), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_691), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_705), .B(n_617), .C(n_656), .Y(n_730) );
NOR2xp67_ASAP7_75t_L g731 ( .A(n_701), .B(n_647), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_692), .Y(n_732) );
AND2x2_ASAP7_75t_SL g733 ( .A(n_697), .B(n_674), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_726), .B(n_647), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_693), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_694), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_723), .B(n_661), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_698), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_711), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_714), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_702), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_699), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_700), .B(n_683), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_706), .B(n_685), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_722), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_707), .B(n_672), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_713), .B(n_644), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_697), .B(n_665), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_687), .B(n_684), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_713), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_710), .Y(n_751) );
OAI21xp33_ASAP7_75t_L g752 ( .A1(n_724), .A2(n_678), .B(n_669), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_751), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_730), .A2(n_690), .B(n_724), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_750), .B(n_688), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_743), .Y(n_756) );
INVxp33_ASAP7_75t_L g757 ( .A(n_731), .Y(n_757) );
NAND5xp2_ASAP7_75t_L g758 ( .A(n_752), .B(n_576), .C(n_577), .D(n_627), .E(n_681), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_737), .B(n_720), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_743), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_747), .Y(n_761) );
OAI21xp33_ASAP7_75t_SL g762 ( .A1(n_733), .A2(n_690), .B(n_709), .Y(n_762) );
OAI322xp33_ASAP7_75t_L g763 ( .A1(n_746), .A2(n_722), .A3(n_720), .B1(n_689), .B2(n_696), .C1(n_688), .C2(n_695), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_749), .Y(n_764) );
OAI32xp33_ASAP7_75t_L g765 ( .A1(n_730), .A2(n_712), .A3(n_725), .B1(n_695), .B2(n_716), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_748), .A2(n_734), .B1(n_721), .B2(n_740), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_745), .B(n_708), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_762), .A2(n_747), .B(n_709), .Y(n_768) );
O2A1O1Ixp33_ASAP7_75t_L g769 ( .A1(n_754), .A2(n_744), .B(n_736), .C(n_729), .Y(n_769) );
OAI21xp33_ASAP7_75t_L g770 ( .A1(n_757), .A2(n_742), .B(n_735), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_756), .B(n_728), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_766), .A2(n_633), .B1(n_741), .B2(n_738), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_760), .A2(n_739), .B1(n_732), .B2(n_633), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_758), .A2(n_594), .B(n_710), .Y(n_774) );
AOI221x1_ASAP7_75t_L g775 ( .A1(n_758), .A2(n_607), .B1(n_621), .B2(n_727), .C(n_719), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_753), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_761), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_755), .B(n_718), .Y(n_778) );
AOI21xp33_ASAP7_75t_L g779 ( .A1(n_765), .A2(n_664), .B(n_670), .Y(n_779) );
AOI321xp33_ASAP7_75t_L g780 ( .A1(n_759), .A2(n_715), .A3(n_717), .B1(n_704), .B2(n_703), .C(n_657), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_763), .A2(n_625), .B(n_629), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_L g782 ( .A1(n_755), .A2(n_591), .B(n_619), .C(n_679), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_764), .B(n_668), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_769), .B(n_771), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_768), .A2(n_772), .B(n_770), .Y(n_785) );
NOR4xp25_ASAP7_75t_L g786 ( .A(n_779), .B(n_777), .C(n_782), .D(n_776), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_773), .A2(n_778), .B1(n_774), .B2(n_781), .C(n_783), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_784), .B(n_767), .Y(n_788) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_785), .B(n_622), .Y(n_789) );
NAND4xp25_ASAP7_75t_SL g790 ( .A(n_787), .B(n_775), .C(n_780), .D(n_676), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_788), .B(n_786), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_789), .B(n_767), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_790), .B(n_661), .Y(n_793) );
XNOR2x1_ASAP7_75t_L g794 ( .A(n_791), .B(n_622), .Y(n_794) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_793), .B(n_569), .C(n_621), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_794), .A2(n_792), .B1(n_628), .B2(n_606), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_795), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_797), .A2(n_569), .B(n_603), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_796), .B(n_677), .Y(n_799) );
AOI21xp33_ASAP7_75t_SL g800 ( .A1(n_799), .A2(n_798), .B(n_588), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_800), .A2(n_573), .B(n_568), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_801), .B(n_555), .Y(n_802) );
OAI21xp33_ASAP7_75t_L g803 ( .A1(n_802), .A2(n_660), .B(n_679), .Y(n_803) );
endmodule