module fake_jpeg_15531_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_36),
.B(n_39),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_1),
.Y(n_37)
);

NOR2xp67_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_30),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_48),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_74),
.B1(n_21),
.B2(n_31),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_66),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_37),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_70),
.C(n_30),
.Y(n_77)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_41),
.B(n_26),
.Y(n_73)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_35),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_77),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_96),
.B1(n_60),
.B2(n_71),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_42),
.B1(n_45),
.B2(n_18),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_27),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_19),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_89),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_31),
.B1(n_25),
.B2(n_20),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_55),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_33),
.B1(n_32),
.B2(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_83),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_88),
.B(n_93),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_120),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_49),
.C(n_50),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_118),
.C(n_106),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_98),
.B1(n_100),
.B2(n_33),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_64),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_60),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_50),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_90),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_92),
.B1(n_78),
.B2(n_99),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_132),
.Y(n_143)
);

NOR4xp25_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_82),
.C(n_79),
.D(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_82),
.C(n_100),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_101),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_134),
.C(n_139),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_107),
.B1(n_113),
.B2(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_98),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_49),
.B(n_28),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_148),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_103),
.C(n_112),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_126),
.C(n_139),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_117),
.Y(n_152)
);

XOR2x2_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_106),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_136),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_145),
.Y(n_154)
);

OAI322xp33_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_160),
.A3(n_161),
.B1(n_150),
.B2(n_125),
.C1(n_133),
.C2(n_109),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_138),
.C(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_115),
.C(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_164),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_136),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_137),
.C(n_122),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_136),
.B1(n_144),
.B2(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_167),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_150),
.B(n_151),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_171),
.B(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_151),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_158),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_149),
.A3(n_125),
.B1(n_109),
.B2(n_28),
.C1(n_97),
.C2(n_59),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_176),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_169),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

NOR2x1_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_154),
.Y(n_181)
);

AOI21x1_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_2),
.B(n_4),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_175),
.A3(n_62),
.B1(n_59),
.B2(n_15),
.C1(n_13),
.C2(n_9),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_182),
.B(n_183),
.Y(n_187)
);

AOI332xp33_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_15),
.A3(n_13),
.B1(n_6),
.B2(n_7),
.B3(n_8),
.C1(n_2),
.C2(n_10),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_185),
.A2(n_186),
.B(n_7),
.C(n_8),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_188),
.B(n_7),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_190)
);


endmodule