module fake_jpeg_19517_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_27),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_58),
.C(n_59),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_30),
.B1(n_28),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_55),
.B1(n_33),
.B2(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_30),
.B1(n_20),
.B2(n_19),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_20),
.B(n_17),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_30),
.B1(n_18),
.B2(n_19),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_63),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_31),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_74),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_75),
.B(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_16),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_26),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_86),
.C(n_43),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_90),
.B1(n_101),
.B2(n_32),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_87),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_45),
.C(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_30),
.B1(n_16),
.B2(n_20),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_32),
.B(n_26),
.Y(n_114)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_24),
.B1(n_35),
.B2(n_34),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_32),
.B1(n_28),
.B2(n_33),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_34),
.B1(n_35),
.B2(n_17),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_40),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_122),
.B1(n_132),
.B2(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_0),
.B(n_1),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_117),
.B(n_120),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_128),
.B1(n_91),
.B2(n_21),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_86),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_39),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_103),
.B1(n_88),
.B2(n_87),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_98),
.B1(n_65),
.B2(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_100),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_39),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_147),
.B(n_150),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_138),
.A2(n_141),
.B1(n_146),
.B2(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_142),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_72),
.B1(n_74),
.B2(n_68),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_100),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_161),
.C(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_63),
.B1(n_80),
.B2(n_78),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_121),
.B1(n_108),
.B2(n_130),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_38),
.B1(n_94),
.B2(n_89),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_2),
.B(n_3),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_109),
.B1(n_119),
.B2(n_125),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_40),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_134),
.B1(n_116),
.B2(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_21),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_112),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_158),
.Y(n_168)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_36),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_21),
.B(n_85),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_109),
.B(n_113),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_129),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_106),
.A2(n_95),
.B1(n_82),
.B2(n_12),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_121),
.B1(n_130),
.B2(n_123),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_21),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_25),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_135),
.C(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_112),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_170),
.B1(n_159),
.B2(n_150),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_108),
.B1(n_107),
.B2(n_127),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_180),
.B1(n_190),
.B2(n_150),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_124),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_182),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_181),
.Y(n_223)
);

AO22x1_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_109),
.B1(n_133),
.B2(n_123),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_162),
.Y(n_182)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_183),
.A2(n_2),
.B(n_3),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_109),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_192),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_185),
.B(n_188),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_113),
.B1(n_119),
.B2(n_29),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_187),
.B(n_191),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_113),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_161),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_139),
.B(n_29),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_197),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_144),
.A3(n_149),
.B1(n_160),
.B2(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_216),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_143),
.C(n_137),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_219),
.C(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_194),
.B(n_163),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_213),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

XOR2x1_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_147),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_207),
.B(n_186),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_223),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_137),
.B1(n_136),
.B2(n_158),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_211),
.B1(n_217),
.B2(n_169),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_137),
.B1(n_150),
.B2(n_138),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_183),
.A2(n_168),
.B(n_171),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_212),
.A2(n_178),
.B(n_176),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_148),
.C(n_141),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_185),
.B(n_146),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_227),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_148),
.B1(n_15),
.B2(n_14),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_25),
.C(n_23),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_36),
.C(n_13),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_225),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_170),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_3),
.C(n_4),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_197),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_242),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_208),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_248),
.B1(n_216),
.B2(n_237),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_174),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_249),
.B1(n_204),
.B2(n_174),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_226),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_199),
.Y(n_263)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_202),
.CI(n_207),
.CON(n_253),
.SN(n_253)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_209),
.B1(n_212),
.B2(n_217),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_252),
.A2(n_190),
.B1(n_234),
.B2(n_232),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_204),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_254),
.A2(n_245),
.B1(n_233),
.B2(n_230),
.Y(n_273)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_226),
.C(n_219),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_261),
.C(n_262),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_202),
.C(n_191),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_189),
.C(n_165),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_264),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_175),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_165),
.C(n_187),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_267),
.C(n_181),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_249),
.C(n_233),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_218),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_196),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_275),
.B1(n_252),
.B2(n_270),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_240),
.B1(n_241),
.B2(n_231),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_229),
.B(n_234),
.Y(n_276)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_271),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_232),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_264),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_284),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_193),
.C(n_181),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_267),
.C(n_265),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_221),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_284),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_193),
.B(n_5),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_287),
.B(n_4),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_4),
.C(n_5),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_257),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_294),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_286),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_291),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_274),
.B1(n_285),
.B2(n_281),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_268),
.B1(n_251),
.B2(n_261),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_300),
.B1(n_301),
.B2(n_277),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_297),
.C(n_283),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_253),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_298),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_253),
.B1(n_6),
.B2(n_7),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_8),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_299),
.A2(n_274),
.B1(n_278),
.B2(n_280),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_280),
.B1(n_277),
.B2(n_7),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_308),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_293),
.A2(n_296),
.B1(n_295),
.B2(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_309),
.B(n_295),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_312),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_294),
.C(n_6),
.Y(n_312)
);

AOI211xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_8),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_316),
.B(n_9),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_310),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_312),
.B1(n_317),
.B2(n_302),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_321),
.B(n_314),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_318),
.B(n_303),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_322),
.B(n_10),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_326),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_10),
.B(n_11),
.Y(n_329)
);


endmodule