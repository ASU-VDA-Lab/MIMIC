module real_jpeg_11145_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_302, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_302;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_300;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx24_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_65),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_65),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_3),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_151),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_3),
.A2(n_40),
.B1(n_49),
.B2(n_151),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g77 ( 
.A(n_7),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_8),
.A2(n_36),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_10),
.A2(n_40),
.B1(n_49),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_10),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_100),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_100),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_100),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_11),
.A2(n_40),
.B1(n_49),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_12),
.A2(n_57),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_12),
.B(n_57),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_12),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_12),
.A2(n_27),
.B1(n_33),
.B2(n_162),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_51),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_12),
.A2(n_42),
.B(n_46),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_12),
.A2(n_40),
.B1(n_49),
.B2(n_160),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_14),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_142),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_142),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_14),
.A2(n_40),
.B1(n_49),
.B2(n_142),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_15),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_74),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_15),
.A2(n_40),
.B1(n_49),
.B2(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_20),
.B(n_108),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_21),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_21),
.B(n_293),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_70),
.CI(n_89),
.CON(n_21),
.SN(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_54),
.B2(n_69),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_25),
.A2(n_38),
.B(n_69),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_25),
.A2(n_26),
.B1(n_55),
.B2(n_290),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_27),
.A2(n_33),
.B1(n_141),
.B2(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_27),
.A2(n_94),
.B(n_144),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_27),
.A2(n_34),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_27),
.A2(n_33),
.B1(n_207),
.B2(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_27),
.A2(n_193),
.B(n_229),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_28),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_28),
.A2(n_32),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_29),
.A2(n_30),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_29),
.B(n_63),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_29),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_30),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_152)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_32),
.B(n_35),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_32),
.B(n_93),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_33),
.B(n_160),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_33),
.A2(n_92),
.B(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_47),
.B(n_50),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_39),
.A2(n_99),
.B(n_101),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_39),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_39),
.A2(n_44),
.B1(n_243),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_39),
.A2(n_44),
.B1(n_99),
.B2(n_252),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_40),
.A2(n_41),
.B(n_160),
.C(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_44),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_76),
.B(n_78),
.C(n_79),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_76),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g185 ( 
.A(n_46),
.B(n_160),
.CON(n_185),
.SN(n_185)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_48),
.B(n_51),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_51),
.A2(n_116),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_55),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_64),
.B(n_66),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_62),
.B1(n_64),
.B2(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_56),
.A2(n_62),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_56),
.A2(n_62),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_56),
.A2(n_62),
.B1(n_150),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_56),
.A2(n_62),
.B1(n_175),
.B2(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_56),
.A2(n_82),
.B(n_183),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_58),
.B1(n_76),
.B2(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_57),
.B(n_76),
.Y(n_191)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_58),
.A2(n_78),
.B1(n_185),
.B2(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_62),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_62),
.A2(n_85),
.B(n_96),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_67),
.A2(n_84),
.B(n_87),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_81),
.B(n_88),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_81),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_75),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_75),
.A2(n_79),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_75),
.A2(n_123),
.B(n_255),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_79),
.B(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_110),
.B1(n_111),
.B2(n_128),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_88),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.C(n_102),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_90),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_91),
.B(n_95),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_104),
.B(n_160),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_104),
.A2(n_120),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_104),
.A2(n_120),
.B1(n_203),
.B2(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_129),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_119),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_120),
.A2(n_239),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_280),
.A3(n_292),
.B1(n_294),
.B2(n_300),
.C(n_302),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_245),
.C(n_276),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_219),
.B(n_244),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_196),
.B(n_218),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_178),
.B(n_195),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_169),
.B(n_177),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_157),
.B(n_168),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_145),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_152),
.B2(n_156),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_163),
.B(n_167),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_171),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_172),
.B(n_179),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.CI(n_176),
.CON(n_172),
.SN(n_172)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_189),
.B2(n_194),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_184),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_188),
.C(n_194),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_192),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_212),
.B2(n_213),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_215),
.C(n_216),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_204),
.B1(n_205),
.B2(n_211),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_206),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_208),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_209),
.C(n_211),
.Y(n_230)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_215),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_221),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_223),
.B(n_232),
.C(n_233),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_240),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_237),
.C(n_240),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_263),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_246),
.B(n_263),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_257),
.C(n_261),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_250),
.C(n_256),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_256),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_272),
.C(n_273),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_268),
.C(n_271),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_281),
.A2(n_295),
.B(n_299),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_283),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.C(n_291),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_295)
);


endmodule