module fake_jpeg_799_n_562 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_562);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_562;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_6),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_20),
.Y(n_54)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_59),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_69),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_65),
.B(n_68),
.Y(n_156)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_84),
.Y(n_114)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

OR2x2_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_51),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_78),
.A2(n_103),
.B(n_51),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_80),
.B(n_93),
.Y(n_159)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_38),
.B(n_1),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_36),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_92),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_2),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_95),
.Y(n_149)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_24),
.B(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_32),
.Y(n_163)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_40),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_41),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_21),
.B1(n_47),
.B2(n_43),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_117),
.B(n_33),
.Y(n_173)
);

OR2x4_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_67),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_65),
.B(n_68),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_146),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_82),
.A2(n_45),
.B1(n_47),
.B2(n_21),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_137),
.A2(n_141),
.B1(n_143),
.B2(n_34),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_75),
.A2(n_21),
.B1(n_47),
.B2(n_43),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_142),
.B1(n_28),
.B2(n_97),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_82),
.A2(n_45),
.B1(n_19),
.B2(n_43),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_55),
.A2(n_45),
.B1(n_19),
.B2(n_42),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_67),
.A2(n_32),
.B1(n_42),
.B2(n_22),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_51),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_163),
.C(n_28),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_78),
.B(n_42),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_53),
.A2(n_41),
.B(n_37),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_33),
.B(n_37),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_58),
.A2(n_87),
.B1(n_62),
.B2(n_66),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_153),
.A2(n_154),
.B1(n_162),
.B2(n_95),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_30),
.B1(n_22),
.B2(n_25),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_54),
.B(n_52),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_160),
.B(n_94),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_71),
.A2(n_30),
.B1(n_22),
.B2(n_25),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_79),
.B(n_32),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_30),
.Y(n_169)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_168),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_169),
.B(n_190),
.Y(n_246)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_170),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_171),
.A2(n_180),
.B1(n_229),
.B2(n_128),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_34),
.B1(n_33),
.B2(n_41),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_172),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_173),
.B(n_203),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_81),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_174),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_101),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_175),
.B(n_176),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_112),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_177),
.A2(n_207),
.B1(n_216),
.B2(n_222),
.Y(n_232)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_122),
.A2(n_88),
.B1(n_96),
.B2(n_83),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_210),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_108),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_185),
.B(n_188),
.Y(n_241)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_132),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_77),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_114),
.B(n_64),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_192),
.B(n_201),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_115),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_193),
.B(n_199),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_105),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_197),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_195),
.A2(n_130),
.B(n_13),
.Y(n_263)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_106),
.B(n_37),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_134),
.B(n_61),
.Y(n_201)
);

INVx5_ASAP7_75t_SL g202 ( 
.A(n_113),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_202),
.Y(n_264)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_205),
.B(n_215),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_206),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_72),
.B1(n_63),
.B2(n_34),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_209),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_95),
.C(n_103),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_212),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_121),
.B(n_95),
.C(n_91),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_89),
.C(n_76),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_218),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_121),
.B(n_17),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_137),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_158),
.B(n_3),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_12),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_144),
.B(n_3),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_225),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_143),
.A2(n_141),
.B1(n_127),
.B2(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_223),
.B1(n_155),
.B2(n_130),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_109),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_111),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_123),
.B(n_7),
.C(n_10),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_226),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_128),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_126),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_228),
.Y(n_281)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_165),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_177),
.A2(n_127),
.B1(n_111),
.B2(n_149),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_235),
.A2(n_242),
.B1(n_251),
.B2(n_260),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_236),
.A2(n_250),
.B1(n_265),
.B2(n_269),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_239),
.B(n_248),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_198),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_203),
.A2(n_120),
.B1(n_151),
.B2(n_164),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_175),
.A2(n_155),
.B1(n_164),
.B2(n_151),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_196),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_256),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_197),
.A2(n_164),
.B1(n_151),
.B2(n_120),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_178),
.B(n_149),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_261),
.B(n_214),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_263),
.A2(n_268),
.B(n_280),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_219),
.A2(n_131),
.B1(n_14),
.B2(n_15),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_273),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_173),
.A2(n_131),
.B(n_15),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_193),
.A2(n_180),
.B1(n_208),
.B2(n_176),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_213),
.A2(n_131),
.B1(n_15),
.B2(n_16),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_174),
.B(n_14),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_190),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_276),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_190),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_174),
.A2(n_14),
.B(n_16),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_241),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g341 ( 
.A(n_286),
.B(n_287),
.C(n_292),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_281),
.Y(n_287)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_293),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_281),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_258),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_183),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_295),
.B(n_321),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_SL g297 ( 
.A(n_233),
.B(n_174),
.C(n_187),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_297),
.Y(n_348)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_298),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_189),
.C(n_211),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_299),
.B(n_305),
.C(n_318),
.Y(n_338)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_271),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_315),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_244),
.B(n_208),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_302),
.B(n_231),
.Y(n_344)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_304),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_244),
.B(n_168),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_207),
.B1(n_216),
.B2(n_208),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_307),
.A2(n_310),
.B1(n_326),
.B2(n_282),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_224),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_312),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_232),
.A2(n_229),
.B1(n_209),
.B2(n_186),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g311 ( 
.A1(n_279),
.A2(n_226),
.B(n_212),
.C(n_202),
.Y(n_311)
);

AO21x2_ASAP7_75t_SL g351 ( 
.A1(n_311),
.A2(n_277),
.B(n_278),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_249),
.B(n_226),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

A2O1A1O1Ixp25_ASAP7_75t_L g316 ( 
.A1(n_234),
.A2(n_181),
.B(n_170),
.C(n_179),
.D(n_226),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_316),
.A2(n_256),
.B(n_248),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_279),
.A2(n_232),
.B1(n_239),
.B2(n_233),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_317),
.A2(n_322),
.B1(n_265),
.B2(n_264),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_225),
.C(n_184),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_246),
.B(n_227),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_319),
.B(n_240),
.C(n_237),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_259),
.A2(n_200),
.B(n_228),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_259),
.B(n_280),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_217),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_233),
.A2(n_206),
.B1(n_16),
.B2(n_17),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_257),
.B(n_274),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_323),
.B(n_333),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_272),
.B(n_254),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_327),
.Y(n_368)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_247),
.B(n_268),
.CI(n_257),
.CON(n_325),
.SN(n_325)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_275),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_236),
.A2(n_252),
.B1(n_235),
.B2(n_250),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_271),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_272),
.B(n_253),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_328),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_267),
.B(n_252),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_331),
.Y(n_349)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_330),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_252),
.B(n_262),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_230),
.Y(n_332)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_332),
.Y(n_377)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_230),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_263),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_334),
.B(n_336),
.C(n_347),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_273),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_313),
.A2(n_242),
.B(n_276),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g399 ( 
.A1(n_337),
.A2(n_351),
.B(n_361),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_SL g400 ( 
.A1(n_340),
.A2(n_343),
.B(n_360),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_344),
.B(n_350),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_329),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_231),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_296),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_366),
.Y(n_378)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_375),
.C(n_291),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_371),
.B1(n_352),
.B2(n_354),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_289),
.A2(n_237),
.B1(n_275),
.B2(n_282),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_359),
.A2(n_372),
.B1(n_333),
.B2(n_306),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_307),
.A2(n_277),
.B(n_245),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_278),
.B(n_240),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_294),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_365),
.B(n_298),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_305),
.B(n_245),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_318),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_289),
.A2(n_237),
.B1(n_326),
.B2(n_312),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_310),
.A2(n_309),
.B1(n_311),
.B2(n_284),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_288),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_376),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_317),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_291),
.B(n_302),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_379),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_380),
.B(n_397),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_381),
.A2(n_384),
.B1(n_390),
.B2(n_391),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_327),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_382),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_341),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_392),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_351),
.A2(n_311),
.B1(n_290),
.B2(n_323),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_363),
.B(n_301),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_387),
.B(n_396),
.Y(n_431)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_352),
.Y(n_388)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_351),
.A2(n_311),
.B1(n_285),
.B2(n_316),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_345),
.A2(n_311),
.B1(n_285),
.B2(n_323),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_368),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_346),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_413),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_371),
.A2(n_322),
.B1(n_325),
.B2(n_313),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_394),
.A2(n_404),
.B1(n_415),
.B2(n_407),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_R g426 ( 
.A(n_395),
.B(n_374),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_303),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_300),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_401),
.Y(n_428)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_345),
.B(n_332),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_403),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_360),
.A2(n_351),
.B1(n_375),
.B2(n_340),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_411),
.B1(n_377),
.B2(n_361),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_304),
.Y(n_406)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_406),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_337),
.B(n_330),
.Y(n_407)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_353),
.A2(n_373),
.B1(n_355),
.B2(n_342),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_376),
.A2(n_359),
.B1(n_349),
.B2(n_356),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_348),
.B(n_336),
.Y(n_412)
);

OAI21xp33_ASAP7_75t_L g422 ( 
.A1(n_412),
.A2(n_339),
.B(n_344),
.Y(n_422)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_364),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_348),
.A2(n_335),
.B1(n_343),
.B2(n_360),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_414),
.A2(n_342),
.B(n_384),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_334),
.A2(n_349),
.B1(n_347),
.B2(n_370),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_378),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_422),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_338),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_419),
.B(n_443),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_367),
.C(n_364),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_423),
.B(n_430),
.C(n_436),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_429),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_378),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_367),
.C(n_374),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_406),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_392),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_377),
.C(n_355),
.Y(n_436)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_437),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_441),
.A2(n_402),
.B(n_413),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_380),
.B(n_389),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_409),
.C(n_386),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_447),
.C(n_388),
.Y(n_461)
);

OA22x2_ASAP7_75t_L g445 ( 
.A1(n_404),
.A2(n_414),
.B1(n_399),
.B2(n_410),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_383),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_446),
.A2(n_399),
.B1(n_393),
.B2(n_381),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_386),
.B(n_391),
.C(n_410),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_394),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_444),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_435),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_452),
.B(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_454),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_441),
.A2(n_399),
.B(n_400),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_455),
.A2(n_464),
.B(n_445),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_456),
.A2(n_463),
.B1(n_472),
.B2(n_445),
.Y(n_488)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_458),
.Y(n_491)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_459),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_430),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_461),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_443),
.B(n_401),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_474),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_446),
.A2(n_424),
.B1(n_437),
.B2(n_418),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_425),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_427),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_466),
.Y(n_479)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_467),
.Y(n_494)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_398),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_475),
.Y(n_498)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_428),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_470),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_424),
.A2(n_418),
.B1(n_448),
.B2(n_440),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_419),
.B(n_433),
.C(n_436),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_433),
.C(n_434),
.Y(n_483)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

INVx13_ASAP7_75t_L g477 ( 
.A(n_476),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_451),
.A2(n_440),
.B1(n_447),
.B2(n_427),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_480),
.A2(n_482),
.B1(n_488),
.B2(n_484),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_451),
.A2(n_426),
.B1(n_434),
.B2(n_445),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_485),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_484),
.A2(n_492),
.B(n_498),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_460),
.C(n_473),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_471),
.C(n_461),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_490),
.C(n_499),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_431),
.C(n_420),
.Y(n_490)
);

INVx13_ASAP7_75t_L g497 ( 
.A(n_464),
.Y(n_497)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_497),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_462),
.C(n_472),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_502),
.A2(n_510),
.B1(n_517),
.B2(n_514),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_458),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_506),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_505),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_463),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_479),
.B(n_469),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_509),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_479),
.A2(n_453),
.B(n_455),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_508),
.A2(n_516),
.B(n_489),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_456),
.C(n_449),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_482),
.A2(n_476),
.B(n_467),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_510),
.A2(n_494),
.B1(n_496),
.B2(n_477),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_478),
.B(n_468),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_477),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_478),
.B(n_470),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_495),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_457),
.C(n_475),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_494),
.C(n_496),
.Y(n_529)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_488),
.B(n_491),
.CI(n_497),
.CON(n_514),
.SN(n_514)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_514),
.A2(n_481),
.B1(n_487),
.B2(n_489),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_485),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_517),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_491),
.A2(n_492),
.B(n_498),
.Y(n_516)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_518),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_520),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_521),
.A2(n_516),
.B(n_507),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_505),
.A2(n_504),
.B(n_500),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_522),
.A2(n_508),
.B(n_513),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_481),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_524),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_509),
.B(n_486),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_487),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_525),
.B(n_503),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_529),
.Y(n_533)
);

AOI21xp33_ASAP7_75t_L g539 ( 
.A1(n_531),
.A2(n_514),
.B(n_501),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_515),
.Y(n_540)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_536),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_537),
.A2(n_539),
.B(n_542),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_538),
.B(n_519),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_540),
.B(n_543),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_L g542 ( 
.A(n_526),
.B(n_501),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_526),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g544 ( 
.A(n_534),
.B(n_524),
.Y(n_544)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_544),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_547),
.B(n_550),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_537),
.A2(n_530),
.B(n_527),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_548),
.A2(n_531),
.B(n_541),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_533),
.C(n_519),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_551),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_547),
.Y(n_552)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_552),
.Y(n_556)
);

AOI31xp33_ASAP7_75t_L g557 ( 
.A1(n_554),
.A2(n_549),
.A3(n_545),
.B(n_546),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_557),
.A2(n_541),
.B(n_520),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_556),
.B(n_553),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_558),
.B(n_559),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_555),
.B(n_525),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_523),
.Y(n_562)
);


endmodule