module fake_jpeg_23936_n_68 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_R g14 ( 
.A(n_5),
.B(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_1),
.C(n_3),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_1),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_29),
.B1(n_15),
.B2(n_16),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_10),
.B1(n_16),
.B2(n_20),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_15),
.B1(n_11),
.B2(n_17),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_40),
.B1(n_30),
.B2(n_27),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_12),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_23),
.A2(n_13),
.B1(n_21),
.B2(n_12),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_47),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_49),
.B1(n_32),
.B2(n_36),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_27),
.B(n_22),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_41),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_12),
.CI(n_21),
.CON(n_47),
.SN(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_13),
.B1(n_21),
.B2(n_34),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_53),
.Y(n_60)
);

XOR2x1_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_47),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_45),
.B1(n_49),
.B2(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_59),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_42),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_42),
.C(n_44),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_60),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_50),
.C(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_62),
.C(n_61),
.Y(n_67)
);

AOI211xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_65),
.B(n_61),
.C(n_63),
.Y(n_68)
);


endmodule