module fake_jpeg_29175_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_42),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_3),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_15),
.Y(n_60)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_17),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_47),
.B(n_74),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_23),
.B1(n_31),
.B2(n_21),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_68),
.Y(n_77)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_30),
.B1(n_29),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_63),
.B1(n_7),
.B2(n_10),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_30),
.C(n_32),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_56),
.B(n_70),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_16),
.B1(n_28),
.B2(n_26),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_14),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_21),
.B1(n_31),
.B2(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_32),
.C(n_28),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_35),
.B(n_1),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_4),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_35),
.A2(n_16),
.B1(n_25),
.B2(n_20),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_40),
.B1(n_37),
.B2(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_88),
.Y(n_113)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_98),
.B1(n_59),
.B2(n_67),
.Y(n_126)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_51),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_13),
.B1(n_14),
.B2(n_48),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_106),
.B1(n_59),
.B2(n_62),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_13),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_50),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_51),
.A2(n_57),
.B1(n_71),
.B2(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_112),
.B(n_114),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_57),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_118),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_86),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_136),
.B1(n_92),
.B2(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_49),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_122),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_55),
.C(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_55),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_128),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_67),
.C(n_64),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_88),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_96),
.A2(n_91),
.B1(n_82),
.B2(n_90),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_110),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_102),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_115),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_93),
.B1(n_105),
.B2(n_81),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_78),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_137),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_78),
.C(n_105),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_92),
.B1(n_119),
.B2(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_134),
.B1(n_112),
.B2(n_120),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_112),
.B(n_116),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_161),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_128),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_156),
.B(n_118),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_125),
.B1(n_149),
.B2(n_138),
.C(n_154),
.Y(n_177)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_109),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_108),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_179),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_111),
.Y(n_173)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_172),
.B(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_111),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_153),
.C(n_148),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_173),
.B(n_152),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_125),
.C(n_155),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_158),
.C(n_145),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_176),
.C(n_141),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_194),
.B(n_195),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_148),
.B(n_144),
.C(n_146),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_196),
.B1(n_163),
.B2(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_142),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_185),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_176),
.C(n_163),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_179),
.C(n_178),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_213),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_205),
.A2(n_183),
.B1(n_192),
.B2(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_183),
.B(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_217),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_199),
.C(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_220),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_208),
.C(n_197),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_215),
.B(n_198),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_169),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_169),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_215),
.B1(n_188),
.B2(n_189),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_227),
.Y(n_231)
);

AOI31xp67_ASAP7_75t_L g227 ( 
.A1(n_218),
.A2(n_198),
.A3(n_212),
.B(n_165),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_229),
.B(n_222),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_232),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_222),
.B1(n_151),
.B2(n_157),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_228),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_160),
.B1(n_175),
.B2(n_226),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_234),
.A2(n_225),
.B(n_159),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_236),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_160),
.Y(n_238)
);


endmodule