module fake_netlist_6_4712_n_2611 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_537, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2611);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_537;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2611;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_2496;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_2590;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_2585;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_2203;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_290),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_108),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_208),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_478),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_264),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_500),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_387),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_221),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_45),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_354),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_21),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_114),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_254),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_536),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_89),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_331),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_355),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_432),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_6),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_307),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_523),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_283),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_509),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_528),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_243),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_282),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_133),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_139),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_177),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_470),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_51),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_61),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_401),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_147),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_296),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_139),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_513),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_397),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_442),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_530),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_450),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_516),
.Y(n_581)
);

CKINVDCx16_ASAP7_75t_R g582 ( 
.A(n_253),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_328),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_25),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_196),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_42),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_389),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_484),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_526),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_191),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_15),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_134),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_255),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_79),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_132),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_520),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_158),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_258),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_80),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_47),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_4),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_150),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_506),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_89),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_215),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_443),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_22),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_511),
.Y(n_608)
);

CKINVDCx14_ASAP7_75t_R g609 ( 
.A(n_83),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_372),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_527),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_485),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_120),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_273),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_309),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_188),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_99),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_233),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_87),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_533),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_176),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_263),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_218),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_440),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_435),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_296),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_273),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_515),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_421),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_33),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_72),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_466),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_147),
.Y(n_633)
);

BUFx8_ASAP7_75t_SL g634 ( 
.A(n_287),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_52),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_73),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_371),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_152),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_77),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_345),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_345),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_193),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_501),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_2),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_159),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_107),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_126),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_290),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_217),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_276),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_525),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_102),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_274),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_302),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_211),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_469),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_408),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_192),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_32),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_82),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_529),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_458),
.Y(n_663)
);

INVxp67_ASAP7_75t_SL g664 ( 
.A(n_465),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_201),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_323),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_399),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_268),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_118),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_517),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_512),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_229),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_510),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_481),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_150),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_305),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_534),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_297),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_183),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_158),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_182),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_72),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_334),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_467),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_505),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_16),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_531),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_521),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_378),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_255),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_420),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_204),
.Y(n_692)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_99),
.Y(n_693)
);

CKINVDCx11_ASAP7_75t_R g694 ( 
.A(n_329),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_172),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_30),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_532),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_319),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_55),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_91),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_183),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_503),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_411),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_92),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_359),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_480),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_187),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_462),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_496),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_214),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_502),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_315),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_242),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_522),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_519),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_377),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_176),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_477),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_429),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_105),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_260),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_436),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_472),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_354),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_445),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_82),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_127),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_333),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_80),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_347),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_100),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_518),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_424),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_67),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_310),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_36),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_117),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_330),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_295),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_182),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_514),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_451),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_419),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_488),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_269),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_22),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_476),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_41),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_109),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_487),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_524),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_309),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_209),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_159),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_142),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_372),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_74),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_268),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_64),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_254),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_39),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_344),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_441),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_267),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_3),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_98),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_111),
.Y(n_767)
);

BUFx8_ASAP7_75t_SL g768 ( 
.A(n_507),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_504),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_535),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_461),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_694),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_694),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_724),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_634),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_744),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_634),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_724),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_731),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_610),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_546),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_731),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_553),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_621),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_546),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_542),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_546),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_553),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_609),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_546),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_544),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_552),
.Y(n_792)
);

INVxp33_ASAP7_75t_SL g793 ( 
.A(n_650),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_662),
.B(n_0),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_560),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_584),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_629),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_567),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_584),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_584),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_660),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_584),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_623),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_623),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_623),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_623),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_562),
.Y(n_807)
);

CKINVDCx14_ASAP7_75t_R g808 ( 
.A(n_609),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_612),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_629),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_638),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_638),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_638),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_638),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_567),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_647),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_647),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_647),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_563),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_647),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_745),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_745),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_745),
.Y(n_823)
);

INVxp33_ASAP7_75t_L g824 ( 
.A(n_675),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_745),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_612),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_540),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_547),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_550),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_555),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_558),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_559),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_591),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_565),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_578),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_582),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_595),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_570),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_588),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_589),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_574),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_575),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_583),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_608),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_590),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_592),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_595),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_593),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_620),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_591),
.Y(n_850)
);

CKINVDCx20_ASAP7_75t_R g851 ( 
.A(n_640),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_642),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_594),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_597),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_640),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_549),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_653),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_600),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_605),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_653),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_607),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_690),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_693),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_616),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_617),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_627),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_549),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_631),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_637),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_639),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_646),
.Y(n_871)
);

INVxp67_ASAP7_75t_SL g872 ( 
.A(n_684),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_662),
.B(n_0),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_654),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_625),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_797),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_785),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_787),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_786),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_783),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_791),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_792),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_797),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_790),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_796),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_795),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_799),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_783),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_800),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_807),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_788),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_819),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_835),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_803),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_788),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_810),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_798),
.Y(n_897)
);

INVxp33_ASAP7_75t_SL g898 ( 
.A(n_777),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_839),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_804),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_840),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_844),
.B(n_572),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_805),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_806),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_872),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_849),
.B(n_662),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_798),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_811),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_875),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_812),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_813),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_815),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_814),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_775),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_816),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_775),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_817),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_818),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_781),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_863),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_809),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_821),
.Y(n_922)
);

INVxp67_ASAP7_75t_SL g923 ( 
.A(n_809),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_815),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_822),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_837),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_863),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_789),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_789),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_781),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_823),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_773),
.Y(n_932)
);

CKINVDCx16_ASAP7_75t_R g933 ( 
.A(n_808),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_773),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_772),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_808),
.B(n_684),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_776),
.B(n_733),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_772),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_837),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_847),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_847),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_919),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_896),
.B(n_802),
.Y(n_943)
);

CKINVDCx6p67_ASAP7_75t_R g944 ( 
.A(n_933),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_905),
.B(n_802),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_876),
.Y(n_946)
);

OA21x2_ASAP7_75t_L g947 ( 
.A1(n_919),
.A2(n_820),
.B(n_825),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_877),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_878),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_884),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_883),
.B(n_833),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_879),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_885),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_887),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_881),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_921),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_902),
.B(n_867),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_889),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_921),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_894),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_SL g961 ( 
.A1(n_880),
.A2(n_707),
.B1(n_717),
.B2(n_690),
.Y(n_961)
);

CKINVDCx20_ASAP7_75t_R g962 ( 
.A(n_880),
.Y(n_962)
);

CKINVDCx11_ASAP7_75t_R g963 ( 
.A(n_888),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_900),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_930),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_921),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_928),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_930),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_903),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_921),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_904),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_908),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_910),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_929),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_911),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_906),
.B(n_820),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_937),
.B(n_833),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_913),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_920),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_915),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_936),
.B(n_850),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_917),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_927),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_882),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_918),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_922),
.Y(n_986)
);

AND2x6_ASAP7_75t_L g987 ( 
.A(n_925),
.B(n_545),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_931),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_923),
.Y(n_989)
);

AND2x6_ASAP7_75t_L g990 ( 
.A(n_886),
.B(n_545),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_890),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_SL g992 ( 
.A1(n_888),
.A2(n_717),
.B1(n_735),
.B2(n_707),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_892),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_893),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_899),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_901),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_909),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_898),
.B(n_793),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_891),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_935),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_938),
.B(n_794),
.Y(n_1001)
);

AND2x6_ASAP7_75t_L g1002 ( 
.A(n_932),
.B(n_580),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_891),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_934),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_914),
.Y(n_1005)
);

INVx5_ASAP7_75t_L g1006 ( 
.A(n_916),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_941),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_941),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_895),
.B(n_850),
.Y(n_1009)
);

CKINVDCx16_ASAP7_75t_R g1010 ( 
.A(n_895),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_940),
.B(n_873),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_897),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_940),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_897),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_907),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_907),
.B(n_852),
.Y(n_1016)
);

NOR2x1_ASAP7_75t_L g1017 ( 
.A(n_912),
.B(n_576),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_912),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_939),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_924),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_924),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_926),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_926),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_939),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_896),
.B(n_852),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_896),
.A2(n_793),
.B1(n_801),
.B2(n_824),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_919),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_896),
.B(n_733),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_921),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_936),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_962),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_947),
.Y(n_1032)
);

AND3x1_ASAP7_75t_L g1033 ( 
.A(n_1009),
.B(n_853),
.C(n_836),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_958),
.Y(n_1034)
);

AND2x6_ASAP7_75t_L g1035 ( 
.A(n_977),
.B(n_580),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_SL g1036 ( 
.A1(n_961),
.A2(n_855),
.B1(n_857),
.B2(n_851),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_947),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_947),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_958),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_942),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_959),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_969),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_959),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_977),
.B(n_946),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_942),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_970),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_970),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_965),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_969),
.Y(n_1049)
);

AO22x1_ASAP7_75t_L g1050 ( 
.A1(n_1002),
.A2(n_824),
.B1(n_614),
.B2(n_721),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_1009),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_965),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_980),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_980),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_946),
.B(n_780),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_988),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1025),
.B(n_664),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_981),
.B(n_784),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_968),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1030),
.A2(n_587),
.B1(n_596),
.B2(n_576),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_981),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_968),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_990),
.A2(n_596),
.B1(n_603),
.B2(n_587),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_948),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_966),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_980),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1025),
.B(n_606),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_SL g1068 ( 
.A1(n_992),
.A2(n_855),
.B1(n_857),
.B2(n_851),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1027),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_949),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_950),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_951),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1027),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_990),
.A2(n_663),
.B1(n_677),
.B2(n_603),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_953),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_951),
.B(n_606),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_SL g1077 ( 
.A(n_1014),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_954),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_1014),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_980),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_1026),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_960),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_964),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_990),
.A2(n_677),
.B1(n_703),
.B2(n_663),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_972),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_966),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1016),
.B(n_856),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_973),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1016),
.B(n_774),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_SL g1090 ( 
.A(n_1005),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_966),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_978),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_971),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_985),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_1016),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_971),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_943),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_945),
.B(n_556),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_982),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_982),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_982),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_1028),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_979),
.B(n_983),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_976),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_989),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_990),
.A2(n_723),
.B1(n_703),
.B2(n_557),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_975),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_975),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_975),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_980),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_990),
.A2(n_1002),
.B1(n_957),
.B2(n_1011),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_986),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_986),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_986),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_990),
.B(n_688),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_986),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_986),
.Y(n_1117)
);

INVx6_ASAP7_75t_L g1118 ( 
.A(n_991),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_979),
.B(n_778),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1001),
.B(n_993),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_987),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_L g1122 ( 
.A(n_1000),
.B(n_723),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_987),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_987),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_987),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_987),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_991),
.B(n_994),
.Y(n_1127)
);

NAND2x1_ASAP7_75t_L g1128 ( 
.A(n_956),
.B(n_612),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_956),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_956),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_995),
.B(n_630),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_987),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1029),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1029),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1029),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1002),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_1002),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_994),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1002),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1002),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_996),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_997),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_1007),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_997),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_991),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_991),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1007),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_991),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_967),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_962),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_967),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_974),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_998),
.B(n_612),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_974),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_983),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1017),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1008),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_952),
.B(n_688),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1008),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1015),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1021),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1020),
.Y(n_1162)
);

INVx3_ASAP7_75t_SL g1163 ( 
.A(n_944),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1021),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1006),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1006),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_952),
.A2(n_748),
.B1(n_764),
.B2(n_735),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1040),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1044),
.B(n_984),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1159),
.B(n_1006),
.Y(n_1170)
);

INVx6_ASAP7_75t_L g1171 ( 
.A(n_1103),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1041),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1055),
.B(n_984),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1040),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1045),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1045),
.Y(n_1176)
);

CKINVDCx16_ASAP7_75t_R g1177 ( 
.A(n_1077),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1041),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1048),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1058),
.B(n_955),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1048),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1052),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1052),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1051),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1097),
.B(n_955),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1141),
.B(n_1006),
.Y(n_1186)
);

AOI22x1_ASAP7_75t_SL g1187 ( 
.A1(n_1031),
.A2(n_862),
.B1(n_860),
.B2(n_999),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1079),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1102),
.B(n_579),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1093),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1101),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1093),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1051),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1102),
.B(n_581),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1101),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1041),
.Y(n_1196)
);

BUFx4f_ASAP7_75t_L g1197 ( 
.A(n_1163),
.Y(n_1197)
);

AND2x6_ASAP7_75t_L g1198 ( 
.A(n_1137),
.B(n_1005),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1072),
.B(n_611),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1041),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1087),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1120),
.B(n_1022),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1059),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_1118),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1141),
.B(n_1006),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1060),
.B(n_1150),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1100),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1142),
.B(n_1005),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1119),
.B(n_1004),
.Y(n_1209)
);

BUFx10_ASAP7_75t_L g1210 ( 
.A(n_1090),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1095),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1059),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1120),
.B(n_860),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1062),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1090),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1159),
.B(n_1005),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1062),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1131),
.B(n_862),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1043),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1147),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1043),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1035),
.A2(n_716),
.B1(n_628),
.B2(n_632),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1069),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1118),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1043),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1100),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1043),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1163),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1089),
.Y(n_1229)
);

CKINVDCx11_ASAP7_75t_R g1230 ( 
.A(n_1151),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1157),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1161),
.B(n_1005),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_SL g1233 ( 
.A(n_1063),
.B(n_1012),
.C(n_1019),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1142),
.B(n_1004),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1035),
.A2(n_716),
.B1(n_643),
.B2(n_657),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1074),
.A2(n_1013),
.B1(n_1018),
.B2(n_1023),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1077),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1161),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1072),
.B(n_624),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1104),
.B(n_674),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1065),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1096),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1118),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_L g1244 ( 
.A(n_1156),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1069),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1035),
.A2(n_711),
.B1(n_722),
.B2(n_709),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1034),
.Y(n_1247)
);

AND2x6_ASAP7_75t_L g1248 ( 
.A(n_1137),
.B(n_1004),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1057),
.B(n_725),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1131),
.B(n_1023),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1061),
.B(n_944),
.Y(n_1251)
);

AND2x6_ASAP7_75t_L g1252 ( 
.A(n_1137),
.B(n_1024),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1039),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1164),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1053),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1073),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1151),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1123),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1152),
.B(n_1024),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1081),
.B(n_1010),
.Y(n_1260)
);

AO22x2_ASAP7_75t_L g1261 ( 
.A1(n_1081),
.A2(n_551),
.B1(n_721),
.B2(n_614),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1099),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1046),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1145),
.B(n_827),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1053),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1046),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1035),
.A2(n_742),
.B1(n_750),
.B2(n_741),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1047),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1061),
.B(n_771),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1047),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1032),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1123),
.Y(n_1272)
);

AND2x6_ASAP7_75t_L g1273 ( 
.A(n_1137),
.B(n_569),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1152),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1138),
.B(n_1012),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1042),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1143),
.B(n_1019),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1032),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1038),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1065),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1123),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1123),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1038),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1056),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1086),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1145),
.B(n_577),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1086),
.Y(n_1287)
);

NAND3xp33_ASAP7_75t_L g1288 ( 
.A(n_1167),
.B(n_541),
.C(n_539),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1160),
.Y(n_1289)
);

NAND2xp33_ASAP7_75t_L g1290 ( 
.A(n_1035),
.B(n_651),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1049),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1144),
.B(n_1003),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1143),
.B(n_1149),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1107),
.B(n_715),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1160),
.B(n_1003),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1162),
.B(n_963),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1107),
.B(n_718),
.Y(n_1297)
);

INVx5_ASAP7_75t_L g1298 ( 
.A(n_1053),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1091),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1091),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1036),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1108),
.B(n_732),
.Y(n_1302)
);

AND2x6_ASAP7_75t_L g1303 ( 
.A(n_1136),
.B(n_642),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1108),
.B(n_656),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1064),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1084),
.A2(n_757),
.B1(n_764),
.B2(n_748),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1068),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1053),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1154),
.B(n_779),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1106),
.A2(n_757),
.B1(n_667),
.B2(n_670),
.Y(n_1310)
);

NOR2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1155),
.B(n_782),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1162),
.B(n_1127),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1146),
.B(n_661),
.Y(n_1313)
);

BUFx4f_ASAP7_75t_L g1314 ( 
.A(n_1148),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1098),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1070),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1054),
.Y(n_1317)
);

NAND2xp33_ASAP7_75t_L g1318 ( 
.A(n_1126),
.B(n_671),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1071),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1075),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1054),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1078),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1136),
.B(n_644),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1122),
.B(n_963),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1033),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1054),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1082),
.B(n_828),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1083),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1085),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1050),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1054),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1066),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1088),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1092),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1127),
.B(n_673),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1094),
.B(n_829),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1105),
.B(n_685),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1098),
.A2(n_551),
.B1(n_737),
.B2(n_726),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1037),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_SL g1340 ( 
.A(n_1165),
.B(n_768),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1158),
.B(n_635),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1109),
.Y(n_1342)
);

AND2x6_ASAP7_75t_L g1343 ( 
.A(n_1139),
.B(n_644),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1066),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1158),
.B(n_641),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1066),
.B(n_830),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1037),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1098),
.B(n_687),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1037),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1037),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1167),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1110),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1076),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1126),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1129),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1066),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1080),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1112),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_SL g1359 ( 
.A(n_1126),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1067),
.B(n_689),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1135),
.B(n_691),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1135),
.B(n_697),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1113),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1153),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1165),
.B(n_831),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1130),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1111),
.B(n_702),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1258),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1218),
.A2(n_1153),
.B1(n_1140),
.B2(n_1139),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1250),
.A2(n_1115),
.B(n_1140),
.C(n_659),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1247),
.Y(n_1371)
);

AND2x6_ASAP7_75t_SL g1372 ( 
.A(n_1296),
.B(n_655),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1253),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1353),
.B(n_1271),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1276),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_1172),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1185),
.B(n_1080),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1291),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1209),
.B(n_1169),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1180),
.B(n_1080),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1289),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1174),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1220),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1173),
.B(n_1080),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1271),
.B(n_1114),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1278),
.B(n_1117),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1345),
.A2(n_1121),
.B(n_1125),
.C(n_1124),
.Y(n_1387)
);

OR2x6_ASAP7_75t_L g1388 ( 
.A(n_1171),
.B(n_1126),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1172),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1312),
.B(n_1166),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1202),
.B(n_1166),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1238),
.Y(n_1392)
);

OR2x6_ASAP7_75t_SL g1393 ( 
.A(n_1351),
.B(n_543),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1216),
.B(n_1116),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1174),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1216),
.B(n_1130),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1175),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1232),
.B(n_1189),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1316),
.B(n_1229),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1232),
.B(n_1133),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1194),
.B(n_1133),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1175),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1244),
.B(n_1116),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1274),
.B(n_549),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1176),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1201),
.B(n_1132),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1176),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1244),
.B(n_1116),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1179),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1322),
.B(n_1116),
.Y(n_1410)
);

AOI22x1_ASAP7_75t_L g1411 ( 
.A1(n_1285),
.A2(n_1134),
.B1(n_706),
.B2(n_714),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1306),
.A2(n_708),
.B1(n_743),
.B2(n_719),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1179),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1181),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1181),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1213),
.B(n_648),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1182),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1305),
.B(n_658),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1231),
.B(n_1254),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1172),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1329),
.B(n_747),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1319),
.B(n_699),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1320),
.B(n_700),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1182),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1277),
.B(n_739),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1257),
.B(n_751),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1278),
.B(n_1128),
.Y(n_1427)
);

BUFx8_ASAP7_75t_L g1428 ( 
.A(n_1188),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1260),
.A2(n_769),
.B1(n_770),
.B2(n_763),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1349),
.B(n_666),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1293),
.Y(n_1431)
);

INVx8_ASAP7_75t_L g1432 ( 
.A(n_1198),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1249),
.B(n_672),
.Y(n_1433)
);

INVx8_ASAP7_75t_L g1434 ( 
.A(n_1198),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1328),
.B(n_548),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1171),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1284),
.B(n_832),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1251),
.B(n_834),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1170),
.B(n_838),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1183),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_1228),
.B(n_374),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1183),
.Y(n_1442)
);

AND2x2_ASAP7_75t_SL g1443 ( 
.A(n_1197),
.B(n_680),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1327),
.B(n_841),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1223),
.Y(n_1445)
);

AOI22x1_ASAP7_75t_L g1446 ( 
.A1(n_1285),
.A2(n_680),
.B1(n_710),
.B2(n_842),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1223),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1170),
.B(n_843),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1365),
.A2(n_768),
.B1(n_710),
.B2(n_678),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1314),
.B(n_845),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1333),
.B(n_554),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1334),
.B(n_561),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1191),
.B(n_682),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1314),
.B(n_1294),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1191),
.B(n_692),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1178),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1206),
.B(n_564),
.Y(n_1457)
);

INVxp67_ASAP7_75t_SL g1458 ( 
.A(n_1178),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1297),
.B(n_846),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1315),
.A2(n_854),
.B1(n_858),
.B2(n_848),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1302),
.B(n_566),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1199),
.B(n_568),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1258),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1184),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1310),
.B(n_1292),
.C(n_1295),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1330),
.B(n_859),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1311),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1298),
.B(n_861),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1193),
.B(n_571),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1298),
.B(n_864),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1239),
.B(n_573),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1195),
.B(n_695),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1168),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1258),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1301),
.A2(n_622),
.B1(n_665),
.B2(n_599),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_SL g1476 ( 
.A(n_1210),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1190),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1192),
.Y(n_1478)
);

NOR3xp33_ASAP7_75t_L g1479 ( 
.A(n_1233),
.B(n_866),
.C(n_865),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1269),
.B(n_585),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1298),
.B(n_868),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1195),
.B(n_698),
.Y(n_1482)
);

INVx8_ASAP7_75t_L g1483 ( 
.A(n_1198),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1203),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1262),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1240),
.B(n_586),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1264),
.B(n_598),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1275),
.A2(n_701),
.B(n_705),
.C(n_704),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1262),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1272),
.Y(n_1490)
);

INVx8_ASAP7_75t_L g1491 ( 
.A(n_1198),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1264),
.B(n_601),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1207),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1211),
.B(n_869),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1341),
.B(n_1236),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1178),
.B(n_870),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1288),
.B(n_604),
.C(n_602),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1364),
.B(n_613),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1200),
.B(n_1219),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1242),
.B(n_615),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1309),
.B(n_648),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1200),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1339),
.B(n_712),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1259),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1222),
.A2(n_728),
.B1(n_729),
.B2(n_727),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1272),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1200),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1307),
.B(n_618),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1226),
.Y(n_1509)
);

O2A1O1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1348),
.A2(n_740),
.B(n_753),
.C(n_752),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1212),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1327),
.A2(n_874),
.B1(n_871),
.B2(n_626),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1347),
.B(n_755),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1272),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1219),
.B(n_619),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1214),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1217),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1350),
.B(n_1279),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1235),
.A2(n_765),
.B1(n_767),
.B2(n_760),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1365),
.A2(n_648),
.B1(n_636),
.B2(n_645),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1340),
.A2(n_649),
.B1(n_652),
.B2(n_633),
.Y(n_1521)
);

INVx8_ASAP7_75t_L g1522 ( 
.A(n_1359),
.Y(n_1522)
);

BUFx8_ASAP7_75t_L g1523 ( 
.A(n_1325),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1245),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1342),
.A2(n_669),
.B(n_676),
.C(n_668),
.Y(n_1525)
);

NAND2xp33_ASAP7_75t_L g1526 ( 
.A(n_1248),
.B(n_762),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_SL g1527 ( 
.A(n_1359),
.B(n_686),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1336),
.B(n_1259),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1336),
.A2(n_681),
.B1(n_683),
.B2(n_679),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1324),
.B(n_696),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1360),
.B(n_713),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1221),
.B(n_720),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1187),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1252),
.A2(n_734),
.B1(n_736),
.B2(n_730),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1256),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1221),
.B(n_1225),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1234),
.B(n_738),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1252),
.A2(n_1273),
.B1(n_1335),
.B2(n_1323),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1252),
.A2(n_749),
.B1(n_754),
.B2(n_746),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1252),
.A2(n_758),
.B1(n_759),
.B2(n_756),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1221),
.B(n_761),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1337),
.B(n_766),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1273),
.A2(n_1323),
.B1(n_1343),
.B2(n_1303),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1355),
.B(n_1),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1366),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1230),
.B(n_1),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1358),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1263),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1225),
.B(n_809),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1279),
.B(n_1283),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1283),
.B(n_1241),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1281),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1241),
.B(n_375),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1358),
.B(n_376),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1225),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1215),
.B(n_2),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1227),
.B(n_809),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1266),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1227),
.B(n_826),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1227),
.B(n_826),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1338),
.B(n_3),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1243),
.B(n_826),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1261),
.B(n_4),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1268),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1243),
.B(n_1204),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1270),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1363),
.B(n_379),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1204),
.B(n_380),
.Y(n_1568)
);

INVxp67_ASAP7_75t_SL g1569 ( 
.A(n_1281),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1224),
.B(n_381),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1281),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1261),
.B(n_5),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1495),
.A2(n_1273),
.B1(n_1286),
.B2(n_1313),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1431),
.B(n_1177),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1374),
.B(n_1208),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1382),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1374),
.B(n_1273),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1428),
.Y(n_1579)
);

AOI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1465),
.A2(n_1352),
.B1(n_1363),
.B2(n_1248),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1457),
.A2(n_1323),
.B1(n_1343),
.B2(n_1303),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1508),
.A2(n_1323),
.B1(n_1343),
.B2(n_1303),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1381),
.B(n_1237),
.Y(n_1583)
);

INVx2_ASAP7_75t_SL g1584 ( 
.A(n_1428),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1419),
.B(n_1196),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1383),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1485),
.Y(n_1587)
);

INVx4_ASAP7_75t_L g1588 ( 
.A(n_1522),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1379),
.B(n_1462),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1419),
.B(n_1210),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1489),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1522),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1416),
.A2(n_1267),
.B(n_1246),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1371),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1464),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1533),
.B(n_1205),
.C(n_1186),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1399),
.B(n_1361),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1528),
.B(n_1196),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1561),
.A2(n_1303),
.B1(n_1343),
.B2(n_1367),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1412),
.A2(n_1280),
.B1(n_1300),
.B2(n_1299),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1471),
.B(n_1304),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1395),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1522),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1373),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1375),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1444),
.A2(n_1248),
.B1(n_1290),
.B2(n_1287),
.Y(n_1606)
);

NAND2xp33_ASAP7_75t_SL g1607 ( 
.A(n_1476),
.B(n_1282),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1444),
.A2(n_1248),
.B1(n_1287),
.B2(n_1318),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1398),
.A2(n_1362),
.B(n_1346),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1480),
.B(n_1308),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1425),
.B(n_1308),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1397),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1378),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1461),
.B(n_1317),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1402),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_SL g1616 ( 
.A(n_1443),
.B(n_1282),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1392),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1389),
.Y(n_1618)
);

NOR3xp33_ASAP7_75t_SL g1619 ( 
.A(n_1556),
.B(n_1546),
.C(n_1521),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1486),
.B(n_1317),
.Y(n_1620)
);

AND2x2_ASAP7_75t_SL g1621 ( 
.A(n_1527),
.B(n_1255),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1527),
.B(n_1282),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1477),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1449),
.A2(n_1354),
.B1(n_1265),
.B2(n_1331),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1433),
.B(n_1321),
.Y(n_1625)
);

NOR2x2_ASAP7_75t_L g1626 ( 
.A(n_1388),
.B(n_5),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1405),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1466),
.A2(n_1326),
.B1(n_1344),
.B2(n_1321),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1409),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1523),
.Y(n_1630)
);

OR2x6_ASAP7_75t_L g1631 ( 
.A(n_1432),
.B(n_1354),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1436),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1504),
.Y(n_1633)
);

BUFx4f_ASAP7_75t_SL g1634 ( 
.A(n_1523),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1432),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1530),
.B(n_1354),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1413),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1418),
.B(n_1326),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1415),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1404),
.B(n_1255),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1433),
.B(n_1344),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1497),
.A2(n_1356),
.B1(n_1331),
.B2(n_1332),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1501),
.B(n_1265),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1391),
.B(n_1531),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1467),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1479),
.A2(n_1356),
.B1(n_1357),
.B2(n_1332),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1389),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1542),
.B(n_1357),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1478),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1407),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1438),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1469),
.B(n_7),
.Y(n_1652)
);

NOR2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1422),
.B(n_382),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1417),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1414),
.Y(n_1655)
);

NOR2x2_ASAP7_75t_L g1656 ( 
.A(n_1388),
.B(n_8),
.Y(n_1656)
);

NOR2x2_ASAP7_75t_L g1657 ( 
.A(n_1388),
.B(n_9),
.Y(n_1657)
);

NAND2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1420),
.B(n_383),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1424),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1525),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1434),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1440),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1476),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1563),
.B(n_10),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1445),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1442),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1447),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1423),
.B(n_1460),
.Y(n_1668)
);

INVx4_ASAP7_75t_L g1669 ( 
.A(n_1434),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1473),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_R g1671 ( 
.A(n_1434),
.B(n_384),
.Y(n_1671)
);

NAND2x1p5_ASAP7_75t_L g1672 ( 
.A(n_1420),
.B(n_385),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1534),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_SL g1674 ( 
.A(n_1510),
.B(n_12),
.C(n_13),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1493),
.Y(n_1675)
);

BUFx4f_ASAP7_75t_L g1676 ( 
.A(n_1389),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1450),
.B(n_14),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_SL g1678 ( 
.A(n_1441),
.B(n_386),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1401),
.B(n_14),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1483),
.B(n_388),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1456),
.Y(n_1681)
);

BUFx4f_ASAP7_75t_L g1682 ( 
.A(n_1456),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1572),
.B(n_15),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1509),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1456),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1498),
.B(n_16),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1384),
.B(n_390),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1380),
.B(n_538),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1516),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1453),
.B(n_17),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1483),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1487),
.B(n_17),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1483),
.B(n_391),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1439),
.B(n_392),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1453),
.B(n_18),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1484),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1454),
.B(n_18),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1511),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1455),
.B(n_19),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1517),
.Y(n_1700)
);

INVx5_ASAP7_75t_L g1701 ( 
.A(n_1491),
.Y(n_1701)
);

CKINVDCx8_ASAP7_75t_R g1702 ( 
.A(n_1372),
.Y(n_1702)
);

BUFx12f_ASAP7_75t_L g1703 ( 
.A(n_1502),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1535),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1503),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1494),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1539),
.A2(n_1540),
.B1(n_1448),
.B2(n_1475),
.Y(n_1707)
);

AND2x6_ASAP7_75t_SL g1708 ( 
.A(n_1435),
.B(n_19),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1455),
.B(n_20),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1503),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1472),
.B(n_20),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1513),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1472),
.B(n_21),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1512),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1482),
.B(n_23),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1513),
.Y(n_1716)
);

AND2x6_ASAP7_75t_SL g1717 ( 
.A(n_1451),
.B(n_24),
.Y(n_1717)
);

OAI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1429),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1529),
.B(n_26),
.Y(n_1719)
);

OR2x6_ASAP7_75t_L g1720 ( 
.A(n_1491),
.B(n_393),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1437),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1406),
.B(n_394),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1524),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1502),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1502),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1482),
.B(n_27),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1545),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_SL g1728 ( 
.A(n_1520),
.B(n_28),
.C(n_29),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1548),
.B(n_537),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1430),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1558),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1564),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1492),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1430),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1377),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1550),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1507),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1459),
.B(n_34),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1452),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1385),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1385),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1369),
.B(n_35),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1566),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1537),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1386),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1386),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1518),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1518),
.Y(n_1748)
);

INVx5_ASAP7_75t_L g1749 ( 
.A(n_1507),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1390),
.B(n_37),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1551),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_SL g1752 ( 
.A(n_1376),
.B(n_395),
.Y(n_1752)
);

OR2x4_ASAP7_75t_L g1753 ( 
.A(n_1507),
.B(n_37),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1368),
.Y(n_1754)
);

NOR3xp33_ASAP7_75t_L g1755 ( 
.A(n_1515),
.B(n_38),
.C(n_39),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1368),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1500),
.B(n_38),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1463),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_R g1759 ( 
.A(n_1526),
.B(n_396),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1421),
.B(n_1426),
.Y(n_1760)
);

NOR3xp33_ASAP7_75t_SL g1761 ( 
.A(n_1532),
.B(n_40),
.C(n_41),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_SL g1762 ( 
.A(n_1396),
.B(n_40),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1400),
.B(n_42),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1744),
.B(n_1644),
.Y(n_1764)
);

NAND2xp33_ASAP7_75t_R g1765 ( 
.A(n_1759),
.B(n_1553),
.Y(n_1765)
);

NAND2xp33_ASAP7_75t_SL g1766 ( 
.A(n_1619),
.B(n_1403),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1664),
.B(n_1393),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1611),
.B(n_1541),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1707),
.B(n_1408),
.Y(n_1769)
);

NAND2xp33_ASAP7_75t_SL g1770 ( 
.A(n_1592),
.B(n_1554),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1730),
.B(n_1544),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1734),
.B(n_1554),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1683),
.B(n_1496),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1652),
.B(n_1589),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1621),
.B(n_1553),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1705),
.B(n_1538),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1710),
.B(n_1458),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1712),
.B(n_1370),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1716),
.B(n_1568),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1760),
.B(n_1570),
.Y(n_1781)
);

NAND2xp33_ASAP7_75t_SL g1782 ( 
.A(n_1592),
.B(n_1468),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1648),
.B(n_1410),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1668),
.B(n_1543),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1640),
.B(n_1488),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1736),
.B(n_1505),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_SL g1788 ( 
.A(n_1592),
.B(n_1470),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1694),
.B(n_1551),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1694),
.B(n_1481),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1686),
.B(n_1411),
.Y(n_1791)
);

NAND2xp33_ASAP7_75t_SL g1792 ( 
.A(n_1588),
.B(n_1565),
.Y(n_1792)
);

NAND2xp33_ASAP7_75t_SL g1793 ( 
.A(n_1596),
.B(n_1463),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1573),
.B(n_1427),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1747),
.B(n_1505),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1748),
.B(n_1519),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1638),
.B(n_1616),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1643),
.B(n_1427),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1692),
.B(n_1519),
.Y(n_1799)
);

NAND2xp33_ASAP7_75t_SL g1800 ( 
.A(n_1671),
.B(n_1474),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1595),
.B(n_1387),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1636),
.B(n_1394),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1577),
.B(n_1499),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1597),
.B(n_1536),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1757),
.B(n_1474),
.Y(n_1805)
);

NAND2xp33_ASAP7_75t_SL g1806 ( 
.A(n_1761),
.B(n_1490),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1687),
.B(n_1490),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1687),
.B(n_1506),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1598),
.B(n_1506),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1688),
.B(n_1514),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1740),
.B(n_1569),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1688),
.B(n_1514),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1741),
.B(n_1552),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1745),
.B(n_1552),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1746),
.B(n_1620),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1729),
.B(n_1571),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1729),
.B(n_1571),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1614),
.B(n_1446),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1610),
.B(n_1562),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1624),
.B(n_1549),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1598),
.B(n_1557),
.Y(n_1821)
);

NAND2xp33_ASAP7_75t_SL g1822 ( 
.A(n_1586),
.B(n_1559),
.Y(n_1822)
);

NAND2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1632),
.B(n_1560),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1624),
.B(n_43),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1677),
.B(n_43),
.Y(n_1825)
);

NAND2xp33_ASAP7_75t_SL g1826 ( 
.A(n_1669),
.B(n_44),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1751),
.B(n_44),
.Y(n_1827)
);

NAND2x1p5_ASAP7_75t_L g1828 ( 
.A(n_1635),
.B(n_398),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1585),
.B(n_400),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_SL g1830 ( 
.A(n_1690),
.B(n_45),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1585),
.B(n_402),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1695),
.B(n_46),
.Y(n_1832)
);

NAND2xp33_ASAP7_75t_SL g1833 ( 
.A(n_1669),
.B(n_46),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1699),
.B(n_47),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1603),
.B(n_403),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1709),
.B(n_1711),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1706),
.B(n_48),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1590),
.B(n_48),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1575),
.B(n_49),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1713),
.B(n_49),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1715),
.B(n_50),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1726),
.B(n_50),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1663),
.B(n_51),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1593),
.B(n_52),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1593),
.B(n_1719),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1721),
.B(n_53),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1697),
.B(n_1609),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1635),
.B(n_404),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1739),
.B(n_53),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1678),
.B(n_54),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1574),
.B(n_54),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1635),
.B(n_405),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1750),
.B(n_55),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1722),
.B(n_56),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1679),
.B(n_56),
.Y(n_1855)
);

NAND2xp33_ASAP7_75t_SL g1856 ( 
.A(n_1630),
.B(n_57),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1755),
.B(n_57),
.Y(n_1857)
);

NAND2xp33_ASAP7_75t_SL g1858 ( 
.A(n_1653),
.B(n_58),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1625),
.B(n_58),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1641),
.B(n_59),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1622),
.B(n_59),
.Y(n_1861)
);

NAND2xp33_ASAP7_75t_SL g1862 ( 
.A(n_1653),
.B(n_60),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1738),
.B(n_62),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_SL g1864 ( 
.A(n_1731),
.B(n_62),
.Y(n_1864)
);

NAND2xp33_ASAP7_75t_SL g1865 ( 
.A(n_1584),
.B(n_63),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1732),
.B(n_64),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1743),
.B(n_65),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1594),
.B(n_65),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1763),
.B(n_66),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_SL g1870 ( 
.A(n_1689),
.B(n_66),
.Y(n_1870)
);

NAND2xp33_ASAP7_75t_SL g1871 ( 
.A(n_1579),
.B(n_67),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_SL g1872 ( 
.A(n_1700),
.B(n_68),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1604),
.B(n_68),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1704),
.B(n_69),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1582),
.B(n_69),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1580),
.B(n_1576),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1580),
.B(n_70),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1602),
.B(n_70),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1605),
.B(n_71),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1670),
.B(n_71),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1612),
.B(n_73),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1615),
.B(n_74),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1613),
.B(n_75),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1627),
.B(n_75),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1629),
.B(n_76),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1633),
.B(n_76),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1637),
.B(n_77),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1578),
.B(n_78),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1639),
.B(n_78),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1654),
.B(n_79),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1659),
.B(n_81),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1666),
.B(n_81),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1583),
.B(n_83),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1714),
.B(n_1696),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1587),
.B(n_1591),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1701),
.B(n_406),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1698),
.B(n_84),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1714),
.B(n_84),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1723),
.B(n_85),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1727),
.B(n_85),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_SL g1901 ( 
.A(n_1646),
.B(n_86),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1762),
.B(n_86),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1733),
.B(n_88),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1733),
.B(n_90),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1617),
.B(n_90),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1752),
.B(n_91),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1623),
.B(n_92),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1649),
.B(n_93),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1675),
.B(n_94),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1684),
.B(n_1718),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1701),
.B(n_94),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_SL g1912 ( 
.A(n_1661),
.B(n_1691),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1650),
.B(n_95),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1655),
.B(n_95),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1701),
.B(n_96),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1608),
.B(n_96),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1608),
.B(n_1599),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_SL g1918 ( 
.A(n_1606),
.B(n_97),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1651),
.B(n_97),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1606),
.B(n_1660),
.Y(n_1920)
);

NAND2xp33_ASAP7_75t_SL g1921 ( 
.A(n_1691),
.B(n_98),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1742),
.B(n_101),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1581),
.B(n_101),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1662),
.B(n_102),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1665),
.B(n_1667),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1600),
.B(n_1607),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1735),
.B(n_103),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1618),
.B(n_104),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1895),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1925),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1814),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1809),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1847),
.B(n_1735),
.Y(n_1933)
);

O2A1O1Ixp33_ASAP7_75t_L g1934 ( 
.A1(n_1857),
.A2(n_1927),
.B(n_1825),
.C(n_1898),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1785),
.Y(n_1935)
);

BUFx12f_ASAP7_75t_L g1936 ( 
.A(n_1835),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1821),
.Y(n_1937)
);

A2O1A1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1858),
.A2(n_1862),
.B(n_1927),
.C(n_1766),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1785),
.Y(n_1939)
);

AND3x1_ASAP7_75t_SL g1940 ( 
.A(n_1843),
.B(n_1702),
.C(n_1708),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1815),
.Y(n_1941)
);

AO22x1_ASAP7_75t_L g1942 ( 
.A1(n_1903),
.A2(n_1904),
.B1(n_1852),
.B2(n_1896),
.Y(n_1942)
);

BUFx8_ASAP7_75t_SL g1943 ( 
.A(n_1767),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1764),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1835),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1848),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1827),
.Y(n_1947)
);

O2A1O1Ixp33_ASAP7_75t_SL g1948 ( 
.A1(n_1854),
.A2(n_1728),
.B(n_1674),
.C(n_1725),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1876),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1765),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1829),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_R g1952 ( 
.A(n_1765),
.B(n_1634),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1829),
.B(n_1720),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1831),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1888),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1774),
.B(n_1647),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1831),
.Y(n_1957)
);

INVx2_ASAP7_75t_SL g1958 ( 
.A(n_1848),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1852),
.B(n_1720),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1771),
.B(n_1658),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1778),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1896),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1807),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1800),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1797),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1811),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1768),
.B(n_1645),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1808),
.Y(n_1968)
);

BUFx3_ASAP7_75t_L g1969 ( 
.A(n_1880),
.Y(n_1969)
);

NOR2x1_ASAP7_75t_L g1970 ( 
.A(n_1775),
.B(n_1720),
.Y(n_1970)
);

BUFx3_ASAP7_75t_L g1971 ( 
.A(n_1899),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1913),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1772),
.B(n_1673),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1897),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1801),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1845),
.B(n_1754),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_1810),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1856),
.Y(n_1978)
);

AOI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1770),
.A2(n_1693),
.B(n_1680),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1914),
.Y(n_1980)
);

AO221x1_ASAP7_75t_L g1981 ( 
.A1(n_1824),
.A2(n_1685),
.B1(n_1681),
.B2(n_1618),
.C(n_1754),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1868),
.Y(n_1982)
);

AO32x2_ASAP7_75t_L g1983 ( 
.A1(n_1917),
.A2(n_1918),
.A3(n_1836),
.B1(n_1916),
.B2(n_1920),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1873),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1795),
.B(n_1758),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1879),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1900),
.Y(n_1987)
);

BUFx2_ASAP7_75t_L g1988 ( 
.A(n_1773),
.Y(n_1988)
);

INVxp67_ASAP7_75t_SL g1989 ( 
.A(n_1779),
.Y(n_1989)
);

AND2x2_ASAP7_75t_SL g1990 ( 
.A(n_1849),
.B(n_1676),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1813),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1828),
.Y(n_1992)
);

BUFx3_ASAP7_75t_L g1993 ( 
.A(n_1886),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1912),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1883),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1917),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1804),
.Y(n_1997)
);

INVx4_ASAP7_75t_L g1998 ( 
.A(n_1828),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1893),
.B(n_1753),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1877),
.A2(n_1693),
.B1(n_1628),
.B2(n_1672),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1812),
.B(n_1724),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1919),
.B(n_1799),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1796),
.B(n_1758),
.Y(n_2003)
);

INVx5_ASAP7_75t_L g2004 ( 
.A(n_1782),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1837),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1844),
.B(n_1749),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1816),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1859),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1793),
.Y(n_2009)
);

AOI21x1_ASAP7_75t_L g2010 ( 
.A1(n_1784),
.A2(n_1631),
.B(n_1642),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1905),
.Y(n_2011)
);

BUFx12f_ASAP7_75t_L g2012 ( 
.A(n_1865),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1817),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1908),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1839),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1781),
.B(n_1708),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1787),
.B(n_1749),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1803),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1894),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1822),
.Y(n_2020)
);

INVx3_ASAP7_75t_L g2021 ( 
.A(n_1902),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1805),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1918),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1769),
.B(n_1676),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1802),
.Y(n_2025)
);

CKINVDCx20_ASAP7_75t_R g2026 ( 
.A(n_1871),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1846),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1855),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1916),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1853),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1841),
.B(n_1756),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1789),
.B(n_1749),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_1911),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1926),
.B(n_1682),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1851),
.B(n_1717),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1777),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1869),
.B(n_1717),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1819),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1790),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1823),
.Y(n_2040)
);

INVx2_ASAP7_75t_SL g2041 ( 
.A(n_1915),
.Y(n_2041)
);

A2O1A1Ixp33_ASAP7_75t_L g2042 ( 
.A1(n_1791),
.A2(n_1682),
.B(n_1737),
.C(n_1626),
.Y(n_2042)
);

A2O1A1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_1920),
.A2(n_1656),
.B(n_1657),
.C(n_1756),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1860),
.Y(n_2044)
);

INVx5_ASAP7_75t_L g2045 ( 
.A(n_1788),
.Y(n_2045)
);

INVx2_ASAP7_75t_SL g2046 ( 
.A(n_1863),
.Y(n_2046)
);

AO22x1_ASAP7_75t_L g2047 ( 
.A1(n_1826),
.A2(n_1756),
.B1(n_1681),
.B2(n_1685),
.Y(n_2047)
);

OAI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1938),
.A2(n_1850),
.B(n_1906),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1929),
.Y(n_2049)
);

INVx2_ASAP7_75t_SL g2050 ( 
.A(n_1936),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1961),
.B(n_1776),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1979),
.A2(n_1960),
.B(n_1970),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1930),
.Y(n_2053)
);

O2A1O1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_1934),
.A2(n_1922),
.B(n_1830),
.C(n_1834),
.Y(n_2054)
);

OAI21x1_ASAP7_75t_L g2055 ( 
.A1(n_2010),
.A2(n_1794),
.B(n_1818),
.Y(n_2055)
);

OAI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1950),
.A2(n_1922),
.B1(n_1901),
.B2(n_1875),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1935),
.Y(n_2057)
);

AO21x2_ASAP7_75t_L g2058 ( 
.A1(n_1989),
.A2(n_1820),
.B(n_1786),
.Y(n_2058)
);

OR2x6_ASAP7_75t_L g2059 ( 
.A(n_1979),
.B(n_1910),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1934),
.A2(n_1780),
.B(n_1832),
.Y(n_2060)
);

BUFx8_ASAP7_75t_L g2061 ( 
.A(n_2012),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2043),
.A2(n_1840),
.B1(n_1842),
.B2(n_1923),
.Y(n_2062)
);

BUFx6f_ASAP7_75t_L g2063 ( 
.A(n_1962),
.Y(n_2063)
);

INVx6_ASAP7_75t_L g2064 ( 
.A(n_1962),
.Y(n_2064)
);

O2A1O1Ixp33_ASAP7_75t_L g2065 ( 
.A1(n_2016),
.A2(n_1861),
.B(n_1909),
.C(n_1907),
.Y(n_2065)
);

INVx5_ASAP7_75t_L g2066 ( 
.A(n_2020),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1970),
.A2(n_1798),
.B(n_1783),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_2000),
.A2(n_1792),
.B(n_1921),
.Y(n_2068)
);

OAI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_2009),
.A2(n_1924),
.B1(n_1872),
.B2(n_1874),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1939),
.B(n_1618),
.Y(n_2070)
);

BUFx2_ASAP7_75t_SL g2071 ( 
.A(n_1969),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1941),
.Y(n_2072)
);

INVx5_ASAP7_75t_L g2073 ( 
.A(n_2004),
.Y(n_2073)
);

INVx3_ASAP7_75t_SL g2074 ( 
.A(n_1978),
.Y(n_2074)
);

AO32x2_ASAP7_75t_L g2075 ( 
.A1(n_2005),
.A2(n_2027),
.A3(n_2046),
.B1(n_2033),
.B2(n_2041),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1996),
.Y(n_2076)
);

AOI221x1_ASAP7_75t_L g2077 ( 
.A1(n_2035),
.A2(n_1806),
.B1(n_1838),
.B2(n_1928),
.C(n_1833),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1996),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_1988),
.Y(n_2079)
);

OAI21xp5_ASAP7_75t_L g2080 ( 
.A1(n_1989),
.A2(n_1866),
.B(n_1864),
.Y(n_2080)
);

AND2x6_ASAP7_75t_L g2081 ( 
.A(n_1953),
.B(n_1681),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1933),
.A2(n_1867),
.B(n_1870),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_SL g2083 ( 
.A1(n_1959),
.A2(n_1881),
.B(n_1878),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2004),
.A2(n_1884),
.B(n_1882),
.Y(n_2084)
);

NAND3x1_ASAP7_75t_L g2085 ( 
.A(n_2037),
.B(n_104),
.C(n_105),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1999),
.A2(n_1887),
.B1(n_1889),
.B2(n_1885),
.Y(n_2086)
);

INVxp67_ASAP7_75t_L g2087 ( 
.A(n_1967),
.Y(n_2087)
);

NOR2x1_ASAP7_75t_R g2088 ( 
.A(n_1993),
.B(n_1703),
.Y(n_2088)
);

AO31x2_ASAP7_75t_L g2089 ( 
.A1(n_1998),
.A2(n_1949),
.A3(n_2029),
.B(n_2023),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1966),
.B(n_1890),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2004),
.A2(n_1892),
.B(n_1891),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1965),
.Y(n_2092)
);

OAI21x1_ASAP7_75t_L g2093 ( 
.A1(n_1976),
.A2(n_1631),
.B(n_1685),
.Y(n_2093)
);

A2O1A1Ixp33_ASAP7_75t_L g2094 ( 
.A1(n_1933),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_1976),
.A2(n_409),
.B(n_407),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_SL g2096 ( 
.A(n_2045),
.B(n_410),
.Y(n_2096)
);

AOI21xp5_ASAP7_75t_L g2097 ( 
.A1(n_2045),
.A2(n_1953),
.B(n_1959),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_SL g2098 ( 
.A(n_2045),
.B(n_412),
.Y(n_2098)
);

O2A1O1Ixp33_ASAP7_75t_SL g2099 ( 
.A1(n_2042),
.A2(n_110),
.B(n_106),
.C(n_109),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2039),
.A2(n_1975),
.B1(n_1990),
.B2(n_2024),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2047),
.A2(n_1948),
.B(n_2034),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2026),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_2102)
);

AO31x2_ASAP7_75t_L g2103 ( 
.A1(n_2036),
.A2(n_114),
.A3(n_112),
.B(n_113),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_1935),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_2031),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_1985),
.A2(n_414),
.B(n_413),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2019),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_1985),
.A2(n_416),
.B(n_415),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_2039),
.A2(n_116),
.B1(n_113),
.B2(n_115),
.Y(n_2109)
);

AOI221xp5_ASAP7_75t_SL g2110 ( 
.A1(n_1944),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.C(n_118),
.Y(n_2110)
);

BUFx10_ASAP7_75t_L g2111 ( 
.A(n_2028),
.Y(n_2111)
);

O2A1O1Ixp5_ASAP7_75t_SL g2112 ( 
.A1(n_2044),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_2112)
);

INVx2_ASAP7_75t_SL g2113 ( 
.A(n_1971),
.Y(n_2113)
);

OA21x2_ASAP7_75t_L g2114 ( 
.A1(n_1981),
.A2(n_119),
.B(n_121),
.Y(n_2114)
);

AOI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_2002),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2092),
.B(n_1937),
.Y(n_2116)
);

OAI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2068),
.A2(n_2015),
.B(n_2040),
.Y(n_2117)
);

BUFx2_ASAP7_75t_R g2118 ( 
.A(n_2074),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2053),
.Y(n_2119)
);

AND2x2_ASAP7_75t_SL g2120 ( 
.A(n_2096),
.B(n_2002),
.Y(n_2120)
);

OA21x2_ASAP7_75t_L g2121 ( 
.A1(n_2055),
.A2(n_2017),
.B(n_2003),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_2056),
.A2(n_2021),
.B1(n_2008),
.B2(n_1947),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2076),
.Y(n_2123)
);

OA21x2_ASAP7_75t_L g2124 ( 
.A1(n_2052),
.A2(n_2017),
.B(n_2003),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2072),
.B(n_1944),
.Y(n_2125)
);

AO21x2_ASAP7_75t_L g2126 ( 
.A1(n_2067),
.A2(n_1952),
.B(n_2022),
.Y(n_2126)
);

OAI21x1_ASAP7_75t_L g2127 ( 
.A1(n_2106),
.A2(n_2108),
.B(n_2097),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_2095),
.A2(n_2018),
.B(n_2038),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2078),
.Y(n_2129)
);

NOR2xp33_ASAP7_75t_L g2130 ( 
.A(n_2059),
.B(n_2039),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_2098),
.A2(n_1942),
.B(n_1973),
.Y(n_2131)
);

AO32x2_ASAP7_75t_L g2132 ( 
.A1(n_2062),
.A2(n_1983),
.A3(n_1958),
.B1(n_2021),
.B2(n_2030),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_2093),
.A2(n_2107),
.B(n_2101),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2089),
.Y(n_2134)
);

INVxp67_ASAP7_75t_L g2135 ( 
.A(n_2071),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_2112),
.A2(n_1992),
.B(n_2025),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2089),
.Y(n_2137)
);

AO21x1_ASAP7_75t_L g2138 ( 
.A1(n_2060),
.A2(n_1972),
.B(n_1955),
.Y(n_2138)
);

OAI21xp5_ASAP7_75t_L g2139 ( 
.A1(n_2054),
.A2(n_1973),
.B(n_1980),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2079),
.B(n_1956),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2049),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2075),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_2073),
.B(n_1935),
.Y(n_2143)
);

OA21x2_ASAP7_75t_L g2144 ( 
.A1(n_2080),
.A2(n_2006),
.B(n_1991),
.Y(n_2144)
);

AOI21xp33_ASAP7_75t_L g2145 ( 
.A1(n_2065),
.A2(n_2059),
.B(n_2048),
.Y(n_2145)
);

AOI221xp5_ASAP7_75t_L g2146 ( 
.A1(n_2099),
.A2(n_1986),
.B1(n_1995),
.B2(n_1984),
.C(n_1982),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2115),
.A2(n_2085),
.B1(n_2094),
.B2(n_2100),
.Y(n_2147)
);

INVx1_ASAP7_75t_SL g2148 ( 
.A(n_2113),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2075),
.Y(n_2149)
);

OAI22xp33_ASAP7_75t_L g2150 ( 
.A1(n_2077),
.A2(n_2102),
.B1(n_2086),
.B2(n_2066),
.Y(n_2150)
);

OAI21x1_ASAP7_75t_L g2151 ( 
.A1(n_2112),
.A2(n_1992),
.B(n_1997),
.Y(n_2151)
);

OA21x2_ASAP7_75t_L g2152 ( 
.A1(n_2084),
.A2(n_2006),
.B(n_1994),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2105),
.B(n_2011),
.Y(n_2153)
);

OAI21x1_ASAP7_75t_L g2154 ( 
.A1(n_2051),
.A2(n_2091),
.B(n_2090),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_2111),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2087),
.B(n_1932),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_2069),
.A2(n_2014),
.B1(n_1974),
.B2(n_1987),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2058),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_2082),
.A2(n_1954),
.B1(n_1957),
.B2(n_1951),
.Y(n_2159)
);

OAI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_2147),
.A2(n_2066),
.B1(n_2073),
.B2(n_1963),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2140),
.B(n_2057),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2150),
.A2(n_2110),
.B1(n_1946),
.B2(n_1957),
.Y(n_2162)
);

CKINVDCx6p67_ASAP7_75t_R g2163 ( 
.A(n_2120),
.Y(n_2163)
);

AOI21xp33_ASAP7_75t_L g2164 ( 
.A1(n_2126),
.A2(n_2088),
.B(n_2114),
.Y(n_2164)
);

OAI221xp5_ASAP7_75t_L g2165 ( 
.A1(n_2145),
.A2(n_2109),
.B1(n_2083),
.B2(n_2050),
.C(n_1964),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_2124),
.Y(n_2166)
);

AOI22xp33_ASAP7_75t_L g2167 ( 
.A1(n_2122),
.A2(n_2114),
.B1(n_1951),
.B2(n_1957),
.Y(n_2167)
);

OAI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2122),
.A2(n_2073),
.B1(n_1946),
.B2(n_1968),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_2143),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_2120),
.A2(n_1951),
.B1(n_1968),
.B2(n_1963),
.Y(n_2170)
);

AOI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_2139),
.A2(n_1963),
.B1(n_1977),
.B2(n_1968),
.Y(n_2171)
);

CKINVDCx16_ASAP7_75t_R g2172 ( 
.A(n_2156),
.Y(n_2172)
);

NAND2x1p5_ASAP7_75t_L g2173 ( 
.A(n_2152),
.B(n_2124),
.Y(n_2173)
);

AOI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_2157),
.A2(n_1977),
.B1(n_2013),
.B2(n_2007),
.Y(n_2174)
);

OAI21x1_ASAP7_75t_L g2175 ( 
.A1(n_2127),
.A2(n_2104),
.B(n_1931),
.Y(n_2175)
);

HB1xp67_ASAP7_75t_L g2176 ( 
.A(n_2124),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2119),
.Y(n_2177)
);

INVx4_ASAP7_75t_L g2178 ( 
.A(n_2155),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_2116),
.B(n_2070),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2123),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_R g2181 ( 
.A(n_2155),
.B(n_2061),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2129),
.Y(n_2182)
);

CKINVDCx20_ASAP7_75t_R g2183 ( 
.A(n_2148),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_2118),
.Y(n_2184)
);

AND2x4_ASAP7_75t_L g2185 ( 
.A(n_2133),
.B(n_2063),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_2154),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_2169),
.Y(n_2187)
);

BUFx3_ASAP7_75t_L g2188 ( 
.A(n_2183),
.Y(n_2188)
);

OAI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2163),
.A2(n_2159),
.B1(n_2157),
.B2(n_2131),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2160),
.A2(n_2117),
.B1(n_2138),
.B2(n_2146),
.Y(n_2190)
);

AOI222xp33_ASAP7_75t_L g2191 ( 
.A1(n_2165),
.A2(n_2149),
.B1(n_2153),
.B2(n_2135),
.C1(n_2142),
.C2(n_2159),
.Y(n_2191)
);

INVx1_ASAP7_75t_SL g2192 ( 
.A(n_2181),
.Y(n_2192)
);

OA21x2_ASAP7_75t_L g2193 ( 
.A1(n_2166),
.A2(n_2137),
.B(n_2134),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2182),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2182),
.Y(n_2195)
);

AOI21xp5_ASAP7_75t_L g2196 ( 
.A1(n_2164),
.A2(n_2126),
.B(n_2168),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2180),
.B(n_2154),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_2187),
.B(n_2178),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_R g2199 ( 
.A(n_2192),
.B(n_2184),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_R g2200 ( 
.A(n_2188),
.B(n_2155),
.Y(n_2200)
);

XNOR2xp5_ASAP7_75t_L g2201 ( 
.A(n_2189),
.B(n_1940),
.Y(n_2201)
);

CKINVDCx20_ASAP7_75t_R g2202 ( 
.A(n_2190),
.Y(n_2202)
);

INVxp67_ASAP7_75t_L g2203 ( 
.A(n_2191),
.Y(n_2203)
);

XNOR2xp5_ASAP7_75t_L g2204 ( 
.A(n_2190),
.B(n_2162),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2198),
.B(n_2187),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2198),
.B(n_2187),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_2201),
.Y(n_2207)
);

INVxp67_ASAP7_75t_SL g2208 ( 
.A(n_2204),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2202),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2203),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2200),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2199),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2198),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2198),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2209),
.B(n_2208),
.Y(n_2215)
);

NAND4xp25_ASAP7_75t_L g2216 ( 
.A(n_2210),
.B(n_2207),
.C(n_2209),
.D(n_2211),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2205),
.B(n_2172),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2210),
.B(n_2196),
.Y(n_2218)
);

OAI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2211),
.A2(n_2170),
.B1(n_2167),
.B2(n_2171),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2205),
.B(n_2181),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2206),
.B(n_2169),
.Y(n_2221)
);

OAI21xp33_ASAP7_75t_L g2222 ( 
.A1(n_2213),
.A2(n_2197),
.B(n_2171),
.Y(n_2222)
);

NAND3xp33_ASAP7_75t_L g2223 ( 
.A(n_2213),
.B(n_2186),
.C(n_2167),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2214),
.B(n_2194),
.Y(n_2224)
);

NAND3xp33_ASAP7_75t_SL g2225 ( 
.A(n_2212),
.B(n_2173),
.C(n_2170),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2220),
.B(n_2212),
.Y(n_2226)
);

OA211x2_ASAP7_75t_L g2227 ( 
.A1(n_2225),
.A2(n_2215),
.B(n_2218),
.C(n_2222),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2217),
.B(n_2206),
.Y(n_2228)
);

AOI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_2216),
.A2(n_2207),
.B1(n_2214),
.B2(n_2176),
.C(n_2173),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_2221),
.Y(n_2230)
);

INVxp67_ASAP7_75t_SL g2231 ( 
.A(n_2223),
.Y(n_2231)
);

AOI221xp5_ASAP7_75t_L g2232 ( 
.A1(n_2219),
.A2(n_2174),
.B1(n_2142),
.B2(n_2158),
.C(n_2195),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2224),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_2220),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2228),
.B(n_2178),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2226),
.B(n_2169),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2234),
.B(n_2230),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_2234),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2237),
.B(n_2231),
.Y(n_2239)
);

OAI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2238),
.A2(n_2229),
.B(n_2232),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2238),
.B(n_2233),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2236),
.B(n_2229),
.Y(n_2242)
);

OAI22xp5_ASAP7_75t_SL g2243 ( 
.A1(n_2240),
.A2(n_2227),
.B1(n_1943),
.B2(n_2232),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_R g2244 ( 
.A(n_2239),
.B(n_2235),
.Y(n_2244)
);

NOR2x1_ASAP7_75t_SL g2245 ( 
.A(n_2241),
.B(n_2169),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_2242),
.B(n_2161),
.Y(n_2246)
);

OAI221xp5_ASAP7_75t_L g2247 ( 
.A1(n_2240),
.A2(n_2174),
.B1(n_2130),
.B2(n_2152),
.C(n_1945),
.Y(n_2247)
);

AO221x2_ASAP7_75t_L g2248 ( 
.A1(n_2241),
.A2(n_2158),
.B1(n_2177),
.B2(n_2125),
.C(n_2141),
.Y(n_2248)
);

NAND4xp25_ASAP7_75t_L g2249 ( 
.A(n_2246),
.B(n_2130),
.C(n_2185),
.D(n_2143),
.Y(n_2249)
);

OAI21xp33_ASAP7_75t_L g2250 ( 
.A1(n_2244),
.A2(n_2185),
.B(n_2133),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2245),
.B(n_2248),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_2243),
.B(n_2179),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2247),
.B(n_2179),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2246),
.Y(n_2254)
);

OAI32xp33_ASAP7_75t_L g2255 ( 
.A1(n_2246),
.A2(n_2132),
.A3(n_2193),
.B1(n_2103),
.B2(n_1983),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2246),
.Y(n_2256)
);

NOR2xp67_ASAP7_75t_L g2257 ( 
.A(n_2246),
.B(n_122),
.Y(n_2257)
);

OR2x6_ASAP7_75t_L g2258 ( 
.A(n_2243),
.B(n_1962),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2257),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2254),
.Y(n_2260)
);

AOI21xp33_ASAP7_75t_SL g2261 ( 
.A1(n_2256),
.A2(n_123),
.B(n_124),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2251),
.Y(n_2262)
);

OR2x2_ASAP7_75t_L g2263 ( 
.A(n_2249),
.B(n_2193),
.Y(n_2263)
);

O2A1O1Ixp33_ASAP7_75t_SL g2264 ( 
.A1(n_2255),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2252),
.B(n_2152),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2253),
.B(n_2185),
.Y(n_2266)
);

AND2x4_ASAP7_75t_L g2267 ( 
.A(n_2258),
.B(n_2116),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2258),
.B(n_2116),
.Y(n_2268)
);

A2O1A1Ixp33_ASAP7_75t_L g2269 ( 
.A1(n_2250),
.A2(n_2127),
.B(n_2175),
.C(n_2136),
.Y(n_2269)
);

OR2x2_ASAP7_75t_L g2270 ( 
.A(n_2254),
.B(n_2144),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_2252),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2271),
.B(n_125),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2262),
.A2(n_2144),
.B1(n_2064),
.B2(n_2143),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2259),
.B(n_2132),
.Y(n_2274)
);

AOI222xp33_ASAP7_75t_L g2275 ( 
.A1(n_2260),
.A2(n_2136),
.B1(n_2151),
.B2(n_130),
.C1(n_132),
.C2(n_128),
.Y(n_2275)
);

INVxp67_ASAP7_75t_SL g2276 ( 
.A(n_2266),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2261),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2267),
.B(n_2132),
.Y(n_2278)
);

OAI221xp5_ASAP7_75t_L g2279 ( 
.A1(n_2263),
.A2(n_2144),
.B1(n_2064),
.B2(n_2121),
.C(n_2013),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2267),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2268),
.B(n_2132),
.Y(n_2281)
);

NAND3xp33_ASAP7_75t_L g2282 ( 
.A(n_2264),
.B(n_128),
.C(n_129),
.Y(n_2282)
);

AOI221xp5_ASAP7_75t_L g2283 ( 
.A1(n_2265),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.C(n_133),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2270),
.A2(n_1977),
.B1(n_2013),
.B2(n_2007),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_2269),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_2259),
.B(n_2063),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2280),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2272),
.B(n_131),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2277),
.B(n_134),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2282),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2276),
.Y(n_2291)
);

INVx1_ASAP7_75t_SL g2292 ( 
.A(n_2286),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2285),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2274),
.Y(n_2294)
);

OAI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2283),
.A2(n_2151),
.B(n_2128),
.Y(n_2295)
);

NOR2xp67_ASAP7_75t_L g2296 ( 
.A(n_2284),
.B(n_135),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2281),
.B(n_2278),
.Y(n_2297)
);

INVx1_ASAP7_75t_SL g2298 ( 
.A(n_2273),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_2275),
.A2(n_2081),
.B1(n_2001),
.B2(n_2121),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2279),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2287),
.A2(n_2081),
.B1(n_2001),
.B2(n_2121),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2289),
.Y(n_2302)
);

AOI222xp33_ASAP7_75t_L g2303 ( 
.A1(n_2293),
.A2(n_137),
.B1(n_140),
.B2(n_135),
.C1(n_136),
.C2(n_138),
.Y(n_2303)
);

INVx2_ASAP7_75t_SL g2304 ( 
.A(n_2291),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2290),
.Y(n_2305)
);

OAI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_2292),
.A2(n_2007),
.B1(n_2032),
.B2(n_2103),
.Y(n_2306)
);

NAND2x1_ASAP7_75t_L g2307 ( 
.A(n_2294),
.B(n_2081),
.Y(n_2307)
);

XNOR2xp5_ASAP7_75t_L g2308 ( 
.A(n_2297),
.B(n_136),
.Y(n_2308)
);

INVxp67_ASAP7_75t_SL g2309 ( 
.A(n_2296),
.Y(n_2309)
);

OAI32xp33_ASAP7_75t_L g2310 ( 
.A1(n_2298),
.A2(n_140),
.A3(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2288),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2300),
.Y(n_2312)
);

OAI21xp33_ASAP7_75t_SL g2313 ( 
.A1(n_2299),
.A2(n_2128),
.B(n_141),
.Y(n_2313)
);

OAI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2295),
.A2(n_142),
.B(n_143),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2287),
.B(n_143),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2287),
.Y(n_2316)
);

OAI322xp33_ASAP7_75t_L g2317 ( 
.A1(n_2293),
.A2(n_144),
.A3(n_145),
.B1(n_146),
.B2(n_148),
.C1(n_149),
.C2(n_151),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2287),
.B(n_144),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_2287),
.Y(n_2319)
);

XNOR2xp5_ASAP7_75t_L g2320 ( 
.A(n_2287),
.B(n_145),
.Y(n_2320)
);

INVx2_ASAP7_75t_SL g2321 ( 
.A(n_2287),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2289),
.A2(n_146),
.B(n_148),
.Y(n_2322)
);

INVxp67_ASAP7_75t_L g2323 ( 
.A(n_2315),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2320),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2308),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2319),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2318),
.Y(n_2327)
);

BUFx4f_ASAP7_75t_SL g2328 ( 
.A(n_2321),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2309),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2316),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2305),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2304),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2310),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2307),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2312),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2317),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2302),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2311),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2314),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2322),
.Y(n_2340)
);

INVxp67_ASAP7_75t_SL g2341 ( 
.A(n_2303),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2313),
.Y(n_2342)
);

INVxp33_ASAP7_75t_L g2343 ( 
.A(n_2301),
.Y(n_2343)
);

INVx1_ASAP7_75t_SL g2344 ( 
.A(n_2306),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2320),
.Y(n_2345)
);

CKINVDCx16_ASAP7_75t_R g2346 ( 
.A(n_2319),
.Y(n_2346)
);

INVxp33_ASAP7_75t_SL g2347 ( 
.A(n_2308),
.Y(n_2347)
);

INVx1_ASAP7_75t_SL g2348 ( 
.A(n_2320),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2320),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2319),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2320),
.Y(n_2351)
);

INVxp67_ASAP7_75t_SL g2352 ( 
.A(n_2320),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2320),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2320),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2319),
.B(n_149),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2320),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2319),
.B(n_151),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2320),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2320),
.Y(n_2359)
);

NAND5xp2_ASAP7_75t_L g2360 ( 
.A(n_2332),
.B(n_154),
.C(n_152),
.D(n_153),
.E(n_155),
.Y(n_2360)
);

AOI21xp33_ASAP7_75t_L g2361 ( 
.A1(n_2343),
.A2(n_153),
.B(n_154),
.Y(n_2361)
);

A2O1A1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_2357),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2362)
);

OAI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2341),
.A2(n_156),
.B(n_157),
.Y(n_2363)
);

OAI322xp33_ASAP7_75t_L g2364 ( 
.A1(n_2329),
.A2(n_160),
.A3(n_161),
.B1(n_162),
.B2(n_163),
.C1(n_164),
.C2(n_165),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2346),
.B(n_160),
.Y(n_2365)
);

OAI211xp5_ASAP7_75t_L g2366 ( 
.A1(n_2333),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_2366)
);

OAI321xp33_ASAP7_75t_L g2367 ( 
.A1(n_2336),
.A2(n_166),
.A3(n_168),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_2367)
);

OAI21xp33_ASAP7_75t_SL g2368 ( 
.A1(n_2342),
.A2(n_166),
.B(n_167),
.Y(n_2368)
);

INVx2_ASAP7_75t_SL g2369 ( 
.A(n_2328),
.Y(n_2369)
);

O2A1O1Ixp33_ASAP7_75t_L g2370 ( 
.A1(n_2355),
.A2(n_170),
.B(n_168),
.C(n_169),
.Y(n_2370)
);

O2A1O1Ixp33_ASAP7_75t_L g2371 ( 
.A1(n_2355),
.A2(n_2326),
.B(n_2350),
.C(n_2331),
.Y(n_2371)
);

AOI21xp33_ASAP7_75t_L g2372 ( 
.A1(n_2330),
.A2(n_169),
.B(n_170),
.Y(n_2372)
);

AOI21xp33_ASAP7_75t_L g2373 ( 
.A1(n_2335),
.A2(n_171),
.B(n_172),
.Y(n_2373)
);

XNOR2xp5_ASAP7_75t_L g2374 ( 
.A(n_2347),
.B(n_171),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_2334),
.Y(n_2375)
);

A2O1A1Ixp33_ASAP7_75t_L g2376 ( 
.A1(n_2344),
.A2(n_2352),
.B(n_2325),
.C(n_2348),
.Y(n_2376)
);

OAI311xp33_ASAP7_75t_L g2377 ( 
.A1(n_2340),
.A2(n_175),
.A3(n_173),
.B1(n_174),
.C1(n_177),
.Y(n_2377)
);

NOR3xp33_ASAP7_75t_L g2378 ( 
.A(n_2348),
.B(n_173),
.C(n_174),
.Y(n_2378)
);

INVxp67_ASAP7_75t_L g2379 ( 
.A(n_2339),
.Y(n_2379)
);

A2O1A1Ixp33_ASAP7_75t_L g2380 ( 
.A1(n_2344),
.A2(n_179),
.B(n_175),
.C(n_178),
.Y(n_2380)
);

INVx2_ASAP7_75t_SL g2381 ( 
.A(n_2324),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2345),
.A2(n_2032),
.B1(n_180),
.B2(n_178),
.Y(n_2382)
);

INVxp67_ASAP7_75t_L g2383 ( 
.A(n_2349),
.Y(n_2383)
);

AOI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_2338),
.A2(n_2337),
.B1(n_2353),
.B2(n_2351),
.Y(n_2384)
);

NAND4xp25_ASAP7_75t_L g2385 ( 
.A(n_2354),
.B(n_2358),
.C(n_2359),
.D(n_2356),
.Y(n_2385)
);

AOI22xp33_ASAP7_75t_L g2386 ( 
.A1(n_2327),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2386)
);

A2O1A1Ixp33_ASAP7_75t_L g2387 ( 
.A1(n_2323),
.A2(n_185),
.B(n_181),
.C(n_184),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2355),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2346),
.B(n_184),
.Y(n_2389)
);

OAI211xp5_ASAP7_75t_L g2390 ( 
.A1(n_2341),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2390)
);

NOR2xp67_ASAP7_75t_L g2391 ( 
.A(n_2355),
.B(n_186),
.Y(n_2391)
);

OAI211xp5_ASAP7_75t_L g2392 ( 
.A1(n_2368),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_2392)
);

OAI222xp33_ASAP7_75t_L g2393 ( 
.A1(n_2369),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.C1(n_192),
.C2(n_193),
.Y(n_2393)
);

AOI221xp5_ASAP7_75t_SL g2394 ( 
.A1(n_2376),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.C(n_197),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2381),
.A2(n_197),
.B1(n_194),
.B2(n_195),
.Y(n_2395)
);

AOI21xp5_ASAP7_75t_L g2396 ( 
.A1(n_2371),
.A2(n_198),
.B(n_199),
.Y(n_2396)
);

AOI221xp5_ASAP7_75t_L g2397 ( 
.A1(n_2380),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.C(n_201),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2374),
.Y(n_2398)
);

A2O1A1Ixp33_ASAP7_75t_SL g2399 ( 
.A1(n_2379),
.A2(n_203),
.B(n_200),
.C(n_202),
.Y(n_2399)
);

AOI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2363),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.C(n_205),
.Y(n_2400)
);

O2A1O1Ixp33_ASAP7_75t_L g2401 ( 
.A1(n_2377),
.A2(n_207),
.B(n_205),
.C(n_206),
.Y(n_2401)
);

NAND4xp25_ASAP7_75t_L g2402 ( 
.A(n_2384),
.B(n_208),
.C(n_206),
.D(n_207),
.Y(n_2402)
);

AOI221xp5_ASAP7_75t_SL g2403 ( 
.A1(n_2383),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.C(n_212),
.Y(n_2403)
);

OAI211xp5_ASAP7_75t_SL g2404 ( 
.A1(n_2388),
.A2(n_213),
.B(n_210),
.C(n_212),
.Y(n_2404)
);

NAND2xp33_ASAP7_75t_R g2405 ( 
.A(n_2375),
.B(n_213),
.Y(n_2405)
);

AO22x2_ASAP7_75t_L g2406 ( 
.A1(n_2365),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_2406)
);

OAI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2389),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_2407)
);

AOI31xp33_ASAP7_75t_L g2408 ( 
.A1(n_2390),
.A2(n_221),
.A3(n_219),
.B(n_220),
.Y(n_2408)
);

AOI211x1_ASAP7_75t_SL g2409 ( 
.A1(n_2385),
.A2(n_222),
.B(n_219),
.C(n_220),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2360),
.B(n_222),
.Y(n_2410)
);

AOI22xp33_ASAP7_75t_L g2411 ( 
.A1(n_2378),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2411)
);

NOR3xp33_ASAP7_75t_L g2412 ( 
.A(n_2367),
.B(n_223),
.C(n_224),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2391),
.Y(n_2413)
);

NAND5xp2_ASAP7_75t_L g2414 ( 
.A(n_2366),
.B(n_2370),
.C(n_2382),
.D(n_2361),
.E(n_2386),
.Y(n_2414)
);

OAI211xp5_ASAP7_75t_SL g2415 ( 
.A1(n_2372),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_2415)
);

AND4x1_ASAP7_75t_L g2416 ( 
.A(n_2362),
.B(n_228),
.C(n_226),
.D(n_227),
.Y(n_2416)
);

NOR2xp33_ASAP7_75t_L g2417 ( 
.A(n_2373),
.B(n_228),
.Y(n_2417)
);

OAI211xp5_ASAP7_75t_L g2418 ( 
.A1(n_2387),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_2418)
);

OAI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2364),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.C(n_233),
.Y(n_2419)
);

NAND3xp33_ASAP7_75t_L g2420 ( 
.A(n_2380),
.B(n_232),
.C(n_234),
.Y(n_2420)
);

NAND2xp33_ASAP7_75t_SL g2421 ( 
.A(n_2365),
.B(n_234),
.Y(n_2421)
);

AOI221xp5_ASAP7_75t_L g2422 ( 
.A1(n_2368),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.C(n_238),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2369),
.B(n_235),
.Y(n_2423)
);

NAND4xp25_ASAP7_75t_L g2424 ( 
.A(n_2384),
.B(n_238),
.C(n_236),
.D(n_237),
.Y(n_2424)
);

OAI221xp5_ASAP7_75t_L g2425 ( 
.A1(n_2368),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.C(n_242),
.Y(n_2425)
);

NAND4xp25_ASAP7_75t_L g2426 ( 
.A(n_2384),
.B(n_241),
.C(n_239),
.D(n_240),
.Y(n_2426)
);

O2A1O1Ixp33_ASAP7_75t_L g2427 ( 
.A1(n_2380),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_2427)
);

AOI222xp33_ASAP7_75t_L g2428 ( 
.A1(n_2375),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.C1(n_247),
.C2(n_248),
.Y(n_2428)
);

AOI221xp5_ASAP7_75t_L g2429 ( 
.A1(n_2368),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.C(n_249),
.Y(n_2429)
);

AOI211x1_ASAP7_75t_SL g2430 ( 
.A1(n_2376),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_2430)
);

OAI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_2376),
.A2(n_250),
.B(n_251),
.Y(n_2431)
);

O2A1O1Ixp33_ASAP7_75t_L g2432 ( 
.A1(n_2380),
.A2(n_256),
.B(n_252),
.C(n_253),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2374),
.Y(n_2433)
);

NAND4xp75_ASAP7_75t_L g2434 ( 
.A(n_2368),
.B(n_257),
.C(n_252),
.D(n_256),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2369),
.B(n_257),
.Y(n_2435)
);

OAI211xp5_ASAP7_75t_L g2436 ( 
.A1(n_2368),
.A2(n_260),
.B(n_258),
.C(n_259),
.Y(n_2436)
);

OAI221xp5_ASAP7_75t_L g2437 ( 
.A1(n_2368),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.C(n_263),
.Y(n_2437)
);

AOI221xp5_ASAP7_75t_L g2438 ( 
.A1(n_2368),
.A2(n_261),
.B1(n_262),
.B2(n_264),
.C(n_265),
.Y(n_2438)
);

BUFx3_ASAP7_75t_L g2439 ( 
.A(n_2375),
.Y(n_2439)
);

OAI211xp5_ASAP7_75t_SL g2440 ( 
.A1(n_2431),
.A2(n_2430),
.B(n_2413),
.C(n_2398),
.Y(n_2440)
);

OAI21xp5_ASAP7_75t_L g2441 ( 
.A1(n_2401),
.A2(n_265),
.B(n_266),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2434),
.Y(n_2442)
);

A2O1A1Ixp33_ASAP7_75t_L g2443 ( 
.A1(n_2427),
.A2(n_2432),
.B(n_2410),
.C(n_2396),
.Y(n_2443)
);

OAI211xp5_ASAP7_75t_L g2444 ( 
.A1(n_2422),
.A2(n_2429),
.B(n_2438),
.C(n_2436),
.Y(n_2444)
);

A2O1A1Ixp33_ASAP7_75t_L g2445 ( 
.A1(n_2439),
.A2(n_269),
.B(n_266),
.C(n_267),
.Y(n_2445)
);

O2A1O1Ixp33_ASAP7_75t_L g2446 ( 
.A1(n_2399),
.A2(n_272),
.B(n_270),
.C(n_271),
.Y(n_2446)
);

AND4x1_ASAP7_75t_L g2447 ( 
.A(n_2409),
.B(n_272),
.C(n_270),
.D(n_271),
.Y(n_2447)
);

NAND3xp33_ASAP7_75t_L g2448 ( 
.A(n_2394),
.B(n_274),
.C(n_275),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2412),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_2449)
);

XNOR2xp5_ASAP7_75t_L g2450 ( 
.A(n_2416),
.B(n_277),
.Y(n_2450)
);

AOI221xp5_ASAP7_75t_L g2451 ( 
.A1(n_2408),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.C(n_281),
.Y(n_2451)
);

A2O1A1Ixp33_ASAP7_75t_L g2452 ( 
.A1(n_2417),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_2452)
);

OAI221xp5_ASAP7_75t_SL g2453 ( 
.A1(n_2419),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.C(n_284),
.Y(n_2453)
);

OAI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2411),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2454)
);

AOI211xp5_ASAP7_75t_L g2455 ( 
.A1(n_2392),
.A2(n_287),
.B(n_285),
.C(n_286),
.Y(n_2455)
);

XOR2x2_ASAP7_75t_L g2456 ( 
.A(n_2403),
.B(n_288),
.Y(n_2456)
);

AOI222xp33_ASAP7_75t_L g2457 ( 
.A1(n_2433),
.A2(n_2420),
.B1(n_2421),
.B2(n_2397),
.C1(n_2415),
.C2(n_2437),
.Y(n_2457)
);

OAI211xp5_ASAP7_75t_SL g2458 ( 
.A1(n_2423),
.A2(n_2435),
.B(n_2425),
.C(n_2400),
.Y(n_2458)
);

AOI211xp5_ASAP7_75t_L g2459 ( 
.A1(n_2418),
.A2(n_292),
.B(n_289),
.C(n_291),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2406),
.Y(n_2460)
);

OAI221xp5_ASAP7_75t_L g2461 ( 
.A1(n_2405),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.C(n_293),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2402),
.B(n_293),
.Y(n_2462)
);

A2O1A1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2404),
.A2(n_297),
.B(n_294),
.C(n_295),
.Y(n_2463)
);

OAI22xp5_ASAP7_75t_L g2464 ( 
.A1(n_2395),
.A2(n_299),
.B1(n_294),
.B2(n_298),
.Y(n_2464)
);

XOR2x2_ASAP7_75t_L g2465 ( 
.A(n_2407),
.B(n_2414),
.Y(n_2465)
);

AOI211x1_ASAP7_75t_L g2466 ( 
.A1(n_2424),
.A2(n_300),
.B(n_298),
.C(n_299),
.Y(n_2466)
);

OAI211xp5_ASAP7_75t_L g2467 ( 
.A1(n_2428),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_2467)
);

OAI221xp5_ASAP7_75t_L g2468 ( 
.A1(n_2426),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.C(n_305),
.Y(n_2468)
);

AOI21xp5_ASAP7_75t_L g2469 ( 
.A1(n_2393),
.A2(n_303),
.B(n_304),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2406),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_2470)
);

OAI31xp33_ASAP7_75t_L g2471 ( 
.A1(n_2392),
.A2(n_310),
.A3(n_306),
.B(n_308),
.Y(n_2471)
);

OAI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2401),
.A2(n_311),
.B(n_312),
.Y(n_2472)
);

OAI21xp33_ASAP7_75t_SL g2473 ( 
.A1(n_2434),
.A2(n_311),
.B(n_312),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_L g2474 ( 
.A1(n_2439),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_2474)
);

AND4x2_ASAP7_75t_L g2475 ( 
.A(n_2396),
.B(n_313),
.C(n_314),
.D(n_316),
.Y(n_2475)
);

OAI211xp5_ASAP7_75t_SL g2476 ( 
.A1(n_2431),
.A2(n_316),
.B(n_317),
.C(n_318),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2439),
.Y(n_2477)
);

O2A1O1Ixp33_ASAP7_75t_L g2478 ( 
.A1(n_2399),
.A2(n_317),
.B(n_318),
.C(n_319),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2406),
.Y(n_2479)
);

OA22x2_ASAP7_75t_L g2480 ( 
.A1(n_2431),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_2480)
);

AOI221x1_ASAP7_75t_L g2481 ( 
.A1(n_2431),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.C(n_323),
.Y(n_2481)
);

OAI211xp5_ASAP7_75t_SL g2482 ( 
.A1(n_2431),
.A2(n_324),
.B(n_325),
.C(n_326),
.Y(n_2482)
);

OAI221xp5_ASAP7_75t_L g2483 ( 
.A1(n_2394),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.C(n_327),
.Y(n_2483)
);

NOR2x1_ASAP7_75t_L g2484 ( 
.A(n_2460),
.B(n_327),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2480),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2477),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2470),
.B(n_331),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2475),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_SL g2489 ( 
.A(n_2477),
.B(n_332),
.Y(n_2489)
);

NOR2x2_ASAP7_75t_L g2490 ( 
.A(n_2479),
.B(n_2450),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2477),
.Y(n_2491)
);

AOI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_2462),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2456),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2446),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2478),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2466),
.Y(n_2496)
);

NAND3xp33_ASAP7_75t_L g2497 ( 
.A(n_2451),
.B(n_335),
.C(n_336),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2471),
.B(n_335),
.Y(n_2498)
);

AOI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2442),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_2465),
.Y(n_2500)
);

AO22x2_ASAP7_75t_L g2501 ( 
.A1(n_2448),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_2501)
);

AOI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2440),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2447),
.Y(n_2503)
);

AOI22xp5_ASAP7_75t_L g2504 ( 
.A1(n_2476),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_2504)
);

AOI22xp33_ASAP7_75t_L g2505 ( 
.A1(n_2482),
.A2(n_2483),
.B1(n_2458),
.B2(n_2441),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2472),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2461),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2468),
.Y(n_2508)
);

HB1xp67_ASAP7_75t_L g2509 ( 
.A(n_2481),
.Y(n_2509)
);

AOI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2454),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_2510)
);

AOI22xp5_ASAP7_75t_L g2511 ( 
.A1(n_2467),
.A2(n_343),
.B1(n_346),
.B2(n_347),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2463),
.Y(n_2512)
);

AOI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2444),
.A2(n_346),
.B1(n_348),
.B2(n_349),
.Y(n_2513)
);

AO22x1_ASAP7_75t_L g2514 ( 
.A1(n_2464),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2443),
.B(n_350),
.Y(n_2515)
);

AOI22xp5_ASAP7_75t_L g2516 ( 
.A1(n_2473),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_2516)
);

NOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2445),
.B(n_351),
.Y(n_2517)
);

AOI22xp5_ASAP7_75t_L g2518 ( 
.A1(n_2449),
.A2(n_352),
.B1(n_353),
.B2(n_355),
.Y(n_2518)
);

INVxp67_ASAP7_75t_SL g2519 ( 
.A(n_2455),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_2453),
.B(n_356),
.Y(n_2520)
);

HB1xp67_ASAP7_75t_L g2521 ( 
.A(n_2459),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2484),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2501),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_L g2524 ( 
.A(n_2491),
.B(n_2452),
.C(n_2469),
.Y(n_2524)
);

NAND4xp75_ASAP7_75t_L g2525 ( 
.A(n_2494),
.B(n_2457),
.C(n_2474),
.D(n_358),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2501),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2515),
.B(n_356),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2514),
.B(n_357),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2509),
.Y(n_2529)
);

AOI21xp5_ASAP7_75t_L g2530 ( 
.A1(n_2498),
.A2(n_357),
.B(n_358),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2490),
.Y(n_2531)
);

NOR2x1_ASAP7_75t_L g2532 ( 
.A(n_2488),
.B(n_359),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2503),
.Y(n_2533)
);

AND3x2_ASAP7_75t_L g2534 ( 
.A(n_2495),
.B(n_360),
.C(n_361),
.Y(n_2534)
);

INVxp67_ASAP7_75t_L g2535 ( 
.A(n_2489),
.Y(n_2535)
);

NOR3xp33_ASAP7_75t_L g2536 ( 
.A(n_2506),
.B(n_2493),
.C(n_2519),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2487),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2496),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2511),
.Y(n_2539)
);

AND2x2_ASAP7_75t_SL g2540 ( 
.A(n_2520),
.B(n_360),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2502),
.B(n_361),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2516),
.Y(n_2542)
);

AND2x4_ASAP7_75t_L g2543 ( 
.A(n_2485),
.B(n_362),
.Y(n_2543)
);

AOI22xp5_ASAP7_75t_L g2544 ( 
.A1(n_2500),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_2544)
);

HB1xp67_ASAP7_75t_L g2545 ( 
.A(n_2517),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_R g2546 ( 
.A(n_2529),
.B(n_2522),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2543),
.B(n_2492),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_R g2548 ( 
.A(n_2540),
.B(n_2512),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_R g2549 ( 
.A(n_2523),
.B(n_2507),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_R g2550 ( 
.A(n_2542),
.B(n_2508),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_L g2551 ( 
.A(n_2536),
.B(n_2505),
.C(n_2521),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2527),
.B(n_2497),
.Y(n_2552)
);

NAND2xp33_ASAP7_75t_SL g2553 ( 
.A(n_2528),
.B(n_2513),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2543),
.B(n_2504),
.Y(n_2554)
);

NAND2xp33_ASAP7_75t_SL g2555 ( 
.A(n_2541),
.B(n_2510),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_R g2556 ( 
.A(n_2539),
.B(n_2518),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2534),
.B(n_2499),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_2531),
.B(n_2486),
.Y(n_2558)
);

NAND2xp33_ASAP7_75t_SL g2559 ( 
.A(n_2545),
.B(n_363),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2532),
.B(n_364),
.Y(n_2560)
);

NAND3xp33_ASAP7_75t_L g2561 ( 
.A(n_2524),
.B(n_365),
.C(n_366),
.Y(n_2561)
);

NAND2xp33_ASAP7_75t_SL g2562 ( 
.A(n_2526),
.B(n_365),
.Y(n_2562)
);

NAND2xp33_ASAP7_75t_SL g2563 ( 
.A(n_2538),
.B(n_366),
.Y(n_2563)
);

XNOR2x1_ASAP7_75t_L g2564 ( 
.A(n_2525),
.B(n_367),
.Y(n_2564)
);

NAND3xp33_ASAP7_75t_SL g2565 ( 
.A(n_2530),
.B(n_367),
.C(n_368),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2553),
.A2(n_2533),
.B1(n_2535),
.B2(n_2537),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2564),
.Y(n_2567)
);

OAI222xp33_ASAP7_75t_L g2568 ( 
.A1(n_2560),
.A2(n_2544),
.B1(n_369),
.B2(n_370),
.C1(n_371),
.C2(n_373),
.Y(n_2568)
);

NAND3xp33_ASAP7_75t_L g2569 ( 
.A(n_2551),
.B(n_368),
.C(n_369),
.Y(n_2569)
);

AO22x2_ASAP7_75t_L g2570 ( 
.A1(n_2558),
.A2(n_370),
.B1(n_373),
.B2(n_417),
.Y(n_2570)
);

NAND5xp2_ASAP7_75t_L g2571 ( 
.A(n_2552),
.B(n_418),
.C(n_422),
.D(n_423),
.E(n_425),
.Y(n_2571)
);

NOR4xp25_ASAP7_75t_L g2572 ( 
.A(n_2565),
.B(n_426),
.C(n_427),
.D(n_430),
.Y(n_2572)
);

NOR2x1_ASAP7_75t_L g2573 ( 
.A(n_2561),
.B(n_431),
.Y(n_2573)
);

AOI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2562),
.A2(n_433),
.B1(n_434),
.B2(n_437),
.Y(n_2574)
);

NOR4xp25_ASAP7_75t_L g2575 ( 
.A(n_2557),
.B(n_2547),
.C(n_2554),
.D(n_2546),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2559),
.B(n_438),
.Y(n_2576)
);

AND4x1_ASAP7_75t_L g2577 ( 
.A(n_2549),
.B(n_439),
.C(n_444),
.D(n_446),
.Y(n_2577)
);

NAND3xp33_ASAP7_75t_SL g2578 ( 
.A(n_2575),
.B(n_2550),
.C(n_2548),
.Y(n_2578)
);

NOR4xp25_ASAP7_75t_L g2579 ( 
.A(n_2567),
.B(n_2556),
.C(n_2555),
.D(n_2563),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_2570),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2572),
.B(n_447),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2569),
.Y(n_2582)
);

CKINVDCx20_ASAP7_75t_R g2583 ( 
.A(n_2566),
.Y(n_2583)
);

NOR2x1p5_ASAP7_75t_L g2584 ( 
.A(n_2576),
.B(n_448),
.Y(n_2584)
);

HB1xp67_ASAP7_75t_L g2585 ( 
.A(n_2570),
.Y(n_2585)
);

AOI221xp5_ASAP7_75t_L g2586 ( 
.A1(n_2568),
.A2(n_449),
.B1(n_452),
.B2(n_453),
.C(n_454),
.Y(n_2586)
);

NAND4xp25_ASAP7_75t_L g2587 ( 
.A(n_2578),
.B(n_2573),
.C(n_2574),
.D(n_2571),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2585),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2584),
.Y(n_2589)
);

OAI22x1_ASAP7_75t_L g2590 ( 
.A1(n_2580),
.A2(n_2577),
.B1(n_456),
.B2(n_457),
.Y(n_2590)
);

INVx2_ASAP7_75t_SL g2591 ( 
.A(n_2581),
.Y(n_2591)
);

CKINVDCx20_ASAP7_75t_R g2592 ( 
.A(n_2583),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2590),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2588),
.B(n_2579),
.Y(n_2594)
);

NAND2x1p5_ASAP7_75t_L g2595 ( 
.A(n_2589),
.B(n_2582),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2592),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2594),
.Y(n_2597)
);

INVx4_ASAP7_75t_L g2598 ( 
.A(n_2595),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2596),
.Y(n_2599)
);

AOI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2598),
.A2(n_2593),
.B1(n_2591),
.B2(n_2587),
.Y(n_2600)
);

AOI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2599),
.A2(n_2586),
.B1(n_459),
.B2(n_460),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_2597),
.A2(n_455),
.B1(n_463),
.B2(n_464),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2600),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2601),
.Y(n_2604)
);

OAI22xp33_ASAP7_75t_L g2605 ( 
.A1(n_2603),
.A2(n_2602),
.B1(n_471),
.B2(n_473),
.Y(n_2605)
);

AOI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2605),
.A2(n_2604),
.B1(n_474),
.B2(n_475),
.Y(n_2606)
);

XNOR2xp5_ASAP7_75t_L g2607 ( 
.A(n_2606),
.B(n_468),
.Y(n_2607)
);

AOI322xp5_ASAP7_75t_L g2608 ( 
.A1(n_2607),
.A2(n_479),
.A3(n_482),
.B1(n_483),
.B2(n_486),
.C1(n_489),
.C2(n_490),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2608),
.A2(n_491),
.B1(n_492),
.B2(n_493),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2609),
.A2(n_494),
.B(n_495),
.Y(n_2610)
);

AOI211xp5_ASAP7_75t_L g2611 ( 
.A1(n_2610),
.A2(n_497),
.B(n_498),
.C(n_499),
.Y(n_2611)
);


endmodule