module fake_jpeg_12814_n_667 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_667);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_667;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_66),
.Y(n_141)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_22),
.B(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_35),
.Y(n_136)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_73),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_29),
.B(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_74),
.B(n_79),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_22),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_75),
.B(n_82),
.Y(n_167)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_10),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_81),
.B(n_43),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_30),
.B(n_34),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_31),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_85),
.A2(n_28),
.B1(n_55),
.B2(n_46),
.Y(n_197)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_86),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_87),
.Y(n_226)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_92),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_95),
.Y(n_184)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_38),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g206 ( 
.A(n_98),
.Y(n_206)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_30),
.B(n_11),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_104),
.B(n_109),
.Y(n_177)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_33),
.B(n_13),
.Y(n_109)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_38),
.B(n_0),
.CON(n_110),
.SN(n_110)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_26),
.B(n_40),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_113),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g205 ( 
.A(n_115),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_24),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g217 ( 
.A(n_116),
.Y(n_217)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_36),
.Y(n_125)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_127),
.B(n_59),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_136),
.B(n_144),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_39),
.B1(n_58),
.B2(n_42),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_139),
.A2(n_159),
.B1(n_165),
.B2(n_0),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_74),
.B(n_40),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_149),
.B(n_168),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_41),
.B1(n_28),
.B2(n_56),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_152),
.A2(n_182),
.B1(n_197),
.B2(n_28),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_59),
.B(n_26),
.C(n_34),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_154),
.A2(n_0),
.B(n_6),
.C(n_7),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_155),
.B(n_194),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_65),
.A2(n_23),
.B1(n_58),
.B2(n_27),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_87),
.A2(n_23),
.B1(n_58),
.B2(n_27),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_79),
.B(n_57),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_64),
.A2(n_21),
.B1(n_20),
.B2(n_56),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_174),
.A2(n_176),
.B1(n_191),
.B2(n_165),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_33),
.B1(n_57),
.B2(n_35),
.Y(n_176)
);

INVx6_ASAP7_75t_SL g178 ( 
.A(n_98),
.Y(n_178)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_178),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_81),
.A2(n_113),
.B1(n_61),
.B2(n_91),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_186),
.A2(n_0),
.B(n_2),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_50),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_187),
.B(n_21),
.Y(n_247)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_188),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_68),
.A2(n_20),
.B1(n_56),
.B2(n_55),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_117),
.A2(n_43),
.B(n_50),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_195),
.B(n_215),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_88),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_123),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_124),
.Y(n_209)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_125),
.B(n_18),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_128),
.Y(n_219)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_73),
.B(n_41),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_37),
.Y(n_246)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_129),
.Y(n_224)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_107),
.Y(n_225)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_169),
.A2(n_94),
.A3(n_83),
.B1(n_37),
.B2(n_55),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_227),
.B(n_243),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_132),
.A2(n_20),
.B1(n_46),
.B2(n_42),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_228),
.A2(n_235),
.B1(n_258),
.B2(n_296),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_139),
.A2(n_21),
.B1(n_46),
.B2(n_42),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_229),
.A2(n_260),
.B1(n_299),
.B2(n_217),
.Y(n_345)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_230),
.Y(n_346)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_231),
.Y(n_356)
);

BUFx8_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

BUFx8_ASAP7_75t_L g321 ( 
.A(n_232),
.Y(n_321)
);

OA22x2_ASAP7_75t_L g352 ( 
.A1(n_234),
.A2(n_280),
.B1(n_133),
.B2(n_223),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_160),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_236),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_137),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_238),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_242),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_134),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_246),
.B(n_275),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_247),
.A2(n_307),
.B(n_218),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_135),
.B(n_59),
.C(n_2),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_248),
.B(n_283),
.C(n_222),
.Y(n_359)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_249),
.Y(n_348)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_138),
.Y(n_250)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_251),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_258),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_257),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_206),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_134),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_259),
.B(n_262),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_177),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_140),
.Y(n_261)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_226),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_263),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_264),
.Y(n_343)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_143),
.Y(n_265)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_180),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_267),
.B(n_274),
.Y(n_340)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_268),
.Y(n_334)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_270),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_212),
.Y(n_272)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_272),
.Y(n_354)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_147),
.Y(n_273)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_213),
.Y(n_275)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_158),
.Y(n_278)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_167),
.B(n_13),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_279),
.B(n_285),
.Y(n_335)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_141),
.Y(n_281)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_281),
.Y(n_360)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_150),
.Y(n_282)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_215),
.B(n_14),
.C(n_4),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_190),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_286),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_151),
.B(n_14),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_141),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_208),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_289),
.Y(n_333)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_153),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g320 ( 
.A1(n_290),
.A2(n_148),
.B(n_196),
.Y(n_320)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_196),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_291),
.B(n_293),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_154),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_292),
.A2(n_296),
.B1(n_297),
.B2(n_301),
.Y(n_317)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_208),
.Y(n_293)
);

BUFx12f_ASAP7_75t_L g294 ( 
.A(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_294),
.B(n_295),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_174),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_161),
.A2(n_6),
.B1(n_8),
.B2(n_14),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_161),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_170),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_298),
.B(n_300),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_191),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_162),
.B(n_152),
.Y(n_300)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_222),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_148),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_302),
.A2(n_303),
.B1(n_305),
.B2(n_133),
.Y(n_351)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_164),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_163),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_304),
.Y(n_350)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_217),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_306),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_192),
.B(n_19),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_309),
.B(n_284),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_211),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_327),
.C(n_363),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_234),
.A2(n_159),
.B1(n_184),
.B2(n_205),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_311),
.A2(n_315),
.B1(n_316),
.B2(n_326),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_280),
.A2(n_184),
.B1(n_205),
.B2(n_200),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_292),
.A2(n_200),
.B1(n_175),
.B2(n_146),
.Y(n_316)
);

AO22x1_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_193),
.B1(n_183),
.B2(n_157),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_318),
.B(n_367),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_320),
.A2(n_368),
.B(n_322),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_324),
.B(n_321),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_227),
.A2(n_256),
.B1(n_283),
.B2(n_241),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_237),
.B(n_145),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_237),
.B(n_202),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_329),
.B(n_297),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_355),
.B1(n_268),
.B2(n_239),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_340),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_244),
.A2(n_183),
.B(n_189),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_353),
.A2(n_232),
.B(n_288),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_260),
.A2(n_193),
.B1(n_146),
.B2(n_157),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_363),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_248),
.B(n_175),
.C(n_181),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_302),
.A2(n_142),
.B1(n_179),
.B2(n_181),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_365),
.A2(n_242),
.B1(n_253),
.B2(n_257),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_238),
.A2(n_179),
.B1(n_164),
.B2(n_223),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_366),
.A2(n_267),
.B1(n_278),
.B2(n_291),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_273),
.B(n_142),
.Y(n_367)
);

OA21x2_ASAP7_75t_L g368 ( 
.A1(n_288),
.A2(n_259),
.B(n_232),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_369),
.B(n_374),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_314),
.A2(n_252),
.B1(n_240),
.B2(n_301),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_370),
.A2(n_380),
.B1(n_392),
.B2(n_417),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_371),
.A2(n_397),
.B(n_412),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_373),
.A2(n_383),
.B1(n_393),
.B2(n_322),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_310),
.B(n_233),
.C(n_269),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_387),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_319),
.A2(n_277),
.B(n_276),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_376),
.A2(n_415),
.B(n_348),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_305),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_378),
.B(n_385),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_379),
.B(n_407),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_345),
.A2(n_263),
.B1(n_298),
.B2(n_236),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_381),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_271),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_403),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_311),
.A2(n_270),
.B1(n_249),
.B2(n_303),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_353),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_367),
.Y(n_386)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_231),
.C(n_230),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_294),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_391),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_389),
.A2(n_390),
.B1(n_410),
.B2(n_416),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_245),
.B1(n_251),
.B2(n_254),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_333),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_315),
.A2(n_272),
.B1(n_294),
.B2(n_365),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_340),
.A2(n_344),
.B1(n_352),
.B2(n_316),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_395),
.Y(n_442)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_413),
.Y(n_429)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_399),
.Y(n_422)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_332),
.Y(n_402)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_358),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_327),
.B(n_335),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_408),
.Y(n_433)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_406),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_313),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_409),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_320),
.A2(n_352),
.B1(n_318),
.B2(n_319),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_411),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_318),
.B(n_319),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_352),
.A2(n_320),
.B1(n_368),
.B2(n_338),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_414),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_368),
.A2(n_328),
.B(n_317),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_337),
.A2(n_364),
.B1(n_338),
.B2(n_334),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_SL g472 ( 
.A(n_419),
.B(n_441),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g421 ( 
.A(n_374),
.B(n_321),
.CI(n_343),
.CON(n_421),
.SN(n_421)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_421),
.B(n_440),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_384),
.A2(n_337),
.B1(n_331),
.B2(n_364),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_423),
.A2(n_380),
.B1(n_396),
.B2(n_399),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_413),
.A2(n_339),
.B(n_348),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_430),
.A2(n_441),
.B(n_446),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_434),
.B(n_398),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_436),
.A2(n_450),
.B(n_394),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_416),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_371),
.A2(n_339),
.B(n_354),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_382),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_451),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_397),
.A2(n_354),
.B(n_321),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_397),
.A2(n_349),
.B1(n_361),
.B2(n_312),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_381),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_411),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_454),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_377),
.A2(n_349),
.B1(n_334),
.B2(n_342),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_453),
.A2(n_455),
.B1(n_389),
.B2(n_390),
.Y(n_481)
);

OAI32xp33_ASAP7_75t_L g454 ( 
.A1(n_377),
.A2(n_308),
.A3(n_357),
.B1(n_346),
.B2(n_341),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_370),
.A2(n_325),
.B1(n_341),
.B2(n_361),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_446),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_467),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_447),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_459),
.B(n_474),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_469),
.C(n_470),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_434),
.B(n_403),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_462),
.B(n_421),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_463),
.A2(n_442),
.B1(n_456),
.B2(n_423),
.Y(n_518)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_465),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_415),
.B(n_412),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_466),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_449),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_478),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_387),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_429),
.B(n_375),
.C(n_404),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

OAI21xp33_ASAP7_75t_L g531 ( 
.A1(n_472),
.A2(n_492),
.B(n_454),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_473),
.A2(n_445),
.B1(n_440),
.B2(n_456),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_453),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_439),
.A2(n_379),
.B(n_394),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_479),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_424),
.B(n_369),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_476),
.B(n_477),
.C(n_480),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_427),
.B(n_400),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_419),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_430),
.A2(n_417),
.B(n_376),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_427),
.B(n_386),
.Y(n_480)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_481),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_424),
.B(n_410),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_482),
.B(n_485),
.C(n_488),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_432),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_483),
.B(n_487),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_436),
.A2(n_417),
.B(n_384),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_433),
.B(n_391),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_438),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_486),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_432),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_433),
.B(n_409),
.C(n_408),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_438),
.A2(n_406),
.B(n_405),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_457),
.Y(n_491)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_491),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g492 ( 
.A(n_455),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_494),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_422),
.Y(n_495)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_496),
.A2(n_481),
.B1(n_452),
.B2(n_451),
.Y(n_559)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_501),
.B(n_480),
.Y(n_538)
);

MAJx2_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_421),
.C(n_425),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_476),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_460),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_511),
.B(n_515),
.Y(n_545)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_460),
.Y(n_513)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_513),
.Y(n_551)
);

BUFx4f_ASAP7_75t_SL g514 ( 
.A(n_483),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_514),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_487),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_418),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_516),
.B(n_522),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_518),
.A2(n_464),
.B(n_484),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_490),
.A2(n_442),
.B1(n_448),
.B2(n_418),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_490),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_488),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_463),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_461),
.B(n_425),
.Y(n_522)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_471),
.Y(n_525)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_525),
.Y(n_558)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_494),
.Y(n_527)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_527),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_462),
.B(n_444),
.C(n_450),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_528),
.B(n_482),
.C(n_485),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_467),
.A2(n_445),
.B1(n_443),
.B2(n_448),
.Y(n_529)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_529),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_531),
.B(n_475),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_509),
.B(n_468),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_532),
.B(n_540),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_533),
.B(n_535),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_534),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_493),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_536),
.B(n_538),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_512),
.B(n_477),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_537),
.B(n_539),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_526),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_524),
.B(n_489),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_541),
.B(n_513),
.Y(n_564)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_542),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_506),
.B(n_478),
.C(n_466),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_544),
.C(n_547),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_506),
.B(n_458),
.C(n_479),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_526),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_546),
.B(n_507),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_524),
.B(n_464),
.C(n_495),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_516),
.B(n_431),
.C(n_491),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_553),
.C(n_510),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_523),
.Y(n_549)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_549),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_503),
.B(n_510),
.Y(n_550)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_550),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_521),
.B(n_431),
.C(n_443),
.Y(n_553)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_554),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_522),
.B(n_443),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_555),
.B(n_557),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_501),
.B(n_473),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_559),
.A2(n_518),
.B1(n_525),
.B2(n_527),
.Y(n_584)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_561),
.A2(n_499),
.B1(n_503),
.B2(n_507),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_566),
.A2(n_581),
.B1(n_559),
.B2(n_541),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_570),
.B(n_569),
.Y(n_606)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_573),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_553),
.B(n_508),
.C(n_528),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_580),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_535),
.B(n_517),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_576),
.B(n_533),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_545),
.B(n_514),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_579),
.B(n_582),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_530),
.C(n_500),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_551),
.A2(n_499),
.B1(n_519),
.B2(n_504),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_550),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_584),
.A2(n_542),
.B1(n_560),
.B2(n_558),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_544),
.B(n_504),
.C(n_505),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_585),
.B(n_587),
.C(n_555),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_586),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_543),
.B(n_505),
.C(n_498),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_565),
.B(n_536),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_588),
.B(n_604),
.Y(n_622)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_SL g619 ( 
.A(n_591),
.B(n_568),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_577),
.B(n_562),
.Y(n_592)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_592),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_593),
.B(n_594),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_570),
.B(n_556),
.C(n_557),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_562),
.Y(n_595)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_595),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_556),
.C(n_538),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_596),
.B(n_601),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_571),
.A2(n_534),
.B(n_542),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_598),
.A2(n_592),
.B(n_599),
.Y(n_618)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_599),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_567),
.B(n_585),
.C(n_587),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_583),
.B(n_514),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_576),
.B(n_498),
.C(n_552),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_605),
.B(n_607),
.C(n_563),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_606),
.B(n_568),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_575),
.B(n_552),
.C(n_502),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_584),
.A2(n_437),
.B1(n_435),
.B2(n_426),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_608),
.A2(n_581),
.B1(n_578),
.B2(n_566),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_609),
.B(n_623),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_610),
.A2(n_428),
.B1(n_426),
.B2(n_435),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_601),
.B(n_603),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_611),
.B(n_612),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_598),
.A2(n_574),
.B(n_564),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_597),
.A2(n_574),
.B1(n_580),
.B2(n_569),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_614),
.B(n_624),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_618),
.B(n_595),
.Y(n_631)
);

XNOR2x1_ASAP7_75t_L g632 ( 
.A(n_619),
.B(n_625),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_600),
.B(n_497),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_SL g625 ( 
.A(n_591),
.B(n_563),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_593),
.B(n_437),
.C(n_428),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_626),
.B(n_401),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_620),
.B(n_602),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_628),
.B(n_630),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_621),
.A2(n_589),
.B(n_607),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_629),
.A2(n_638),
.B(n_634),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_623),
.B(n_606),
.C(n_594),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_631),
.B(n_640),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_622),
.B(n_605),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_633),
.B(n_634),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_609),
.B(n_596),
.C(n_608),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_635),
.B(n_637),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_614),
.B(n_457),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_636),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g637 ( 
.A(n_615),
.B(n_372),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_641),
.A2(n_644),
.B(n_643),
.Y(n_651)
);

AOI21xp33_ASAP7_75t_L g642 ( 
.A1(n_627),
.A2(n_612),
.B(n_616),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g657 ( 
.A1(n_642),
.A2(n_647),
.B(n_646),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_630),
.A2(n_618),
.B(n_626),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_631),
.B(n_613),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_648),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_639),
.B(n_624),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_649),
.B(n_617),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_651),
.B(n_657),
.C(n_625),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_650),
.B(n_636),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_652),
.B(n_654),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_645),
.A2(n_617),
.B(n_632),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_655),
.B(n_656),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_645),
.A2(n_632),
.B(n_619),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_658),
.B(n_659),
.C(n_660),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_653),
.B(n_654),
.Y(n_661)
);

AO21x1_ASAP7_75t_L g662 ( 
.A1(n_661),
.A2(n_346),
.B(n_357),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_662),
.B(n_663),
.C(n_372),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_664),
.B(n_402),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_665),
.B(n_401),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_666),
.A2(n_402),
.B(n_325),
.Y(n_667)
);


endmodule