module fake_jpeg_29970_n_94 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_11),
.C(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_45),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_48),
.Y(n_62)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_42),
.B1(n_47),
.B2(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_37),
.B1(n_31),
.B2(n_29),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_28),
.C(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_56),
.B(n_52),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_66),
.B1(n_59),
.B2(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_66),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_51),
.B1(n_4),
.B2(n_6),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_73),
.C(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_12),
.C(n_21),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_78),
.B1(n_80),
.B2(n_75),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_82),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_88),
.A2(n_86),
.B1(n_4),
.B2(n_6),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_13),
.A3(n_19),
.B1(n_8),
.B2(n_9),
.C1(n_25),
.C2(n_15),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_91),
.C(n_16),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_2),
.Y(n_94)
);


endmodule