module real_jpeg_19873_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx13_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_59),
.B1(n_69),
.B2(n_84),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_84),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_84),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_3),
.A2(n_64),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_3),
.B(n_72),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_37),
.B(n_41),
.C(n_130),
.D(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_3),
.B(n_37),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_82),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_3),
.A2(n_24),
.B(n_145),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g175 ( 
.A1(n_3),
.A2(n_65),
.B(n_77),
.C(n_96),
.D(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_3),
.B(n_65),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_4),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_87),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_87),
.Y(n_174)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_6),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_6),
.A2(n_25),
.B1(n_105),
.B2(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_6),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_47),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_10),
.A2(n_55),
.B1(n_59),
.B2(n_69),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_10),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_55),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_107),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_88),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_24),
.A2(n_28),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_24),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_25),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_25),
.B(n_146),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_27),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_26),
.B(n_42),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_26),
.B(n_164),
.Y(n_163)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_27),
.A2(n_43),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_32),
.A2(n_151),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_32),
.A2(n_160),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_48),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_37),
.A2(n_38),
.B1(n_78),
.B2(n_79),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_37),
.B(n_78),
.Y(n_182)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_38),
.A2(n_81),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_40),
.A2(n_48),
.B1(n_142),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_40),
.A2(n_174),
.B(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_53),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_48),
.B(n_54),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_48),
.A2(n_52),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_48),
.B(n_68),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.C(n_74),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_51),
.B1(n_74),
.B2(n_75),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B(n_70),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_61),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_61),
.B(n_68),
.C(n_102),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_78),
.B(n_81),
.C(n_82),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_68),
.B(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_86),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_85),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B1(n_94),
.B2(n_98),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_112),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_108),
.B(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_119),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_115),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_119),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_120),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_200),
.B(n_205),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_187),
.B(n_199),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_168),
.B(n_186),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_147),
.B(n_167),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_136),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_131),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_144),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_156),
.B(n_166),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_154),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_161),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_159),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_170),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_179),
.B2(n_185),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_178),
.C(n_185),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_183),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_189),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_195),
.C(n_197),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_191),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);


endmodule