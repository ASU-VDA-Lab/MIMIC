module fake_jpeg_1942_n_174 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_67),
.Y(n_75)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_0),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_54),
.CON(n_70),
.SN(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_78),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_67),
.B1(n_52),
.B2(n_61),
.Y(n_87)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_92),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_62),
.B(n_45),
.C(n_47),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_88),
.B(n_90),
.C(n_74),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_89),
.B1(n_93),
.B2(n_36),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_56),
.B(n_59),
.C(n_55),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_53),
.B1(n_57),
.B2(n_65),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_76),
.B(n_60),
.C(n_53),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_58),
.B1(n_48),
.B2(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_62),
.B1(n_61),
.B2(n_52),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_77),
.B1(n_74),
.B2(n_21),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_1),
.B(n_2),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_3),
.B(n_4),
.Y(n_116)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_80),
.B1(n_74),
.B2(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_115),
.B1(n_113),
.B2(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_106),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_85),
.B1(n_81),
.B2(n_96),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_22),
.Y(n_118)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_113),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_116),
.B(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_2),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_104),
.A2(n_88),
.B(n_9),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_134),
.B(n_14),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_118),
.A2(n_133),
.B1(n_116),
.B2(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_8),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_8),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_23),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_130),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_10),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_24),
.B1(n_34),
.B2(n_32),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_136),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_29),
.C(n_28),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_138),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_25),
.C(n_12),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_142),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

XOR2x1_ASAP7_75t_SL g143 ( 
.A(n_128),
.B(n_11),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_145),
.B(n_133),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_14),
.C(n_15),
.Y(n_147)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_135),
.B(n_117),
.C(n_119),
.D(n_134),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_19),
.B1(n_128),
.B2(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_156),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_145),
.B1(n_150),
.B2(n_143),
.Y(n_163)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_137),
.C(n_136),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_160),
.C(n_152),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_144),
.C(n_146),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_155),
.C(n_127),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_165),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_161),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_166),
.CI(n_156),
.CON(n_170),
.SN(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_171),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_138),
.B(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.Y(n_174)
);


endmodule