module real_jpeg_18700_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_423),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_0),
.B(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_1),
.A2(n_299),
.B1(n_303),
.B2(n_304),
.Y(n_298)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_1),
.A2(n_305),
.B1(n_410),
.B2(n_414),
.Y(n_409)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_4),
.A2(n_54),
.B1(n_123),
.B2(n_126),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_4),
.A2(n_54),
.B1(n_144),
.B2(n_147),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_54),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_30),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_5),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_5),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_5),
.A2(n_30),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_5),
.B(n_128),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_5),
.B(n_231),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_6),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_7),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_7),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_7),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_8),
.A2(n_308),
.B1(n_313),
.B2(n_314),
.Y(n_307)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_8),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_8),
.A2(n_199),
.B1(n_313),
.B2(n_351),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_9),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_12),
.Y(n_156)
);

BUFx4f_ASAP7_75t_L g312 ( 
.A(n_12),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

XOR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_398),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

AO221x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_292),
.B1(n_391),
.B2(n_396),
.C(n_397),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_222),
.B(n_291),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_185),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_20),
.B(n_185),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_129),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_21),
.B(n_130),
.C(n_163),
.Y(n_387)
);

XOR2x1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_58),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_23),
.B(n_336),
.C(n_341),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_23),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_24),
.A2(n_25),
.B1(n_342),
.B2(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_24),
.B(n_60),
.C(n_85),
.Y(n_385)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_34),
.B1(n_44),
.B2(n_52),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g317 ( 
.A1(n_26),
.A2(n_34),
.B1(n_44),
.B2(n_52),
.Y(n_317)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_26),
.Y(n_358)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_42),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_30),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_30),
.B(n_57),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_30),
.B(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_34),
.B(n_44),
.Y(n_359)
);

OAI21x1_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_41),
.B(n_44),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_35),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_44),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_45),
.Y(n_175)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_45),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_85),
.B2(n_86),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_70),
.B(n_79),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_61),
.A2(n_70),
.B1(n_79),
.B2(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_61),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_61),
.B(n_70),
.Y(n_407)
);

NAND2x1p5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_70),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_65),
.Y(n_215)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_69),
.Y(n_256)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_70),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_70),
.A2(n_321),
.B(n_331),
.Y(n_320)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_73),
.Y(n_268)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_77),
.Y(n_250)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_79),
.Y(n_229)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_85),
.A2(n_86),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_85),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_85),
.A2(n_86),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22x1_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_110),
.B1(n_122),
.B2(n_128),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_87),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_87),
.A2(n_110),
.B(n_128),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_87),
.A2(n_110),
.B1(n_128),
.B2(n_409),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_103),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_94),
.B1(n_98),
.B2(n_102),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_99),
.Y(n_208)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

OA22x2_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_105),
.Y(n_244)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_105),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_116),
.A2(n_203),
.A3(n_205),
.B1(n_206),
.B2(n_209),
.Y(n_202)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_121),
.Y(n_417)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_163),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.C(n_137),
.Y(n_130)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_131),
.B(n_349),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_131),
.A2(n_193),
.B1(n_317),
.B2(n_318),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_137),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_137),
.B(n_259),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_142),
.B(n_150),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_151),
.B1(n_157),
.B2(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_146),
.Y(n_314)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_150),
.A2(n_298),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_151),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_151),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_153),
.Y(n_340)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_159),
.Y(n_252)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_179),
.B2(n_180),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_165),
.B(n_179),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_176),
.B2(n_178),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_179),
.A2(n_180),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_180),
.B(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_180),
.B(n_270),
.Y(n_271)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_194),
.C(n_201),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_186),
.A2(n_187),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_191),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_191),
.B(n_240),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_192),
.B(n_317),
.C(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21x1_ASAP7_75t_L g347 ( 
.A1(n_193),
.A2(n_348),
.B(n_353),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_235),
.C(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_194),
.A2(n_236),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_194),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_194),
.A2(n_201),
.B1(n_278),
.B2(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_194),
.A2(n_278),
.B1(n_297),
.B2(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_201),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_216),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_SL g333 ( 
.A(n_218),
.B(n_307),
.Y(n_333)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_282),
.B(n_290),
.Y(n_222)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_237),
.B(n_281),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_234),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_233),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_227),
.A2(n_228),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_227),
.A2(n_228),
.B1(n_338),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_R g274 ( 
.A(n_228),
.B(n_242),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_228),
.B(n_338),
.Y(n_337)
);

AO22x2_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_229),
.B(n_230),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_230),
.A2(n_231),
.B1(n_322),
.B2(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_284),
.C(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_236),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_273),
.B(n_280),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_257),
.B(n_272),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_245),
.A3(n_249),
.B1(n_251),
.B2(n_253),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_269),
.B(n_271),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_267),
.Y(n_303)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_275),
.Y(n_280)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_361),
.C(n_374),
.Y(n_292)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_293),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_343),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_294),
.B(n_343),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_319),
.C(n_335),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_295),
.B(n_319),
.Y(n_373)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_316),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_317),
.C(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_306),
.B1(n_307),
.B2(n_315),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_323),
.B1(n_327),
.B2(n_330),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_320),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_333),
.Y(n_355)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_333),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g419 ( 
.A1(n_333),
.A2(n_355),
.B(n_357),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_373),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_338),
.Y(n_383)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_344),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_354),
.C(n_401),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_407),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_404),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_392),
.B(n_393),
.C(n_395),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_372),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_372),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_368),
.C(n_370),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_364),
.A2(n_365),
.B1(n_368),
.B2(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_368),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_377),
.Y(n_376)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_386),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_379),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_382),
.C(n_384),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_382),
.A2(n_384),
.B1(n_385),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_382),
.Y(n_390)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NOR2x1_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_388),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_421),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_400),
.B(n_402),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_402)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);


endmodule