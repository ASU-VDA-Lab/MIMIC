module fake_jpeg_17037_n_139 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_10),
.B(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_13),
.B(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NAND3xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_22),
.C(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_14),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_20),
.B1(n_19),
.B2(n_13),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_20),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_26),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_31),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_42),
.Y(n_66)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_27),
.C(n_36),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_37),
.C(n_22),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_11),
.B1(n_31),
.B2(n_22),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_56),
.Y(n_59)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_68),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_54),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_84),
.B1(n_88),
.B2(n_91),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_42),
.C(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_47),
.B1(n_34),
.B2(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_87),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_47),
.B(n_52),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_53),
.B(n_18),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_34),
.B1(n_24),
.B2(n_58),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_23),
.B(n_28),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_72),
.C(n_65),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_2),
.B(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_81),
.B(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_73),
.C(n_68),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_101),
.C(n_86),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_79),
.C(n_81),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_104),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_106),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_89),
.B(n_84),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_103),
.B(n_95),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_112),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_66),
.C(n_60),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_66),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_18),
.B(n_70),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_100),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_67),
.C(n_29),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_93),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_102),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

AOI31xp67_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_102),
.A3(n_67),
.B(n_23),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_114),
.B1(n_120),
.B2(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_29),
.C(n_71),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_4),
.C(n_9),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_119),
.B1(n_2),
.B2(n_5),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_4),
.B(n_7),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_131),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_9),
.C(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_136),
.Y(n_139)
);


endmodule