module fake_jpeg_14688_n_328 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_328);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_44),
.B1(n_31),
.B2(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_60),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_26),
.Y(n_53)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_1),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_42),
.B1(n_32),
.B2(n_24),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_32),
.Y(n_98)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_23),
.B(n_3),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_23),
.Y(n_99)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_34),
.B1(n_24),
.B2(n_42),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_67),
.C(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_97),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_40),
.B1(n_30),
.B2(n_55),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_83),
.A2(n_103),
.B1(n_104),
.B2(n_73),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_40),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_68),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_101),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_49),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_44),
.B1(n_20),
.B2(n_31),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_34),
.B1(n_70),
.B2(n_72),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_141)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_113),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_65),
.B1(n_47),
.B2(n_63),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_137),
.B1(n_138),
.B2(n_96),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_121),
.B1(n_125),
.B2(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_27),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx4f_ASAP7_75t_SL g155 ( 
.A(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_58),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_133),
.Y(n_156)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_132),
.B(n_136),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_99),
.Y(n_129)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_27),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_66),
.Y(n_133)
);

AO22x2_ASAP7_75t_L g135 ( 
.A1(n_74),
.A2(n_66),
.B1(n_48),
.B2(n_62),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_135),
.A2(n_129),
.B1(n_133),
.B2(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_83),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_131),
.B1(n_125),
.B2(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_56),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_109),
.B1(n_135),
.B2(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_128),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_84),
.B1(n_91),
.B2(n_69),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_52),
.B1(n_87),
.B2(n_76),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_104),
.B(n_64),
.C(n_67),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_59),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_134),
.B1(n_121),
.B2(n_126),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_163),
.A2(n_165),
.B(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_116),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_164),
.B(n_167),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_110),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_75),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_170),
.C(n_173),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_147),
.B(n_156),
.Y(n_169)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_141),
.A3(n_145),
.B1(n_142),
.B2(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_118),
.C(n_137),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_153),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_156),
.A2(n_117),
.B(n_108),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_156),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_75),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_177),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_146),
.A2(n_107),
.B1(n_127),
.B2(n_114),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_179),
.B(n_154),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_189),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_183),
.A2(n_155),
.B(n_35),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_192),
.B1(n_196),
.B2(n_79),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_160),
.B1(n_149),
.B2(n_157),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_191),
.B1(n_195),
.B2(n_180),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_157),
.B1(n_143),
.B2(n_123),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_174),
.B1(n_173),
.B2(n_165),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_143),
.B1(n_140),
.B2(n_87),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_168),
.B1(n_178),
.B2(n_167),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_172),
.B(n_162),
.C(n_164),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_200),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_201),
.C(n_209),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_178),
.B1(n_177),
.B2(n_155),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_207),
.B1(n_210),
.B2(n_180),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_194),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_206),
.B(n_212),
.Y(n_224)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_154),
.B(n_33),
.C(n_81),
.D(n_27),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_155),
.B1(n_78),
.B2(n_76),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_155),
.C(n_59),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_43),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_186),
.B(n_190),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_208),
.B1(n_211),
.B2(n_79),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_220),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_196),
.B1(n_182),
.B2(n_184),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_222),
.A2(n_227),
.B1(n_206),
.B2(n_197),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_191),
.C(n_195),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_199),
.C(n_202),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_187),
.Y(n_226)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_187),
.B1(n_185),
.B2(n_78),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_27),
.CI(n_39),
.CON(n_228),
.SN(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_213),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_207),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_238),
.C(n_244),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_226),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_236),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_221),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_219),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_248),
.B1(n_221),
.B2(n_222),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_154),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_244),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_223),
.B(n_3),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_254),
.C(n_247),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_263),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_214),
.B1(n_215),
.B2(n_225),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_260),
.B1(n_5),
.B2(n_8),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_230),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_256),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_214),
.B(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_224),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_9),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_228),
.B1(n_217),
.B2(n_81),
.Y(n_260)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_228),
.B1(n_43),
.B2(n_41),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_239),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_240),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_240),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_41),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_265),
.C(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_264),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_278),
.B(n_281),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_262),
.B1(n_249),
.B2(n_15),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_275),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_9),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_256),
.C(n_253),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_293),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_262),
.C(n_61),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_272),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_303),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_289),
.A2(n_280),
.B1(n_271),
.B2(n_15),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_12),
.B(n_13),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_285),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_307),
.C(n_313),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_288),
.B(n_284),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_285),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_309),
.B(n_312),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_292),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_303),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_295),
.C(n_283),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_319),
.B(n_310),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_300),
.B(n_16),
.Y(n_316)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_316),
.A2(n_320),
.B(n_35),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_12),
.Y(n_319)
);

AOI21x1_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_17),
.B(n_18),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_323),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_314),
.B(n_17),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_37),
.B(n_39),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_37),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_325),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_317),
.B(n_61),
.Y(n_328)
);


endmodule