module fake_jpeg_30683_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_48),
.Y(n_141)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_28),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_81),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_56),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_28),
.A2(n_8),
.B1(n_13),
.B2(n_3),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_58),
.A2(n_35),
.B1(n_82),
.B2(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_32),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_73),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_17),
.B(n_14),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_82),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_80),
.Y(n_111)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_87),
.Y(n_121)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_32),
.B(n_6),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_6),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_31),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_30),
.B1(n_23),
.B2(n_22),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_106),
.B1(n_114),
.B2(n_118),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_11),
.B(n_13),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_103),
.B(n_107),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_23),
.B1(n_43),
.B2(n_36),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_19),
.B(n_41),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_47),
.A2(n_42),
.B1(n_36),
.B2(n_19),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_139),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_125),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_39),
.B1(n_37),
.B2(n_31),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_126),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_37),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_38),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_35),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_135),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_54),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_140),
.B1(n_69),
.B2(n_55),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_51),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_4),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_48),
.B(n_51),
.CON(n_139),
.SN(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_63),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_147),
.A2(n_155),
.B1(n_156),
.B2(n_161),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_153),
.Y(n_204)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_68),
.B1(n_53),
.B2(n_77),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_91),
.A2(n_59),
.B1(n_72),
.B2(n_71),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_75),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_168),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_160),
.B(n_172),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_81),
.B1(n_57),
.B2(n_46),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_69),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_167),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_175),
.Y(n_201)
);

AOI22x1_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_52),
.B1(n_60),
.B2(n_65),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_176),
.B1(n_182),
.B2(n_174),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_118),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_178),
.B1(n_181),
.B2(n_187),
.Y(n_197)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_10),
.C(n_11),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_10),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_106),
.A2(n_11),
.B1(n_114),
.B2(n_138),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_130),
.B1(n_131),
.B2(n_149),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_92),
.B(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_97),
.B(n_111),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_96),
.A2(n_99),
.B1(n_102),
.B2(n_136),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_102),
.A2(n_96),
.B1(n_95),
.B2(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_111),
.B(n_110),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_186),
.Y(n_215)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_95),
.A2(n_128),
.B1(n_141),
.B2(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_188),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_184),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_93),
.B(n_143),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_94),
.B(n_123),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_94),
.A2(n_123),
.B1(n_112),
.B2(n_115),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_120),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_160),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_101),
.B(n_140),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_194),
.A2(n_214),
.B1(n_206),
.B2(n_197),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_163),
.B1(n_152),
.B2(n_151),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_203),
.B1(n_210),
.B2(n_212),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_207),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_149),
.B1(n_175),
.B2(n_176),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_214),
.B1(n_197),
.B2(n_222),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_172),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_146),
.A2(n_179),
.B1(n_149),
.B2(n_162),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_162),
.A2(n_164),
.B1(n_157),
.B2(n_176),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_164),
.A2(n_180),
.B1(n_188),
.B2(n_150),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_217),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_158),
.A2(n_145),
.B1(n_167),
.B2(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_173),
.B1(n_198),
.B2(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_166),
.B(n_148),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_173),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_226),
.A2(n_247),
.B1(n_206),
.B2(n_204),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_201),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_238),
.Y(n_265)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_231),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g231 ( 
.A(n_195),
.B(n_215),
.C(n_211),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_210),
.B(n_219),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_239),
.A2(n_227),
.B1(n_249),
.B2(n_248),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_218),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_212),
.B(n_192),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_191),
.C(n_223),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_193),
.C(n_208),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_190),
.B(n_214),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_206),
.B(n_204),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_208),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_269),
.B1(n_242),
.B2(n_225),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_266),
.C(n_246),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_257),
.A2(n_269),
.B(n_250),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_200),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_200),
.C(n_238),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_235),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_232),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

AO22x1_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_248),
.B1(n_239),
.B2(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_275),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_263),
.B1(n_252),
.B2(n_241),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_228),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_233),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_283),
.C(n_285),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_233),
.C(n_231),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_281),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_237),
.B(n_240),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_224),
.C(n_237),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_260),
.B1(n_264),
.B2(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_224),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_275),
.B(n_273),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_264),
.B1(n_256),
.B2(n_265),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_294),
.B1(n_295),
.B2(n_297),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_270),
.B1(n_279),
.B2(n_285),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_287),
.B1(n_290),
.B2(n_294),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_251),
.B1(n_252),
.B2(n_236),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_255),
.C(n_229),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_283),
.C(n_276),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_277),
.A2(n_254),
.B1(n_268),
.B2(n_255),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_300),
.C(n_305),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_280),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_301),
.A2(n_302),
.B1(n_299),
.B2(n_307),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_272),
.B1(n_254),
.B2(n_245),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_272),
.B(n_245),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_292),
.B(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_288),
.B1(n_297),
.B2(n_293),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_289),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_311),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_292),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_313),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_315),
.B(n_302),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_321),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

OAI221xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_298),
.B1(n_305),
.B2(n_308),
.C(n_311),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_312),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_315),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_325),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_314),
.B(n_320),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_309),
.B(n_312),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_327),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_309),
.Y(n_333)
);


endmodule