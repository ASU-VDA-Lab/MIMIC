module fake_jpeg_6701_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_44),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_23),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_64),
.B1(n_66),
.B2(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_55),
.Y(n_86)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_29),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_24),
.B1(n_31),
.B2(n_23),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_70),
.Y(n_71)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_24),
.B1(n_31),
.B2(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_31),
.B1(n_24),
.B2(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_37),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_92),
.C(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_26),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_26),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_55),
.B1(n_47),
.B2(n_63),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_102),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_34),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_39),
.B1(n_58),
.B2(n_46),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_107),
.B1(n_30),
.B2(n_91),
.Y(n_148)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_58),
.B1(n_46),
.B2(n_36),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_112),
.Y(n_127)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_110),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_37),
.B1(n_65),
.B2(n_36),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_108),
.Y(n_139)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_76),
.A2(n_37),
.B1(n_42),
.B2(n_38),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_76),
.A2(n_38),
.B1(n_42),
.B2(n_59),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_73),
.B(n_75),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_76),
.A2(n_42),
.B1(n_38),
.B2(n_32),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_85),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_141),
.C(n_118),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_135),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_93),
.B1(n_79),
.B2(n_72),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_130),
.B1(n_30),
.B2(n_121),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_93),
.B1(n_79),
.B2(n_74),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_92),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_93),
.B1(n_86),
.B2(n_95),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_145),
.B1(n_148),
.B2(n_77),
.Y(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_29),
.B(n_27),
.Y(n_162)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_88),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_97),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_95),
.B1(n_83),
.B2(n_82),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_83),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_169),
.C(n_142),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_117),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_160),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_174),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_110),
.B1(n_102),
.B2(n_115),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_144),
.B1(n_143),
.B2(n_129),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_123),
.A2(n_116),
.B1(n_115),
.B2(n_78),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_161),
.B1(n_168),
.B2(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_34),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_162),
.B(n_165),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_78),
.B1(n_97),
.B2(n_91),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_18),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_128),
.A2(n_78),
.B1(n_16),
.B2(n_17),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_18),
.Y(n_167)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_56),
.C(n_38),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_171),
.B(n_172),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_56),
.B(n_22),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_0),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_173),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_18),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_133),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_178),
.B(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_130),
.B1(n_129),
.B2(n_131),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_196),
.B1(n_150),
.B2(n_166),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_188),
.B1(n_33),
.B2(n_17),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_148),
.B1(n_134),
.B2(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_103),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_149),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_192),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_127),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_127),
.B1(n_134),
.B2(n_142),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_21),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_169),
.C(n_160),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_22),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_217),
.C(n_215),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_194),
.B(n_189),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_208),
.A2(n_210),
.B1(n_212),
.B2(n_221),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_153),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_150),
.B1(n_162),
.B2(n_159),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_153),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_157),
.B1(n_172),
.B2(n_144),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_198),
.B1(n_180),
.B2(n_187),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_18),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_42),
.C(n_52),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_18),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_21),
.B1(n_42),
.B2(n_17),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_22),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_189),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_21),
.B1(n_33),
.B2(n_45),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_183),
.B1(n_33),
.B2(n_21),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_230),
.C(n_215),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_200),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_183),
.C(n_177),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_0),
.B(n_1),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_22),
.B1(n_52),
.B2(n_45),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_244),
.B(n_223),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_243),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_178),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_22),
.B(n_1),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_204),
.B1(n_218),
.B2(n_203),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_69),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_226),
.C(n_230),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_211),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_227),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_202),
.B1(n_212),
.B2(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_255),
.B1(n_241),
.B2(n_242),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_245),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_257),
.B(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_221),
.B1(n_222),
.B2(n_69),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_225),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_259),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_22),
.B(n_1),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_245),
.B1(n_228),
.B2(n_234),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_250),
.B(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_266),
.C(n_271),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_231),
.B(n_237),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_278),
.B1(n_258),
.B2(n_2),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_247),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_249),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_275),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_259),
.B(n_255),
.C(n_256),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_233),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_260),
.C(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_254),
.A2(n_52),
.B1(n_45),
.B2(n_3),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_288),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_281),
.A2(n_268),
.B1(n_278),
.B2(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_274),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_260),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_6),
.C(n_14),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_273),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_15),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_9),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_10),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_289),
.B(n_13),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_292),
.B(n_294),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_271),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_296),
.C(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_297),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_0),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_285),
.B(n_6),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_281),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_6),
.Y(n_306)
);

AOI31xp33_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_287),
.A3(n_280),
.B(n_284),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_12),
.B(n_13),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_SL g302 ( 
.A1(n_291),
.A2(n_290),
.B(n_280),
.C(n_11),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND4xp25_ASAP7_75t_SL g303 ( 
.A(n_296),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_15),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_12),
.C(n_13),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_309),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_301),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_307),
.C(n_313),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_4),
.A3(n_5),
.B1(n_304),
.B2(n_315),
.C1(n_301),
.C2(n_299),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.Y(n_319)
);


endmodule