module fake_netlist_5_471_n_2840 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2840);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2840;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_680;
wire n_1587;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1534;
wire n_1354;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_1312;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_2097;
wire n_1834;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_2722;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_698;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_733;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_597;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_52),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_135),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_553),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_510),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_8),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_193),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_466),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_69),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_259),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_574),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_308),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_468),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_543),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_555),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_79),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_447),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_163),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_259),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_407),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_552),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_250),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_193),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_325),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_222),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_363),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_191),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_576),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_106),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_252),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_324),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_539),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_268),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_257),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_164),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_208),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_422),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_118),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_423),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_220),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_9),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_406),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_384),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_386),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_462),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_403),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_268),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_401),
.Y(n_633)
);

CKINVDCx14_ASAP7_75t_R g634 ( 
.A(n_505),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_1),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_171),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_498),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_203),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_22),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_316),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_26),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_500),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_63),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_192),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_27),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_285),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_345),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_385),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_421),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_547),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_177),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_331),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_104),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_467),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_521),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_294),
.Y(n_656)
);

CKINVDCx14_ASAP7_75t_R g657 ( 
.A(n_171),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_118),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_550),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_173),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_565),
.Y(n_661)
);

CKINVDCx14_ASAP7_75t_R g662 ( 
.A(n_506),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_360),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_560),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_247),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_377),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_572),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_114),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_174),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_531),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_463),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_382),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_31),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_76),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_290),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_447),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_402),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_571),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_488),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_437),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_302),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_419),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_140),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_469),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_340),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_453),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_308),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_212),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_162),
.Y(n_689)
);

CKINVDCx11_ASAP7_75t_R g690 ( 
.A(n_64),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_361),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_333),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_134),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_43),
.Y(n_695)
);

CKINVDCx16_ASAP7_75t_R g696 ( 
.A(n_396),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_566),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_485),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_146),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_209),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_181),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_481),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_579),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_57),
.Y(n_704)
);

BUFx5_ASAP7_75t_L g705 ( 
.A(n_463),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_373),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_419),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_385),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_491),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_48),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_219),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_460),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_424),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_548),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_542),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_242),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_452),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_33),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_205),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_176),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_204),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_143),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_561),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_114),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_465),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_50),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_399),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_437),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_395),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_151),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_103),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_88),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_315),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_289),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_144),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_457),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_241),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_556),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_557),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_191),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_562),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_559),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_253),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_68),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_567),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_494),
.Y(n_746)
);

CKINVDCx14_ASAP7_75t_R g747 ( 
.A(n_195),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_493),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_135),
.Y(n_749)
);

BUFx5_ASAP7_75t_L g750 ( 
.A(n_584),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_178),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_522),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_255),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_406),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_427),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_546),
.Y(n_756)
);

CKINVDCx14_ASAP7_75t_R g757 ( 
.A(n_337),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_332),
.Y(n_758)
);

CKINVDCx14_ASAP7_75t_R g759 ( 
.A(n_527),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_184),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_214),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_538),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_346),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_134),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_517),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_507),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_465),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_104),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_312),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_545),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_194),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_476),
.Y(n_772)
);

BUFx10_ASAP7_75t_L g773 ( 
.A(n_316),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_404),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_241),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_328),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_196),
.Y(n_777)
);

BUFx10_ASAP7_75t_L g778 ( 
.A(n_66),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_583),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_218),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_317),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_549),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_21),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_554),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_13),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_326),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_281),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_294),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_128),
.Y(n_789)
);

CKINVDCx16_ASAP7_75t_R g790 ( 
.A(n_249),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_477),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_520),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_462),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_266),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_461),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_164),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_111),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_13),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_351),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_67),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_427),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_528),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_237),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_140),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_158),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_249),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_537),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_269),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_178),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_558),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_360),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_369),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_530),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_332),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_464),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_315),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_34),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_89),
.Y(n_818)
);

BUFx10_ASAP7_75t_L g819 ( 
.A(n_366),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_551),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_302),
.Y(n_821)
);

BUFx8_ASAP7_75t_SL g822 ( 
.A(n_153),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_209),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_433),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_99),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_271),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_55),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_393),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_279),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_570),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_534),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_454),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_470),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_508),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_46),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_590),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_705),
.Y(n_837)
);

INVxp33_ASAP7_75t_SL g838 ( 
.A(n_690),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_705),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_690),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_705),
.Y(n_841)
);

CKINVDCx14_ASAP7_75t_R g842 ( 
.A(n_634),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_705),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_705),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_705),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_705),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_822),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_650),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_621),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_822),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_621),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_646),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_638),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_750),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_657),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_638),
.Y(n_856)
);

INVxp33_ASAP7_75t_L g857 ( 
.A(n_626),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_768),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_813),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_768),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_646),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_646),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_646),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_589),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_657),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_591),
.Y(n_866)
);

INVxp33_ASAP7_75t_L g867 ( 
.A(n_644),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_593),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_834),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_598),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_602),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_603),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_605),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_612),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_623),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_588),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_600),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_625),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_628),
.Y(n_879)
);

INVxp33_ASAP7_75t_L g880 ( 
.A(n_653),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_834),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_750),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_629),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_633),
.Y(n_884)
);

BUFx5_ASAP7_75t_L g885 ( 
.A(n_596),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_639),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_640),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_696),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_641),
.Y(n_889)
);

INVxp67_ASAP7_75t_SL g890 ( 
.A(n_834),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_652),
.Y(n_891)
);

CKINVDCx14_ASAP7_75t_R g892 ( 
.A(n_634),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_663),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_665),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_790),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_668),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_669),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_673),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_666),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_674),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_684),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_750),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_704),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_706),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_685),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_747),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_747),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_707),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_700),
.B(n_0),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_750),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_710),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_711),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_716),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_718),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_720),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_750),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_750),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_728),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_731),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_736),
.Y(n_920)
);

CKINVDCx14_ASAP7_75t_R g921 ( 
.A(n_662),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_743),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_632),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_744),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_751),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_755),
.Y(n_926)
);

INVxp67_ASAP7_75t_SL g927 ( 
.A(n_599),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_606),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_666),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_758),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_666),
.Y(n_931)
);

CKINVDCx14_ASAP7_75t_R g932 ( 
.A(n_662),
.Y(n_932)
);

INVxp33_ASAP7_75t_SL g933 ( 
.A(n_587),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_760),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_661),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_761),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_757),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_888),
.A2(n_757),
.B1(n_759),
.B2(n_741),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_859),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_876),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_852),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_859),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_869),
.B(n_670),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_859),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_852),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_861),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_859),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_855),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_852),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_854),
.Y(n_950)
);

AND2x6_ASAP7_75t_L g951 ( 
.A(n_854),
.B(n_830),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_862),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_863),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_837),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_839),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_895),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_866),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_876),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_881),
.B(n_678),
.Y(n_959)
);

INVxp33_ASAP7_75t_SL g960 ( 
.A(n_855),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_841),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_868),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_933),
.B(n_759),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_843),
.A2(n_697),
.B(n_692),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_SL g965 ( 
.A1(n_847),
.A2(n_624),
.B1(n_635),
.B2(n_588),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_870),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_871),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_890),
.B(n_715),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_872),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_844),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_845),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_873),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_899),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_846),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_882),
.Y(n_975)
);

XOR2xp5_ASAP7_75t_L g976 ( 
.A(n_847),
.B(n_613),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_874),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_864),
.B(n_739),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_931),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_875),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_877),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_882),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_909),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_902),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_878),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_879),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_849),
.B(n_648),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_902),
.Y(n_988)
);

BUFx8_ASAP7_75t_SL g989 ( 
.A(n_850),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_928),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_910),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_865),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_842),
.B(n_752),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_923),
.Y(n_994)
);

AND2x6_ASAP7_75t_L g995 ( 
.A(n_910),
.B(n_830),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_885),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_916),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_883),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_916),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_884),
.Y(n_1000)
);

NOR2x1_ASAP7_75t_L g1001 ( 
.A(n_851),
.B(n_756),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_927),
.B(n_770),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_840),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_943),
.B(n_772),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_997),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_950),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_939),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_943),
.B(n_842),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_997),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_943),
.B(n_779),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_974),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_975),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_974),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_982),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_982),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_959),
.B(n_935),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_959),
.B(n_892),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_982),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_959),
.B(n_784),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_994),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_984),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_984),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_979),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_956),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_941),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_968),
.B(n_892),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_984),
.Y(n_1027)
);

AND3x2_ASAP7_75t_L g1028 ( 
.A(n_963),
.B(n_691),
.C(n_675),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_999),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_999),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_999),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_975),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_968),
.B(n_921),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_938),
.B(n_865),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_968),
.B(n_921),
.Y(n_1035)
);

BUFx8_ASAP7_75t_L g1036 ( 
.A(n_948),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_946),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_952),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_941),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_949),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_945),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_964),
.A2(n_917),
.B(n_820),
.Y(n_1042)
);

BUFx12f_ASAP7_75t_L g1043 ( 
.A(n_981),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_949),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_964),
.A2(n_917),
.B(n_792),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_939),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_975),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_939),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1002),
.B(n_978),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_953),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_975),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1002),
.B(n_932),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1002),
.B(n_932),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_954),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_987),
.B(n_836),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_945),
.B(n_886),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_954),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_954),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_954),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_954),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_955),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_955),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_939),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_975),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_987),
.B(n_848),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_993),
.B(n_907),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_955),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_988),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1001),
.B(n_887),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_988),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_983),
.B(n_853),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_988),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_955),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_983),
.B(n_957),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_939),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_988),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_944),
.B(n_906),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_942),
.A2(n_891),
.B(n_889),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_955),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_948),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_988),
.Y(n_1081)
);

INVx6_ASAP7_75t_L g1082 ( 
.A(n_991),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_940),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_961),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_962),
.B(n_856),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_961),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_991),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_944),
.B(n_906),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_961),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_961),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_961),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_970),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_991),
.Y(n_1093)
);

INVxp33_ASAP7_75t_L g1094 ( 
.A(n_1020),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1049),
.B(n_970),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_1025),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1078),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1014),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1014),
.Y(n_1099)
);

AND3x2_ASAP7_75t_L g1100 ( 
.A(n_1023),
.B(n_992),
.C(n_1003),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1056),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1016),
.B(n_1004),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1018),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1016),
.B(n_981),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1004),
.B(n_970),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1056),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1018),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1056),
.Y(n_1108)
);

OA21x2_ASAP7_75t_L g1109 ( 
.A1(n_1042),
.A2(n_947),
.B(n_942),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1004),
.B(n_990),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_1025),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1078),
.Y(n_1112)
);

INVx6_ASAP7_75t_L g1113 ( 
.A(n_1056),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_1025),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1023),
.B(n_992),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1037),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1071),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1037),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1038),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1038),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1078),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1022),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_R g1123 ( 
.A(n_1043),
.B(n_990),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1050),
.Y(n_1124)
);

AND3x1_ASAP7_75t_L g1125 ( 
.A(n_1074),
.B(n_973),
.C(n_860),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_SL g1126 ( 
.A1(n_1036),
.A2(n_624),
.B1(n_713),
.B2(n_635),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_1004),
.B(n_960),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_SL g1128 ( 
.A(n_1036),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1050),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1078),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1009),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1009),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1005),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1066),
.B(n_933),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1005),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_1006),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1055),
.B(n_973),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1085),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1085),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_SL g1140 ( 
.A(n_1069),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1055),
.B(n_857),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1039),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1010),
.B(n_1019),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1022),
.Y(n_1144)
);

OR2x6_ASAP7_75t_L g1145 ( 
.A(n_1043),
.B(n_965),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1074),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1010),
.B(n_960),
.Y(n_1147)
);

OAI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1052),
.A2(n_867),
.B1(n_880),
.B2(n_857),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1027),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1041),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1080),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1041),
.Y(n_1152)
);

NAND2xp33_ASAP7_75t_L g1153 ( 
.A(n_1053),
.B(n_750),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1065),
.B(n_907),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1010),
.B(n_970),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1011),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1010),
.B(n_970),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1041),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1019),
.B(n_971),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1027),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1019),
.A2(n_675),
.B1(n_712),
.B2(n_648),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1019),
.B(n_971),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1040),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1011),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1040),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1008),
.B(n_971),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1013),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1017),
.A2(n_741),
.B1(n_762),
.B2(n_613),
.Y(n_1169)
);

NOR2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1026),
.B(n_840),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1033),
.B(n_971),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1071),
.B(n_937),
.C(n_905),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1035),
.A2(n_766),
.B1(n_762),
.B2(n_937),
.Y(n_1173)
);

NAND2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1034),
.B(n_766),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_1079),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1044),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_1079),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1054),
.B(n_971),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1044),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1046),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1015),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1015),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1051),
.B(n_813),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1079),
.Y(n_1184)
);

BUFx4f_ASAP7_75t_L g1185 ( 
.A(n_1080),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1077),
.B(n_681),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1021),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1083),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1024),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1046),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1069),
.A2(n_754),
.B1(n_793),
.B2(n_712),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_1028),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1069),
.A2(n_793),
.B1(n_796),
.B2(n_754),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1006),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_1007),
.Y(n_1195)
);

INVx8_ASAP7_75t_L g1196 ( 
.A(n_1069),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1029),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1051),
.B(n_813),
.Y(n_1198)
);

INVx8_ASAP7_75t_L g1199 ( 
.A(n_1007),
.Y(n_1199)
);

AND2x6_ASAP7_75t_L g1200 ( 
.A(n_1064),
.B(n_813),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1082),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1030),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1064),
.B(n_830),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1030),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1082),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1082),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1054),
.B(n_991),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1082),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1031),
.Y(n_1209)
);

CKINVDCx16_ASAP7_75t_R g1210 ( 
.A(n_1088),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1031),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1070),
.B(n_830),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1070),
.Y(n_1213)
);

NAND2xp33_ASAP7_75t_SL g1214 ( 
.A(n_1072),
.B(n_681),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1072),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1076),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1012),
.Y(n_1217)
);

NAND2xp33_ASAP7_75t_R g1218 ( 
.A(n_1042),
.B(n_850),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1036),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1036),
.B(n_929),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1012),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1046),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1076),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1081),
.B(n_1093),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1012),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1081),
.B(n_867),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1093),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1057),
.B(n_991),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1012),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1131),
.Y(n_1230)
);

AO22x2_ASAP7_75t_L g1231 ( 
.A1(n_1169),
.A2(n_976),
.B1(n_622),
.B2(n_627),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1197),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1150),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1156),
.B(n_1057),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1150),
.Y(n_1235)
);

INVx5_ASAP7_75t_L g1236 ( 
.A(n_1180),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1131),
.Y(n_1237)
);

AND2x6_ASAP7_75t_L g1238 ( 
.A(n_1130),
.B(n_1058),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1188),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_1097),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1152),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1211),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1152),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1152),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1156),
.B(n_880),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1132),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1223),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1133),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1133),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1135),
.Y(n_1250)
);

OAI21xp33_ASAP7_75t_L g1251 ( 
.A1(n_1191),
.A2(n_767),
.B(n_763),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1135),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1151),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1191),
.A2(n_727),
.B1(n_764),
.B2(n_713),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1159),
.B(n_966),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1141),
.B(n_858),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1159),
.B(n_967),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1152),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1132),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1102),
.B(n_1058),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1146),
.B(n_1095),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1117),
.B(n_969),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1181),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1134),
.B(n_838),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1182),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1223),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1123),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1154),
.A2(n_1060),
.B1(n_1061),
.B2(n_1059),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1188),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1227),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1185),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1175),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1180),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1227),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1180),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1164),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1123),
.Y(n_1277)
);

NAND3x1_ASAP7_75t_L g1278 ( 
.A(n_1173),
.B(n_958),
.C(n_940),
.Y(n_1278)
);

INVx6_ASAP7_75t_L g1279 ( 
.A(n_1192),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1187),
.Y(n_1280)
);

AND2x6_ASAP7_75t_L g1281 ( 
.A(n_1097),
.B(n_1059),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1166),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1176),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1134),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1128),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1137),
.B(n_958),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1154),
.B(n_972),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1179),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1202),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1113),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1210),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1204),
.Y(n_1292)
);

INVx4_ASAP7_75t_SL g1293 ( 
.A(n_1113),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1101),
.B(n_977),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1175),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1226),
.B(n_980),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1185),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1106),
.B(n_985),
.Y(n_1298)
);

INVx4_ASAP7_75t_SL g1299 ( 
.A(n_1113),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1115),
.Y(n_1300)
);

AND2x6_ASAP7_75t_L g1301 ( 
.A(n_1112),
.B(n_1060),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1209),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1215),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1157),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1108),
.B(n_986),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1138),
.B(n_998),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1165),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1116),
.B(n_1061),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1215),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1098),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1099),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1180),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1103),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1139),
.B(n_1000),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1190),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1118),
.B(n_1119),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1177),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1104),
.B(n_838),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1189),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1193),
.A2(n_814),
.B1(n_833),
.B2(n_796),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1120),
.B(n_1062),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1107),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1143),
.A2(n_1067),
.B1(n_1073),
.B2(n_1062),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1168),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1122),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1142),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1144),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1193),
.A2(n_1162),
.B1(n_1174),
.B2(n_1186),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1124),
.Y(n_1329)
);

AO21x2_ASAP7_75t_L g1330 ( 
.A1(n_1167),
.A2(n_1045),
.B(n_1067),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1129),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1140),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1096),
.B(n_1032),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1125),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1149),
.Y(n_1335)
);

NOR2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1219),
.B(n_989),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1161),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1190),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1096),
.B(n_893),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1190),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1199),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1213),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1171),
.B(n_1073),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1162),
.A2(n_764),
.B1(n_786),
.B2(n_727),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1104),
.B(n_1084),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1216),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1111),
.B(n_894),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1177),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1190),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1217),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1221),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1174),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1111),
.B(n_896),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1222),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1222),
.Y(n_1355)
);

CKINVDCx16_ASAP7_75t_R g1356 ( 
.A(n_1128),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1199),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1229),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1105),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1155),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1192),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1160),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1222),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1112),
.B(n_1084),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1222),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1199),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1170),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1121),
.B(n_1195),
.Y(n_1368)
);

AND2x6_ASAP7_75t_L g1369 ( 
.A(n_1121),
.B(n_1086),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1094),
.B(n_773),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1153),
.B(n_1089),
.C(n_1086),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1126),
.A2(n_786),
.B1(n_808),
.B2(n_803),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1214),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1196),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1163),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1158),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1225),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1158),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1114),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1140),
.Y(n_1380)
);

AND2x6_ASAP7_75t_L g1381 ( 
.A(n_1184),
.B(n_1089),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1109),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1184),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1214),
.Y(n_1384)
);

INVx5_ASAP7_75t_L g1385 ( 
.A(n_1220),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1109),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1220),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1114),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1220),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_SL g1390 ( 
.A(n_1126),
.Y(n_1390)
);

BUFx10_ASAP7_75t_L g1391 ( 
.A(n_1100),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1195),
.B(n_1090),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1094),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1224),
.Y(n_1394)
);

AO22x2_ASAP7_75t_L g1395 ( 
.A1(n_1110),
.A2(n_694),
.B1(n_771),
.B2(n_619),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1110),
.B(n_1090),
.Y(n_1396)
);

AND2x2_ASAP7_75t_SL g1397 ( 
.A(n_1153),
.B(n_814),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1224),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1109),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1196),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1167),
.B(n_1091),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1225),
.B(n_1201),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1201),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1127),
.B(n_897),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1127),
.B(n_773),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1147),
.B(n_773),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1196),
.Y(n_1407)
);

NOR2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1172),
.B(n_989),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1205),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1205),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1206),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1206),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1207),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1208),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1208),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1228),
.Y(n_1416)
);

AND2x6_ASAP7_75t_L g1417 ( 
.A(n_1178),
.B(n_1091),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1147),
.B(n_1100),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1145),
.B(n_778),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1228),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1145),
.B(n_778),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1186),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1183),
.Y(n_1423)
);

INVx4_ASAP7_75t_L g1424 ( 
.A(n_1136),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1145),
.B(n_778),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1136),
.B(n_1092),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1148),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1183),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1198),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1287),
.B(n_1148),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1264),
.B(n_803),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1261),
.B(n_1032),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1253),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1270),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1248),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1407),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1274),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1261),
.B(n_1240),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1400),
.B(n_1293),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1230),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1284),
.B(n_1319),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1249),
.Y(n_1442)
);

BUFx4_ASAP7_75t_L g1443 ( 
.A(n_1356),
.Y(n_1443)
);

INVx5_ASAP7_75t_L g1444 ( 
.A(n_1273),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1237),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1373),
.A2(n_1218),
.B1(n_808),
.B2(n_777),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1284),
.B(n_1136),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1291),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1286),
.B(n_788),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1240),
.B(n_1032),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1293),
.B(n_1092),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1393),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1328),
.A2(n_1218),
.B1(n_1203),
.B2(n_1212),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1234),
.B(n_1296),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1246),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1267),
.B(n_819),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1328),
.A2(n_807),
.B1(n_782),
.B2(n_1198),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1234),
.B(n_1032),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1316),
.B(n_1047),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1376),
.A2(n_1378),
.B1(n_1316),
.B2(n_1396),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1373),
.A2(n_829),
.B1(n_776),
.B2(n_833),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1264),
.B(n_1047),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1300),
.B(n_1047),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1300),
.B(n_1047),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1393),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1273),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1250),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1279),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1345),
.A2(n_1212),
.B1(n_1203),
.B2(n_637),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1374),
.B(n_1068),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1256),
.B(n_1068),
.Y(n_1471)
);

AND2x6_ASAP7_75t_SL g1472 ( 
.A(n_1419),
.B(n_787),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1329),
.B(n_1068),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1331),
.B(n_1068),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1279),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1345),
.B(n_1087),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1259),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1252),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_R g1479 ( 
.A(n_1277),
.B(n_617),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1266),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1359),
.B(n_1087),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1427),
.A2(n_1087),
.B1(n_655),
.B2(n_659),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1339),
.B(n_1136),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1360),
.B(n_1087),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1362),
.B(n_642),
.Y(n_1485)
);

NOR2xp67_ASAP7_75t_L g1486 ( 
.A(n_1374),
.B(n_471),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1384),
.B(n_592),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1375),
.B(n_664),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1396),
.B(n_667),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1247),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1290),
.B(n_1194),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1245),
.B(n_898),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1247),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1245),
.B(n_819),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1304),
.B(n_679),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1307),
.B(n_698),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1377),
.A2(n_1194),
.B1(n_703),
.B2(n_709),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1422),
.A2(n_714),
.B1(n_723),
.B2(n_702),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1324),
.B(n_738),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1239),
.B(n_900),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1404),
.A2(n_1294),
.B1(n_1305),
.B2(n_1298),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1377),
.A2(n_1194),
.B1(n_745),
.B2(n_746),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1413),
.B(n_742),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1404),
.A2(n_765),
.B1(n_791),
.B2(n_748),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1384),
.B(n_594),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_SL g1506 ( 
.A(n_1391),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1339),
.B(n_1194),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1232),
.Y(n_1508)
);

NOR3xp33_ASAP7_75t_L g1509 ( 
.A(n_1372),
.B(n_903),
.C(n_901),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1242),
.B(n_1260),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1347),
.B(n_802),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1334),
.B(n_595),
.Y(n_1512)
);

NOR3xp33_ASAP7_75t_L g1513 ( 
.A(n_1372),
.B(n_908),
.C(n_904),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1276),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1334),
.B(n_597),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1318),
.B(n_601),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1308),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1352),
.A2(n_831),
.B1(n_810),
.B2(n_951),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1326),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1347),
.B(n_1007),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1260),
.B(n_604),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1370),
.B(n_819),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1318),
.B(n_1390),
.Y(n_1523)
);

NOR2xp67_ASAP7_75t_L g1524 ( 
.A(n_1341),
.B(n_472),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1368),
.B(n_607),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_SL g1526 ( 
.A(n_1297),
.B(n_1285),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1368),
.B(n_1306),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1308),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1321),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1263),
.A2(n_951),
.B1(n_995),
.B2(n_1200),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1405),
.B(n_911),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1282),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1269),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1353),
.B(n_608),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1273),
.Y(n_1535)
);

OR2x6_ASAP7_75t_L g1536 ( 
.A(n_1407),
.B(n_1045),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1353),
.B(n_609),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1314),
.B(n_1321),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1233),
.A2(n_1235),
.B1(n_1323),
.B2(n_1268),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1314),
.B(n_610),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1394),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1379),
.B(n_1007),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1379),
.B(n_1007),
.Y(n_1543)
);

AND2x6_ASAP7_75t_SL g1544 ( 
.A(n_1421),
.B(n_789),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1398),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1262),
.B(n_1294),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1406),
.B(n_912),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1275),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1262),
.B(n_611),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1342),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1283),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1298),
.B(n_614),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1305),
.B(n_615),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1390),
.B(n_616),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1265),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1288),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1255),
.A2(n_885),
.B1(n_1200),
.B2(n_1063),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1272),
.B(n_618),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1272),
.B(n_620),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1254),
.B(n_630),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1361),
.Y(n_1561)
);

NAND2x1_ASAP7_75t_L g1562 ( 
.A(n_1381),
.B(n_1046),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1407),
.B(n_913),
.Y(n_1563)
);

O2A1O1Ixp5_ASAP7_75t_L g1564 ( 
.A1(n_1343),
.A2(n_947),
.B(n_815),
.C(n_818),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1254),
.B(n_631),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1379),
.B(n_1063),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1346),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1388),
.B(n_1063),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1303),
.Y(n_1569)
);

AND2x6_ASAP7_75t_SL g1570 ( 
.A(n_1425),
.B(n_801),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1295),
.B(n_636),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1317),
.B(n_643),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1395),
.A2(n_885),
.B1(n_1200),
.B2(n_821),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1388),
.B(n_1063),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1395),
.A2(n_885),
.B1(n_1200),
.B2(n_915),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1243),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1233),
.A2(n_1048),
.B1(n_1075),
.B2(n_1046),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_SL g1578 ( 
.A(n_1344),
.B(n_645),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1293),
.B(n_1299),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1280),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1317),
.B(n_647),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1243),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1271),
.B(n_1418),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1289),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1344),
.B(n_914),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1302),
.A2(n_919),
.B(n_920),
.C(n_918),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1255),
.A2(n_885),
.B1(n_1200),
.B2(n_1063),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1257),
.B(n_922),
.Y(n_1588)
);

NOR2xp67_ASAP7_75t_L g1589 ( 
.A(n_1341),
.B(n_473),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1309),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1292),
.A2(n_885),
.B1(n_925),
.B2(n_924),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1388),
.B(n_1046),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1348),
.B(n_649),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1348),
.B(n_651),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1392),
.B(n_654),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1310),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1335),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1231),
.A2(n_885),
.B1(n_930),
.B2(n_926),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1231),
.A2(n_936),
.B1(n_934),
.B2(n_951),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1290),
.B(n_1257),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1311),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1392),
.B(n_656),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1268),
.B(n_658),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1364),
.B(n_660),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1397),
.A2(n_995),
.B1(n_951),
.B2(n_672),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1275),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1364),
.B(n_1416),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1420),
.B(n_671),
.Y(n_1608)
);

NOR3xp33_ASAP7_75t_L g1609 ( 
.A(n_1367),
.B(n_677),
.C(n_676),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1243),
.Y(n_1610)
);

OAI21xp33_ASAP7_75t_L g1611 ( 
.A1(n_1251),
.A2(n_682),
.B(n_680),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1323),
.A2(n_686),
.B(n_687),
.C(n_683),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1299),
.B(n_474),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1299),
.B(n_1048),
.Y(n_1614)
);

AND2x6_ASAP7_75t_L g1615 ( 
.A(n_1399),
.B(n_1048),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1332),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1244),
.B(n_688),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1275),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1332),
.B(n_689),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1244),
.B(n_693),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1244),
.B(n_695),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1385),
.A2(n_835),
.B1(n_701),
.B2(n_708),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1313),
.A2(n_995),
.B1(n_951),
.B2(n_717),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1385),
.B(n_475),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1322),
.A2(n_995),
.B1(n_951),
.B2(n_719),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1325),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1327),
.A2(n_995),
.B1(n_721),
.B2(n_722),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1337),
.A2(n_995),
.B1(n_724),
.B2(n_725),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1380),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1383),
.B(n_699),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1380),
.Y(n_1631)
);

INVx8_ASAP7_75t_L g1632 ( 
.A(n_1236),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1424),
.A2(n_996),
.B(n_950),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1387),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1433),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1579),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1561),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1517),
.B(n_1281),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1452),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1508),
.Y(n_1640)
);

AND2x2_ASAP7_75t_SL g1641 ( 
.A(n_1431),
.B(n_1320),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1439),
.B(n_1385),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1523),
.B(n_1391),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1632),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1634),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1465),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1528),
.B(n_1281),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1550),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1448),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1516),
.A2(n_1410),
.B1(n_1403),
.B2(n_1251),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1632),
.B(n_1563),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1435),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1500),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1579),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1613),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1449),
.B(n_1389),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1529),
.B(n_1281),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1434),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1554),
.B(n_1408),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1442),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1467),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1519),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1438),
.B(n_1281),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1468),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1583),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1527),
.B(n_1382),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1510),
.A2(n_1236),
.B(n_1424),
.Y(n_1667)
);

CKINVDCx11_ASAP7_75t_R g1668 ( 
.A(n_1472),
.Y(n_1668)
);

AND2x6_ASAP7_75t_SL g1669 ( 
.A(n_1560),
.B(n_1336),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1454),
.B(n_1386),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1588),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1531),
.B(n_1358),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1439),
.B(n_1546),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1475),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1478),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1437),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1547),
.B(n_1320),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1506),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1538),
.B(n_1301),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1533),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1501),
.B(n_1357),
.Y(n_1681)
);

OR2x6_ASAP7_75t_L g1682 ( 
.A(n_1632),
.B(n_1357),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1494),
.B(n_1350),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1607),
.B(n_1301),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1430),
.B(n_1351),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1541),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1565),
.A2(n_1414),
.B1(n_1238),
.B2(n_1412),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1522),
.B(n_1487),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1440),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1545),
.B(n_1460),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1555),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1525),
.B(n_1301),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_1631),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1521),
.B(n_1301),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1445),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1580),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1584),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1492),
.B(n_1414),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1616),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1444),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1629),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1466),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1597),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1455),
.Y(n_1704)
);

BUFx2_ASAP7_75t_SL g1705 ( 
.A(n_1436),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1613),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1477),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1604),
.B(n_1462),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1567),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1578),
.A2(n_1278),
.B1(n_1417),
.B2(n_1412),
.Y(n_1710)
);

AO22x1_ASAP7_75t_L g1711 ( 
.A1(n_1624),
.A2(n_1505),
.B1(n_1515),
.B2(n_1512),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1563),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1446),
.A2(n_1511),
.B1(n_1526),
.B2(n_1456),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1563),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1466),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1595),
.B(n_1369),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1443),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1601),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1617),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1626),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1619),
.B(n_1414),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1514),
.Y(n_1722)
);

NOR2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1585),
.B(n_1534),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1624),
.Y(n_1724)
);

NOR2xp67_ASAP7_75t_L g1725 ( 
.A(n_1620),
.B(n_1241),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1509),
.B(n_1423),
.Y(n_1726)
);

BUFx12f_ASAP7_75t_L g1727 ( 
.A(n_1544),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1532),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1466),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1490),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1535),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1551),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1556),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1596),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1602),
.B(n_1369),
.Y(n_1735)
);

OAI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1603),
.A2(n_1258),
.B1(n_1241),
.B2(n_1366),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1432),
.B(n_1369),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1609),
.A2(n_1417),
.B1(n_1409),
.B2(n_1415),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1463),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1457),
.A2(n_1236),
.B1(n_1315),
.B2(n_1312),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1576),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1436),
.B(n_1366),
.Y(n_1742)
);

NAND2x1_ASAP7_75t_L g1743 ( 
.A(n_1451),
.B(n_1381),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1480),
.Y(n_1744)
);

BUFx4f_ASAP7_75t_SL g1745 ( 
.A(n_1441),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1513),
.A2(n_1238),
.B1(n_1415),
.B2(n_1409),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1598),
.B(n_1549),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1540),
.B(n_1428),
.Y(n_1748)
);

INVx4_ASAP7_75t_L g1749 ( 
.A(n_1444),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1458),
.B(n_1369),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1459),
.B(n_1238),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1600),
.A2(n_1417),
.B1(n_1381),
.B2(n_1258),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1569),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1504),
.A2(n_1238),
.B1(n_1401),
.B2(n_1429),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1590),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1471),
.B(n_1381),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1493),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1473),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1474),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1489),
.B(n_1343),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1451),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1506),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1586),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1481),
.Y(n_1764)
);

INVxp33_ASAP7_75t_L g1765 ( 
.A(n_1479),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1484),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1622),
.B(n_1312),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1464),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1450),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1537),
.A2(n_1417),
.B1(n_1401),
.B2(n_1371),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1539),
.B(n_1312),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1630),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1535),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1476),
.B(n_1315),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1503),
.B(n_1411),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_L g1776 ( 
.A(n_1535),
.B(n_1338),
.Y(n_1776)
);

OR2x6_ASAP7_75t_L g1777 ( 
.A(n_1483),
.B(n_1315),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1482),
.A2(n_1371),
.B1(n_1411),
.B2(n_1426),
.Y(n_1778)
);

INVx5_ASAP7_75t_L g1779 ( 
.A(n_1615),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1576),
.Y(n_1780)
);

BUFx3_ASAP7_75t_L g1781 ( 
.A(n_1548),
.Y(n_1781)
);

AND3x2_ASAP7_75t_SL g1782 ( 
.A(n_1573),
.B(n_8),
.C(n_0),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1444),
.B(n_1338),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1536),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1608),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1582),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1548),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1485),
.B(n_1338),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1582),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1552),
.A2(n_1426),
.B1(n_729),
.B2(n_730),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1548),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1606),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1536),
.Y(n_1793)
);

INVx4_ASAP7_75t_L g1794 ( 
.A(n_1606),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1606),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1610),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1610),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1536),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1618),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1488),
.B(n_1340),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1618),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1618),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1453),
.B(n_1340),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1621),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1553),
.Y(n_1805)
);

BUFx4f_ASAP7_75t_SL g1806 ( 
.A(n_1447),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1562),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1495),
.B(n_1496),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1453),
.B(n_1340),
.Y(n_1809)
);

AND2x4_ASAP7_75t_L g1810 ( 
.A(n_1520),
.B(n_1349),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1558),
.A2(n_732),
.B1(n_733),
.B2(n_726),
.Y(n_1811)
);

NOR3xp33_ASAP7_75t_L g1812 ( 
.A(n_1461),
.B(n_735),
.C(n_734),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1499),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1612),
.B(n_1559),
.Y(n_1814)
);

INVxp67_ASAP7_75t_SL g1815 ( 
.A(n_1592),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1564),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1470),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1542),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1571),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1570),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1543),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1572),
.Y(n_1822)
);

BUFx2_ASAP7_75t_L g1823 ( 
.A(n_1581),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1593),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1594),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1566),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1599),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1708),
.A2(n_1507),
.B(n_1568),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1700),
.B(n_1486),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1808),
.B(n_1611),
.Y(n_1830)
);

A2O1A1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1641),
.A2(n_1518),
.B(n_1469),
.C(n_1575),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1648),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1688),
.B(n_1498),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1708),
.A2(n_1574),
.B(n_1577),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1645),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1640),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1785),
.B(n_1518),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1649),
.B(n_1486),
.Y(n_1838)
);

NOR2xp67_ASAP7_75t_SL g1839 ( 
.A(n_1727),
.B(n_1349),
.Y(n_1839)
);

NOR3xp33_ASAP7_75t_SL g1840 ( 
.A(n_1678),
.B(n_740),
.C(n_737),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1813),
.B(n_1469),
.Y(n_1841)
);

INVx4_ASAP7_75t_L g1842 ( 
.A(n_1700),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1719),
.B(n_1497),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1643),
.A2(n_1502),
.B(n_1614),
.C(n_1627),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1805),
.A2(n_1605),
.B(n_1524),
.C(n_1589),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1635),
.Y(n_1846)
);

NOR3xp33_ASAP7_75t_SL g1847 ( 
.A(n_1762),
.B(n_753),
.C(n_749),
.Y(n_1847)
);

AO22x1_ASAP7_75t_L g1848 ( 
.A1(n_1765),
.A2(n_774),
.B1(n_775),
.B2(n_769),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1719),
.B(n_1713),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1635),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1760),
.A2(n_1402),
.B(n_1524),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_SL g1852 ( 
.A1(n_1775),
.A2(n_1628),
.B(n_1530),
.C(n_1591),
.Y(n_1852)
);

O2A1O1Ixp5_ASAP7_75t_L g1853 ( 
.A1(n_1711),
.A2(n_1633),
.B(n_1615),
.C(n_1628),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1804),
.B(n_780),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1691),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1696),
.Y(n_1856)
);

XOR2x2_ASAP7_75t_L g1857 ( 
.A(n_1717),
.B(n_1),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1653),
.B(n_1354),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1671),
.B(n_1772),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1665),
.B(n_781),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1653),
.B(n_1354),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_L g1862 ( 
.A1(n_1814),
.A2(n_1491),
.B(n_1333),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1823),
.B(n_783),
.Y(n_1863)
);

XOR2xp5_ASAP7_75t_L g1864 ( 
.A(n_1659),
.B(n_1557),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1671),
.B(n_785),
.Y(n_1865)
);

O2A1O1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1767),
.A2(n_1333),
.B(n_1625),
.C(n_1623),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1699),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1665),
.B(n_794),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1685),
.B(n_795),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1697),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1672),
.B(n_797),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1703),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1814),
.A2(n_1355),
.B(n_1354),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1686),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_R g1875 ( 
.A(n_1637),
.B(n_1355),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1827),
.A2(n_1587),
.B1(n_1363),
.B2(n_1365),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1652),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1660),
.Y(n_1878)
);

OAI22xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1745),
.A2(n_799),
.B1(n_800),
.B2(n_798),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1661),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1639),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1812),
.A2(n_1330),
.B(n_805),
.C(n_806),
.Y(n_1882)
);

INVx2_ASAP7_75t_SL g1883 ( 
.A(n_1674),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1724),
.B(n_1363),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1690),
.A2(n_1365),
.B(n_1615),
.Y(n_1885)
);

A2O1A1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1819),
.A2(n_1530),
.B(n_1365),
.C(n_809),
.Y(n_1886)
);

OAI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1822),
.A2(n_812),
.B1(n_816),
.B2(n_811),
.C(n_804),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1721),
.Y(n_1888)
);

AO32x1_ASAP7_75t_L g1889 ( 
.A1(n_1740),
.A2(n_4),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1636),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1824),
.B(n_817),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1825),
.B(n_823),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1709),
.Y(n_1893)
);

O2A1O1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1723),
.A2(n_825),
.B(n_826),
.C(n_824),
.Y(n_1894)
);

O2A1O1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1726),
.A2(n_828),
.B(n_832),
.C(n_827),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1747),
.A2(n_1048),
.B1(n_1075),
.B2(n_950),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1656),
.A2(n_1075),
.B1(n_950),
.B2(n_4),
.Y(n_1897)
);

BUFx10_ASAP7_75t_L g1898 ( 
.A(n_1642),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1677),
.B(n_2),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1693),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1779),
.A2(n_1075),
.B(n_1006),
.Y(n_1901)
);

NAND2x1p5_ASAP7_75t_L g1902 ( 
.A(n_1749),
.B(n_1075),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1779),
.A2(n_577),
.B(n_575),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1683),
.B(n_3),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1701),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1748),
.B(n_5),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1770),
.A2(n_9),
.B(n_6),
.C(n_7),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1698),
.B(n_6),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_SL g1909 ( 
.A1(n_1820),
.A2(n_11),
.B1(n_7),
.B2(n_10),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_SL g1910 ( 
.A(n_1644),
.B(n_478),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1788),
.B(n_10),
.Y(n_1911)
);

NAND2x1p5_ASAP7_75t_L g1912 ( 
.A(n_1749),
.B(n_479),
.Y(n_1912)
);

A2O1A1Ixp33_ASAP7_75t_L g1913 ( 
.A1(n_1710),
.A2(n_14),
.B(n_11),
.C(n_12),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1636),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_R g1915 ( 
.A(n_1655),
.B(n_480),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1744),
.B(n_12),
.Y(n_1916)
);

NOR3xp33_ASAP7_75t_SL g1917 ( 
.A(n_1768),
.B(n_14),
.C(n_15),
.Y(n_1917)
);

AOI21x1_ASAP7_75t_L g1918 ( 
.A1(n_1771),
.A2(n_483),
.B(n_482),
.Y(n_1918)
);

NAND2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1644),
.B(n_484),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1680),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1675),
.Y(n_1921)
);

NAND2xp33_ASAP7_75t_SL g1922 ( 
.A(n_1636),
.B(n_15),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1673),
.B(n_16),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1673),
.B(n_16),
.Y(n_1924)
);

O2A1O1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1739),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1718),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1642),
.B(n_486),
.Y(n_1927)
);

INVx2_ASAP7_75t_SL g1928 ( 
.A(n_1664),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1720),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_1729),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1667),
.A2(n_581),
.B(n_580),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1788),
.B(n_17),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1704),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1730),
.B(n_18),
.Y(n_1934)
);

INVx5_ASAP7_75t_L g1935 ( 
.A(n_1682),
.Y(n_1935)
);

INVx4_ASAP7_75t_L g1936 ( 
.A(n_1682),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1739),
.B(n_19),
.Y(n_1937)
);

BUFx3_ASAP7_75t_L g1938 ( 
.A(n_1781),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_R g1939 ( 
.A(n_1655),
.B(n_487),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1771),
.A2(n_564),
.B(n_563),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1707),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1806),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1800),
.B(n_1646),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1728),
.B(n_20),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1800),
.B(n_1725),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1764),
.B(n_23),
.Y(n_1946)
);

O2A1O1Ixp33_ASAP7_75t_L g1947 ( 
.A1(n_1740),
.A2(n_1694),
.B(n_1662),
.C(n_1716),
.Y(n_1947)
);

NAND3xp33_ASAP7_75t_L g1948 ( 
.A(n_1811),
.B(n_23),
.C(n_24),
.Y(n_1948)
);

A2O1A1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1738),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1692),
.A2(n_578),
.B(n_573),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1722),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1712),
.B(n_489),
.Y(n_1952)
);

CKINVDCx8_ASAP7_75t_R g1953 ( 
.A(n_1669),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_SL g1954 ( 
.A(n_1651),
.B(n_490),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1763),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.C(n_29),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1706),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1956)
);

A2O1A1Ixp33_ASAP7_75t_L g1957 ( 
.A1(n_1694),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1787),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1714),
.B(n_492),
.Y(n_1959)
);

OAI21x1_ASAP7_75t_L g1960 ( 
.A1(n_1737),
.A2(n_496),
.B(n_495),
.Y(n_1960)
);

OAI21x1_ASAP7_75t_L g1961 ( 
.A1(n_1737),
.A2(n_499),
.B(n_497),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1706),
.B(n_501),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1732),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1692),
.A2(n_569),
.B(n_568),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1654),
.Y(n_1965)
);

O2A1O1Ixp33_ASAP7_75t_L g1966 ( 
.A1(n_1716),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1735),
.A2(n_586),
.B(n_585),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1766),
.B(n_35),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1790),
.B(n_1734),
.Y(n_1969)
);

A2O1A1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1735),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1751),
.A2(n_36),
.B(n_37),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1733),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1663),
.A2(n_582),
.B(n_503),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1755),
.B(n_502),
.Y(n_1974)
);

A2O1A1Ixp33_ASAP7_75t_SL g1975 ( 
.A1(n_1807),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1769),
.B(n_38),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1687),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1753),
.B(n_1757),
.Y(n_1978)
);

O2A1O1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1803),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1670),
.B(n_42),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1663),
.A2(n_509),
.B(n_504),
.Y(n_1981)
);

INVx2_ASAP7_75t_SL g1982 ( 
.A(n_1795),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1654),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1666),
.A2(n_512),
.B(n_511),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1666),
.A2(n_514),
.B(n_513),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1670),
.B(n_44),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1741),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1658),
.Y(n_1988)
);

OAI21xp33_ASAP7_75t_SL g1989 ( 
.A1(n_1638),
.A2(n_516),
.B(n_515),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1654),
.Y(n_1990)
);

O2A1O1Ixp5_ASAP7_75t_L g1991 ( 
.A1(n_1816),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1991)
);

OA21x2_ASAP7_75t_L g1992 ( 
.A1(n_1803),
.A2(n_519),
.B(n_518),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1702),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1679),
.A2(n_48),
.B(n_45),
.C(n_47),
.Y(n_1994)
);

INVxp67_ASAP7_75t_SL g1995 ( 
.A(n_1850),
.Y(n_1995)
);

AOI22xp33_ASAP7_75t_L g1996 ( 
.A1(n_1948),
.A2(n_1681),
.B1(n_1793),
.B2(n_1784),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1993),
.Y(n_1997)
);

NOR2x1_ASAP7_75t_R g1998 ( 
.A(n_1900),
.B(n_1668),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1993),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1836),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1930),
.Y(n_2001)
);

BUFx12f_ASAP7_75t_L g2002 ( 
.A(n_1898),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1943),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1935),
.B(n_1798),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1938),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1859),
.B(n_1676),
.Y(n_2006)
);

CKINVDCx14_ASAP7_75t_R g2007 ( 
.A(n_1888),
.Y(n_2007)
);

AOI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1849),
.A2(n_1681),
.B1(n_1651),
.B2(n_1736),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1935),
.B(n_1651),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1958),
.Y(n_2010)
);

OAI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1830),
.A2(n_1746),
.B1(n_1650),
.B2(n_1754),
.Y(n_2011)
);

BUFx2_ASAP7_75t_L g2012 ( 
.A(n_1987),
.Y(n_2012)
);

O2A1O1Ixp33_ASAP7_75t_L g2013 ( 
.A1(n_1907),
.A2(n_1679),
.B(n_1809),
.C(n_1647),
.Y(n_2013)
);

A2O1A1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1895),
.A2(n_1882),
.B(n_1894),
.C(n_1831),
.Y(n_2014)
);

CKINVDCx20_ASAP7_75t_R g2015 ( 
.A(n_1953),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1855),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1856),
.Y(n_2017)
);

A2O1A1Ixp33_ASAP7_75t_L g2018 ( 
.A1(n_1843),
.A2(n_1782),
.B(n_1752),
.C(n_1778),
.Y(n_2018)
);

INVxp67_ASAP7_75t_L g2019 ( 
.A(n_1881),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1837),
.B(n_1689),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1993),
.Y(n_2021)
);

BUFx6f_ASAP7_75t_L g2022 ( 
.A(n_1965),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1841),
.B(n_1758),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1980),
.B(n_1695),
.Y(n_2024)
);

BUFx12f_ASAP7_75t_L g2025 ( 
.A(n_1898),
.Y(n_2025)
);

AO21x2_ASAP7_75t_L g2026 ( 
.A1(n_1851),
.A2(n_1809),
.B(n_1751),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_1864),
.A2(n_1833),
.B1(n_1869),
.B2(n_1913),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1870),
.Y(n_2028)
);

BUFx3_ASAP7_75t_L g2029 ( 
.A(n_1835),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1986),
.B(n_1759),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1862),
.A2(n_1684),
.B(n_1776),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1832),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1846),
.B(n_1684),
.Y(n_2033)
);

NAND2x1p5_ASAP7_75t_L g2034 ( 
.A(n_1935),
.B(n_1742),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1872),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1937),
.B(n_1780),
.Y(n_2036)
);

OAI222xp33_ASAP7_75t_L g2037 ( 
.A1(n_1942),
.A2(n_1782),
.B1(n_1777),
.B2(n_1647),
.C1(n_1657),
.C2(n_1638),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_1945),
.B(n_1682),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1867),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_1883),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1874),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1936),
.B(n_1777),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1899),
.B(n_1797),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1936),
.B(n_1777),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1906),
.B(n_1774),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1891),
.A2(n_1761),
.B1(n_1742),
.B2(n_1705),
.Y(n_2046)
);

NAND2x1_ASAP7_75t_SL g2047 ( 
.A(n_1829),
.B(n_1799),
.Y(n_2047)
);

INVx4_ASAP7_75t_L g2048 ( 
.A(n_1965),
.Y(n_2048)
);

AO22x1_ASAP7_75t_L g2049 ( 
.A1(n_1971),
.A2(n_1815),
.B1(n_1802),
.B2(n_1817),
.Y(n_2049)
);

OAI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_1863),
.A2(n_1657),
.B1(n_1761),
.B2(n_1756),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1877),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1955),
.A2(n_1756),
.B1(n_1810),
.B2(n_1750),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1965),
.Y(n_2053)
);

BUFx8_ASAP7_75t_SL g2054 ( 
.A(n_1983),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1920),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1878),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1969),
.B(n_1774),
.Y(n_2057)
);

INVx3_ASAP7_75t_L g2058 ( 
.A(n_1983),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_1875),
.Y(n_2059)
);

HB1xp67_ASAP7_75t_L g2060 ( 
.A(n_1905),
.Y(n_2060)
);

INVx5_ASAP7_75t_L g2061 ( 
.A(n_1842),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1983),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_1990),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1880),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_1922),
.A2(n_1810),
.B1(n_1750),
.B2(n_1818),
.Y(n_2065)
);

BUFx2_ASAP7_75t_L g2066 ( 
.A(n_1990),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1890),
.B(n_1773),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1854),
.B(n_1871),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_SL g2069 ( 
.A1(n_1966),
.A2(n_1826),
.B(n_1821),
.Y(n_2069)
);

OR2x6_ASAP7_75t_L g2070 ( 
.A(n_1919),
.B(n_1743),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1932),
.B(n_1786),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1890),
.B(n_1773),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1990),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_1914),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1921),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1944),
.B(n_1801),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1982),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1926),
.Y(n_2078)
);

BUFx4_ASAP7_75t_SL g2079 ( 
.A(n_1916),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1893),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1952),
.B(n_1792),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_1928),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1914),
.B(n_1792),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_1884),
.Y(n_2084)
);

BUFx10_ASAP7_75t_L g2085 ( 
.A(n_1959),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1884),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1934),
.B(n_1789),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1909),
.A2(n_1796),
.B1(n_1794),
.B2(n_1715),
.Y(n_2088)
);

AND2x4_ASAP7_75t_L g2089 ( 
.A(n_1929),
.B(n_1794),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1923),
.B(n_1702),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1988),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_1858),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1838),
.B(n_1702),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1954),
.B(n_1845),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1933),
.Y(n_2095)
);

OR2x6_ASAP7_75t_L g2096 ( 
.A(n_1912),
.B(n_1783),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1941),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1976),
.B(n_1791),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1951),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1963),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_1927),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1972),
.Y(n_2102)
);

NOR2xp67_ASAP7_75t_L g2103 ( 
.A(n_1865),
.B(n_1715),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_1962),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1911),
.B(n_1791),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1927),
.Y(n_2106)
);

INVx3_ASAP7_75t_L g2107 ( 
.A(n_1962),
.Y(n_2107)
);

NAND2x1p5_ASAP7_75t_L g2108 ( 
.A(n_1842),
.B(n_1715),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1947),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_1917),
.A2(n_1791),
.B1(n_1731),
.B2(n_50),
.Y(n_2110)
);

A2O1A1Ixp33_ASAP7_75t_L g2111 ( 
.A1(n_1949),
.A2(n_1731),
.B(n_51),
.C(n_47),
.Y(n_2111)
);

BUFx4f_ASAP7_75t_L g2112 ( 
.A(n_1860),
.Y(n_2112)
);

BUFx8_ASAP7_75t_L g2113 ( 
.A(n_1868),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2003),
.B(n_2057),
.Y(n_2114)
);

OAI22xp33_ASAP7_75t_SL g2115 ( 
.A1(n_2094),
.A2(n_1956),
.B1(n_1910),
.B2(n_1977),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2091),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_1995),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2095),
.Y(n_2118)
);

O2A1O1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_2014),
.A2(n_1925),
.B(n_1994),
.C(n_1970),
.Y(n_2119)
);

INVx3_ASAP7_75t_SL g2120 ( 
.A(n_2059),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2000),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_2015),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2097),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2027),
.A2(n_1857),
.B1(n_1897),
.B2(n_1940),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2099),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_2068),
.B(n_2112),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2018),
.A2(n_1834),
.B(n_1885),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2000),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_2031),
.A2(n_1889),
.B(n_1873),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_2092),
.Y(n_2130)
);

NAND2x1p5_ASAP7_75t_L g2131 ( 
.A(n_2038),
.B(n_1839),
.Y(n_2131)
);

O2A1O1Ixp33_ASAP7_75t_SL g2132 ( 
.A1(n_2111),
.A2(n_1975),
.B(n_1957),
.C(n_1979),
.Y(n_2132)
);

A2O1A1Ixp33_ASAP7_75t_L g2133 ( 
.A1(n_2112),
.A2(n_1991),
.B(n_1853),
.C(n_1844),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2016),
.Y(n_2134)
);

OAI21xp33_ASAP7_75t_L g2135 ( 
.A1(n_2109),
.A2(n_1996),
.B(n_2023),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2100),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2011),
.A2(n_1974),
.B1(n_1924),
.B2(n_1887),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2033),
.B(n_1978),
.Y(n_2138)
);

O2A1O1Ixp33_ASAP7_75t_L g2139 ( 
.A1(n_2110),
.A2(n_1946),
.B(n_1968),
.C(n_1904),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_2109),
.A2(n_1985),
.B(n_1984),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_2085),
.B(n_1892),
.Y(n_2141)
);

O2A1O1Ixp33_ASAP7_75t_SL g2142 ( 
.A1(n_2093),
.A2(n_1861),
.B(n_1908),
.C(n_1886),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_2049),
.A2(n_1889),
.B(n_1828),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_2046),
.A2(n_1848),
.B1(n_1989),
.B2(n_1840),
.Y(n_2144)
);

INVx3_ASAP7_75t_SL g2145 ( 
.A(n_2001),
.Y(n_2145)
);

INVx2_ASAP7_75t_SL g2146 ( 
.A(n_2029),
.Y(n_2146)
);

NAND3xp33_ASAP7_75t_L g2147 ( 
.A(n_2050),
.B(n_1981),
.C(n_1973),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2045),
.B(n_1950),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_2085),
.B(n_1879),
.Y(n_2149)
);

AO21x1_ASAP7_75t_L g2150 ( 
.A1(n_2030),
.A2(n_1967),
.B(n_1964),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_2103),
.B(n_1915),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_SL g2152 ( 
.A1(n_2088),
.A2(n_1903),
.B(n_1931),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_L g2153 ( 
.A(n_2065),
.B(n_1847),
.C(n_1992),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_2008),
.B(n_2009),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2016),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2028),
.Y(n_2156)
);

OAI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_2013),
.A2(n_1961),
.B(n_1960),
.Y(n_2157)
);

BUFx10_ASAP7_75t_L g2158 ( 
.A(n_2005),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_2054),
.Y(n_2159)
);

AO31x2_ASAP7_75t_L g2160 ( 
.A1(n_2028),
.A2(n_1876),
.A3(n_1901),
.B(n_1889),
.Y(n_2160)
);

O2A1O1Ixp33_ASAP7_75t_L g2161 ( 
.A1(n_2037),
.A2(n_1852),
.B(n_1866),
.C(n_1992),
.Y(n_2161)
);

O2A1O1Ixp33_ASAP7_75t_SL g2162 ( 
.A1(n_2105),
.A2(n_1939),
.B(n_52),
.C(n_49),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2043),
.B(n_1918),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1997),
.Y(n_2164)
);

AND2x4_ASAP7_75t_L g2165 ( 
.A(n_2009),
.B(n_1731),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_2106),
.B(n_2104),
.Y(n_2166)
);

NOR2xp33_ASAP7_75t_SL g2167 ( 
.A(n_1998),
.B(n_1902),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_2026),
.A2(n_1896),
.B(n_524),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2041),
.Y(n_2169)
);

A2O1A1Ixp33_ASAP7_75t_L g2170 ( 
.A1(n_2101),
.A2(n_53),
.B(n_49),
.C(n_51),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2090),
.B(n_53),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2113),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2172)
);

OAI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_2024),
.A2(n_525),
.B(n_523),
.Y(n_2173)
);

OAI22x1_ASAP7_75t_L g2174 ( 
.A1(n_2012),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_L g2175 ( 
.A(n_1997),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_2007),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_2026),
.A2(n_529),
.B(n_526),
.Y(n_2177)
);

OAI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2052),
.A2(n_533),
.B(n_532),
.Y(n_2178)
);

BUFx6f_ASAP7_75t_L g2179 ( 
.A(n_1997),
.Y(n_2179)
);

BUFx10_ASAP7_75t_L g2180 ( 
.A(n_2010),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_2096),
.A2(n_536),
.B(n_535),
.Y(n_2181)
);

AO31x2_ASAP7_75t_L g2182 ( 
.A1(n_2051),
.A2(n_60),
.A3(n_58),
.B(n_59),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2051),
.Y(n_2183)
);

AOI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_2096),
.A2(n_541),
.B(n_540),
.Y(n_2184)
);

INVxp67_ASAP7_75t_SL g2185 ( 
.A(n_2117),
.Y(n_2185)
);

AOI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2124),
.A2(n_2113),
.B1(n_2106),
.B2(n_2107),
.Y(n_2186)
);

OAI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2178),
.A2(n_2106),
.B1(n_2070),
.B2(n_2104),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_2158),
.Y(n_2188)
);

AOI22xp33_ASAP7_75t_SL g2189 ( 
.A1(n_2115),
.A2(n_2107),
.B1(n_2044),
.B2(n_2042),
.Y(n_2189)
);

OAI21x1_ASAP7_75t_L g2190 ( 
.A1(n_2157),
.A2(n_2069),
.B(n_2034),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2114),
.B(n_2019),
.Y(n_2191)
);

AND2x4_ASAP7_75t_L g2192 ( 
.A(n_2130),
.B(n_2121),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2118),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2163),
.B(n_2039),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_2154),
.A2(n_2081),
.B1(n_2042),
.B2(n_2044),
.Y(n_2195)
);

CKINVDCx6p67_ASAP7_75t_R g2196 ( 
.A(n_2120),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_2122),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2128),
.Y(n_2198)
);

AOI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2137),
.A2(n_2036),
.B1(n_2098),
.B2(n_2076),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2123),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2172),
.A2(n_2060),
.B1(n_2071),
.B2(n_2020),
.Y(n_2201)
);

INVx8_ASAP7_75t_L g2202 ( 
.A(n_2159),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2134),
.B(n_2056),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2125),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2155),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2119),
.A2(n_2006),
.B1(n_2035),
.B2(n_2017),
.Y(n_2206)
);

BUFx5_ASAP7_75t_L g2207 ( 
.A(n_2156),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_2158),
.Y(n_2208)
);

AO22x1_ASAP7_75t_L g2209 ( 
.A1(n_2126),
.A2(n_2061),
.B1(n_2078),
.B2(n_2089),
.Y(n_2209)
);

OAI21x1_ASAP7_75t_L g2210 ( 
.A1(n_2129),
.A2(n_2102),
.B(n_2064),
.Y(n_2210)
);

BUFx2_ASAP7_75t_L g2211 ( 
.A(n_2176),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2136),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2169),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2183),
.B(n_2056),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2116),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2182),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2182),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2182),
.Y(n_2218)
);

INVx4_ASAP7_75t_SL g2219 ( 
.A(n_2145),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_2153),
.A2(n_2004),
.B1(n_2070),
.B2(n_2084),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_2180),
.Y(n_2221)
);

AOI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_2147),
.A2(n_2004),
.B1(n_2025),
.B2(n_2002),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_2127),
.A2(n_2061),
.B(n_2089),
.Y(n_2223)
);

AOI221xp5_ASAP7_75t_L g2224 ( 
.A1(n_2174),
.A2(n_2087),
.B1(n_2082),
.B2(n_2064),
.C(n_2075),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_SL g2225 ( 
.A1(n_2140),
.A2(n_2061),
.B1(n_2055),
.B2(n_2074),
.Y(n_2225)
);

OAI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2133),
.A2(n_2047),
.B(n_2032),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2141),
.A2(n_2040),
.B1(n_2077),
.B2(n_2086),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_L g2228 ( 
.A1(n_2135),
.A2(n_2086),
.B1(n_2066),
.B2(n_2063),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2164),
.Y(n_2229)
);

OAI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2144),
.A2(n_2086),
.B1(n_2075),
.B2(n_2048),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2138),
.B(n_2080),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2148),
.B(n_2053),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2192),
.B(n_2146),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2198),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2207),
.Y(n_2235)
);

INVxp67_ASAP7_75t_SL g2236 ( 
.A(n_2185),
.Y(n_2236)
);

INVx4_ASAP7_75t_L g2237 ( 
.A(n_2219),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2205),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2213),
.Y(n_2239)
);

INVx4_ASAP7_75t_SL g2240 ( 
.A(n_2216),
.Y(n_2240)
);

AOI21x1_ASAP7_75t_L g2241 ( 
.A1(n_2209),
.A2(n_2143),
.B(n_2177),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2207),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2194),
.B(n_2160),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2214),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2192),
.B(n_2166),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2214),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2203),
.Y(n_2247)
);

OAI21x1_ASAP7_75t_L g2248 ( 
.A1(n_2210),
.A2(n_2161),
.B(n_2168),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2191),
.B(n_2180),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2232),
.B(n_2171),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2215),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2211),
.B(n_2160),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2217),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2207),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2207),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2218),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2207),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2193),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2200),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2204),
.Y(n_2260)
);

INVxp67_ASAP7_75t_L g2261 ( 
.A(n_2244),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_SL g2262 ( 
.A1(n_2237),
.A2(n_2201),
.B1(n_2206),
.B2(n_2223),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_2237),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2244),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2246),
.B(n_2245),
.Y(n_2265)
);

BUFx2_ASAP7_75t_L g2266 ( 
.A(n_2237),
.Y(n_2266)
);

OAI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2241),
.A2(n_2206),
.B1(n_2199),
.B2(n_2230),
.Y(n_2267)
);

AOI21xp5_ASAP7_75t_L g2268 ( 
.A1(n_2248),
.A2(n_2132),
.B(n_2142),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2247),
.B(n_2212),
.Y(n_2269)
);

AOI222xp33_ASAP7_75t_L g2270 ( 
.A1(n_2236),
.A2(n_2201),
.B1(n_2224),
.B2(n_2170),
.C1(n_2226),
.C2(n_2220),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_2249),
.A2(n_2189),
.B1(n_2150),
.B2(n_2187),
.Y(n_2271)
);

AOI222xp33_ASAP7_75t_L g2272 ( 
.A1(n_2250),
.A2(n_2226),
.B1(n_2149),
.B2(n_2152),
.C1(n_2186),
.C2(n_2173),
.Y(n_2272)
);

HB1xp67_ASAP7_75t_L g2273 ( 
.A(n_2261),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2262),
.A2(n_2225),
.B1(n_2222),
.B2(n_2195),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2270),
.B(n_2252),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2269),
.Y(n_2276)
);

OAI221xp5_ASAP7_75t_L g2277 ( 
.A1(n_2268),
.A2(n_2199),
.B1(n_2227),
.B2(n_2243),
.C(n_2228),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2266),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2265),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_2263),
.Y(n_2280)
);

NOR4xp25_ASAP7_75t_L g2281 ( 
.A(n_2275),
.B(n_2278),
.C(n_2267),
.D(n_2277),
.Y(n_2281)
);

AOI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2274),
.A2(n_2272),
.B1(n_2271),
.B2(n_2248),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2279),
.A2(n_2265),
.B1(n_2167),
.B2(n_2252),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2273),
.Y(n_2284)
);

NAND4xp25_ASAP7_75t_L g2285 ( 
.A(n_2276),
.B(n_2139),
.C(n_2162),
.D(n_2232),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2280),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2280),
.Y(n_2287)
);

OAI31xp33_ASAP7_75t_L g2288 ( 
.A1(n_2280),
.A2(n_2131),
.A3(n_2243),
.B(n_2249),
.Y(n_2288)
);

OAI31xp33_ASAP7_75t_L g2289 ( 
.A1(n_2274),
.A2(n_2245),
.A3(n_2233),
.B(n_2264),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2273),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2284),
.B(n_2246),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2290),
.Y(n_2292)
);

BUFx3_ASAP7_75t_L g2293 ( 
.A(n_2286),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2287),
.B(n_2219),
.Y(n_2294)
);

AOI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2282),
.A2(n_2202),
.B(n_2197),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2283),
.B(n_2196),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2285),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2288),
.B(n_2289),
.Y(n_2298)
);

BUFx2_ASAP7_75t_L g2299 ( 
.A(n_2281),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2282),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2284),
.B(n_2233),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2284),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2293),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2292),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2302),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2299),
.B(n_2202),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2294),
.B(n_2188),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2294),
.B(n_2221),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2299),
.B(n_2269),
.Y(n_2309)
);

OAI21x1_ASAP7_75t_SL g2310 ( 
.A1(n_2295),
.A2(n_2241),
.B(n_2202),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_2293),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2311),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_2306),
.B(n_2297),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2311),
.Y(n_2314)
);

INVx2_ASAP7_75t_SL g2315 ( 
.A(n_2311),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2315),
.B(n_2303),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2314),
.B(n_2307),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_2312),
.B(n_2309),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2313),
.B(n_2308),
.Y(n_2319)
);

INVx1_ASAP7_75t_SL g2320 ( 
.A(n_2318),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2317),
.B(n_2306),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2319),
.B(n_2303),
.Y(n_2322)
);

NAND2x1p5_ASAP7_75t_L g2323 ( 
.A(n_2316),
.B(n_2304),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2316),
.B(n_2296),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2316),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2325),
.B(n_2297),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2322),
.B(n_2321),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2323),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2323),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2324),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2320),
.B(n_2296),
.Y(n_2331)
);

NOR2xp67_ASAP7_75t_SL g2332 ( 
.A(n_2320),
.B(n_2305),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2323),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2320),
.B(n_2300),
.Y(n_2334)
);

INVxp67_ASAP7_75t_L g2335 ( 
.A(n_2325),
.Y(n_2335)
);

AOI221xp5_ASAP7_75t_L g2336 ( 
.A1(n_2332),
.A2(n_2300),
.B1(n_2298),
.B2(n_2310),
.C(n_2291),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2328),
.B(n_2329),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2327),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2333),
.A2(n_2298),
.B(n_2301),
.Y(n_2339)
);

AOI21xp5_ASAP7_75t_L g2340 ( 
.A1(n_2334),
.A2(n_2301),
.B(n_2291),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_SL g2341 ( 
.A1(n_2326),
.A2(n_2151),
.B(n_2181),
.Y(n_2341)
);

NAND2x1p5_ASAP7_75t_L g2342 ( 
.A(n_2331),
.B(n_2208),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2335),
.A2(n_2208),
.B(n_2184),
.Y(n_2343)
);

AOI21xp5_ASAP7_75t_L g2344 ( 
.A1(n_2326),
.A2(n_2231),
.B(n_2253),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2330),
.B(n_2245),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2327),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2331),
.B(n_2247),
.Y(n_2347)
);

HB1xp67_ASAP7_75t_L g2348 ( 
.A(n_2328),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2348),
.Y(n_2349)
);

OAI321xp33_ASAP7_75t_L g2350 ( 
.A1(n_2337),
.A2(n_2108),
.A3(n_2231),
.B1(n_2256),
.B2(n_2253),
.C(n_2021),
.Y(n_2350)
);

AOI332xp33_ASAP7_75t_L g2351 ( 
.A1(n_2338),
.A2(n_2256),
.A3(n_63),
.B1(n_60),
.B2(n_64),
.B3(n_62),
.C1(n_58),
.C2(n_59),
.Y(n_2351)
);

OR2x2_ASAP7_75t_L g2352 ( 
.A(n_2340),
.B(n_2251),
.Y(n_2352)
);

AOI21xp33_ASAP7_75t_SL g2353 ( 
.A1(n_2342),
.A2(n_61),
.B(n_62),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2345),
.Y(n_2354)
);

INVx2_ASAP7_75t_SL g2355 ( 
.A(n_2347),
.Y(n_2355)
);

NOR2x1_ASAP7_75t_L g2356 ( 
.A(n_2346),
.B(n_61),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2339),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2336),
.B(n_2343),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2341),
.B(n_65),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2344),
.B(n_2251),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2339),
.B(n_2234),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2337),
.B(n_65),
.Y(n_2362)
);

AOI321xp33_ASAP7_75t_L g2363 ( 
.A1(n_2337),
.A2(n_2079),
.A3(n_2165),
.B1(n_2083),
.B2(n_2072),
.C(n_2067),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2356),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2349),
.B(n_2234),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2357),
.B(n_66),
.Y(n_2366)
);

XNOR2x1_ASAP7_75t_L g2367 ( 
.A(n_2354),
.B(n_2358),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_2355),
.B(n_67),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2362),
.B(n_2240),
.Y(n_2369)
);

XNOR2x1_ASAP7_75t_L g2370 ( 
.A(n_2352),
.B(n_68),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2361),
.Y(n_2371)
);

INVx1_ASAP7_75t_SL g2372 ( 
.A(n_2359),
.Y(n_2372)
);

AOI322xp5_ASAP7_75t_L g2373 ( 
.A1(n_2360),
.A2(n_2229),
.A3(n_2238),
.B1(n_2239),
.B2(n_2254),
.C1(n_2242),
.C2(n_2235),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2351),
.A2(n_2240),
.B1(n_2238),
.B2(n_2239),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2353),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2363),
.B(n_2258),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2350),
.Y(n_2377)
);

INVx2_ASAP7_75t_SL g2378 ( 
.A(n_2364),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2375),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2368),
.Y(n_2380)
);

INVxp67_ASAP7_75t_L g2381 ( 
.A(n_2366),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2377),
.A2(n_2240),
.B1(n_2242),
.B2(n_2235),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2370),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2367),
.Y(n_2384)
);

XOR2x2_ASAP7_75t_L g2385 ( 
.A(n_2372),
.B(n_2371),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2369),
.Y(n_2386)
);

AO22x2_ASAP7_75t_L g2387 ( 
.A1(n_2365),
.A2(n_2240),
.B1(n_71),
.B2(n_69),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2374),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2376),
.B(n_2258),
.Y(n_2389)
);

NOR2x1_ASAP7_75t_L g2390 ( 
.A(n_2373),
.B(n_70),
.Y(n_2390)
);

NOR3xp33_ASAP7_75t_L g2391 ( 
.A(n_2375),
.B(n_2048),
.C(n_70),
.Y(n_2391)
);

INVx1_ASAP7_75t_SL g2392 ( 
.A(n_2364),
.Y(n_2392)
);

INVx1_ASAP7_75t_SL g2393 ( 
.A(n_2364),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2364),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2374),
.A2(n_2255),
.B1(n_2257),
.B2(n_2254),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2364),
.Y(n_2396)
);

AOI211xp5_ASAP7_75t_SL g2397 ( 
.A1(n_2375),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_2397)
);

OR2x2_ASAP7_75t_L g2398 ( 
.A(n_2364),
.B(n_72),
.Y(n_2398)
);

NOR2xp33_ASAP7_75t_L g2399 ( 
.A(n_2375),
.B(n_73),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2378),
.B(n_2392),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2398),
.B(n_74),
.Y(n_2401)
);

NOR3xp33_ASAP7_75t_L g2402 ( 
.A(n_2384),
.B(n_74),
.C(n_75),
.Y(n_2402)
);

NOR3xp33_ASAP7_75t_L g2403 ( 
.A(n_2379),
.B(n_75),
.C(n_76),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2393),
.B(n_77),
.Y(n_2404)
);

NAND5xp2_ASAP7_75t_L g2405 ( 
.A(n_2383),
.B(n_79),
.C(n_77),
.D(n_78),
.E(n_80),
.Y(n_2405)
);

NOR2xp33_ASAP7_75t_L g2406 ( 
.A(n_2386),
.B(n_78),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2399),
.Y(n_2407)
);

NOR2xp67_ASAP7_75t_L g2408 ( 
.A(n_2394),
.B(n_80),
.Y(n_2408)
);

NOR3xp33_ASAP7_75t_L g2409 ( 
.A(n_2388),
.B(n_81),
.C(n_82),
.Y(n_2409)
);

AOI221xp5_ASAP7_75t_L g2410 ( 
.A1(n_2395),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.C(n_84),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2396),
.Y(n_2411)
);

NOR2x1_ASAP7_75t_L g2412 ( 
.A(n_2380),
.B(n_83),
.Y(n_2412)
);

NOR2x1_ASAP7_75t_L g2413 ( 
.A(n_2390),
.B(n_84),
.Y(n_2413)
);

NAND4xp25_ASAP7_75t_L g2414 ( 
.A(n_2391),
.B(n_87),
.C(n_85),
.D(n_86),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2381),
.B(n_85),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2385),
.Y(n_2416)
);

NAND4xp25_ASAP7_75t_L g2417 ( 
.A(n_2397),
.B(n_88),
.C(n_86),
.D(n_87),
.Y(n_2417)
);

NAND3xp33_ASAP7_75t_L g2418 ( 
.A(n_2382),
.B(n_2389),
.C(n_2387),
.Y(n_2418)
);

OAI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2387),
.A2(n_2260),
.B1(n_2259),
.B2(n_2257),
.C(n_2255),
.Y(n_2419)
);

OAI211xp5_ASAP7_75t_SL g2420 ( 
.A1(n_2379),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_2420)
);

NOR2x1_ASAP7_75t_L g2421 ( 
.A(n_2398),
.B(n_90),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2397),
.B(n_91),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_L g2423 ( 
.A(n_2391),
.B(n_92),
.C(n_93),
.Y(n_2423)
);

NAND2x1p5_ASAP7_75t_L g2424 ( 
.A(n_2392),
.B(n_1999),
.Y(n_2424)
);

OAI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2382),
.A2(n_2021),
.B1(n_1999),
.B2(n_2260),
.Y(n_2425)
);

NOR4xp25_ASAP7_75t_L g2426 ( 
.A(n_2392),
.B(n_94),
.C(n_92),
.D(n_93),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_2379),
.B(n_2165),
.Y(n_2427)
);

NOR3x1_ASAP7_75t_L g2428 ( 
.A(n_2378),
.B(n_94),
.C(n_95),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2398),
.Y(n_2429)
);

INVxp67_ASAP7_75t_SL g2430 ( 
.A(n_2398),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2378),
.Y(n_2431)
);

NAND3xp33_ASAP7_75t_L g2432 ( 
.A(n_2391),
.B(n_95),
.C(n_96),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2398),
.Y(n_2433)
);

NOR4xp25_ASAP7_75t_L g2434 ( 
.A(n_2392),
.B(n_98),
.C(n_96),
.D(n_97),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2397),
.B(n_97),
.Y(n_2435)
);

NOR3xp33_ASAP7_75t_L g2436 ( 
.A(n_2384),
.B(n_98),
.C(n_99),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2412),
.Y(n_2437)
);

AOI211x1_ASAP7_75t_L g2438 ( 
.A1(n_2400),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_2438)
);

AOI221x1_ASAP7_75t_SL g2439 ( 
.A1(n_2418),
.A2(n_2416),
.B1(n_2411),
.B2(n_2427),
.C(n_2429),
.Y(n_2439)
);

AOI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_2430),
.A2(n_100),
.B(n_101),
.Y(n_2440)
);

XNOR2xp5_ASAP7_75t_L g2441 ( 
.A(n_2417),
.B(n_102),
.Y(n_2441)
);

AOI211xp5_ASAP7_75t_SL g2442 ( 
.A1(n_2406),
.A2(n_106),
.B(n_103),
.C(n_105),
.Y(n_2442)
);

AOI31xp33_ASAP7_75t_L g2443 ( 
.A1(n_2422),
.A2(n_108),
.A3(n_105),
.B(n_107),
.Y(n_2443)
);

A2O1A1Ixp33_ASAP7_75t_L g2444 ( 
.A1(n_2408),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2435),
.Y(n_2445)
);

AOI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2431),
.A2(n_2021),
.B1(n_1999),
.B2(n_2022),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2401),
.Y(n_2447)
);

OAI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2404),
.A2(n_2190),
.B(n_2259),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2421),
.Y(n_2449)
);

O2A1O1Ixp5_ASAP7_75t_L g2450 ( 
.A1(n_2433),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_2450)
);

AOI211xp5_ASAP7_75t_L g2451 ( 
.A1(n_2426),
.A2(n_113),
.B(n_110),
.C(n_112),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2405),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2428),
.Y(n_2453)
);

AOI21xp33_ASAP7_75t_L g2454 ( 
.A1(n_2415),
.A2(n_112),
.B(n_113),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2431),
.Y(n_2455)
);

NOR2xp67_ASAP7_75t_L g2456 ( 
.A(n_2414),
.B(n_115),
.Y(n_2456)
);

NOR3xp33_ASAP7_75t_L g2457 ( 
.A(n_2407),
.B(n_2432),
.C(n_2423),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2413),
.A2(n_115),
.B(n_116),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2424),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2420),
.Y(n_2460)
);

OAI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_2409),
.A2(n_116),
.B(n_117),
.Y(n_2461)
);

AO221x1_ASAP7_75t_L g2462 ( 
.A1(n_2425),
.A2(n_2175),
.B1(n_2179),
.B2(n_2164),
.C(n_2022),
.Y(n_2462)
);

AOI21xp33_ASAP7_75t_L g2463 ( 
.A1(n_2410),
.A2(n_117),
.B(n_119),
.Y(n_2463)
);

O2A1O1Ixp33_ASAP7_75t_L g2464 ( 
.A1(n_2434),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_2464)
);

OAI21xp33_ASAP7_75t_L g2465 ( 
.A1(n_2402),
.A2(n_2058),
.B(n_2053),
.Y(n_2465)
);

NAND2x1p5_ASAP7_75t_L g2466 ( 
.A(n_2436),
.B(n_2022),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2403),
.B(n_120),
.Y(n_2467)
);

NOR2x1_ASAP7_75t_L g2468 ( 
.A(n_2419),
.B(n_121),
.Y(n_2468)
);

AOI22x1_ASAP7_75t_L g2469 ( 
.A1(n_2424),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2469)
);

AOI321xp33_ASAP7_75t_L g2470 ( 
.A1(n_2400),
.A2(n_124),
.A3(n_126),
.B1(n_122),
.B2(n_123),
.C(n_125),
.Y(n_2470)
);

NAND3xp33_ASAP7_75t_L g2471 ( 
.A(n_2409),
.B(n_125),
.C(n_126),
.Y(n_2471)
);

NOR3xp33_ASAP7_75t_SL g2472 ( 
.A(n_2400),
.B(n_127),
.C(n_128),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2417),
.B(n_127),
.Y(n_2473)
);

XOR2x2_ASAP7_75t_L g2474 ( 
.A(n_2413),
.B(n_129),
.Y(n_2474)
);

NOR2x1_ASAP7_75t_L g2475 ( 
.A(n_2437),
.B(n_129),
.Y(n_2475)
);

NOR3xp33_ASAP7_75t_L g2476 ( 
.A(n_2443),
.B(n_130),
.C(n_131),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_2452),
.B(n_130),
.Y(n_2477)
);

NOR3x1_ASAP7_75t_L g2478 ( 
.A(n_2471),
.B(n_131),
.C(n_132),
.Y(n_2478)
);

HB1xp67_ASAP7_75t_L g2479 ( 
.A(n_2474),
.Y(n_2479)
);

NOR2xp67_ASAP7_75t_L g2480 ( 
.A(n_2447),
.B(n_132),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2473),
.B(n_133),
.Y(n_2481)
);

NOR3xp33_ASAP7_75t_L g2482 ( 
.A(n_2449),
.B(n_133),
.C(n_136),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2441),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2472),
.B(n_136),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_2469),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2438),
.Y(n_2486)
);

NAND4xp25_ASAP7_75t_L g2487 ( 
.A(n_2439),
.B(n_139),
.C(n_137),
.D(n_138),
.Y(n_2487)
);

AOI211xp5_ASAP7_75t_L g2488 ( 
.A1(n_2463),
.A2(n_2464),
.B(n_2461),
.C(n_2458),
.Y(n_2488)
);

NAND4xp75_ASAP7_75t_L g2489 ( 
.A(n_2438),
.B(n_139),
.C(n_137),
.D(n_138),
.Y(n_2489)
);

OR3x2_ASAP7_75t_L g2490 ( 
.A(n_2453),
.B(n_141),
.C(n_142),
.Y(n_2490)
);

NOR2x1_ASAP7_75t_L g2491 ( 
.A(n_2444),
.B(n_141),
.Y(n_2491)
);

HB1xp67_ASAP7_75t_L g2492 ( 
.A(n_2456),
.Y(n_2492)
);

NOR2x1_ASAP7_75t_L g2493 ( 
.A(n_2459),
.B(n_142),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_SL g2494 ( 
.A(n_2470),
.B(n_2164),
.Y(n_2494)
);

NOR3xp33_ASAP7_75t_SL g2495 ( 
.A(n_2460),
.B(n_143),
.C(n_144),
.Y(n_2495)
);

AO22x1_ASAP7_75t_L g2496 ( 
.A1(n_2467),
.A2(n_2455),
.B1(n_2457),
.B2(n_2468),
.Y(n_2496)
);

NAND3xp33_ASAP7_75t_L g2497 ( 
.A(n_2451),
.B(n_145),
.C(n_146),
.Y(n_2497)
);

BUFx4f_ASAP7_75t_SL g2498 ( 
.A(n_2445),
.Y(n_2498)
);

NAND3xp33_ASAP7_75t_L g2499 ( 
.A(n_2442),
.B(n_145),
.C(n_147),
.Y(n_2499)
);

OR2x2_ASAP7_75t_L g2500 ( 
.A(n_2466),
.B(n_147),
.Y(n_2500)
);

NAND4xp25_ASAP7_75t_L g2501 ( 
.A(n_2450),
.B(n_150),
.C(n_148),
.D(n_149),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2440),
.Y(n_2502)
);

NOR3xp33_ASAP7_75t_L g2503 ( 
.A(n_2454),
.B(n_148),
.C(n_149),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2465),
.B(n_150),
.Y(n_2504)
);

NOR3xp33_ASAP7_75t_SL g2505 ( 
.A(n_2448),
.B(n_151),
.C(n_152),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2462),
.B(n_152),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2446),
.B(n_153),
.Y(n_2507)
);

INVx2_ASAP7_75t_SL g2508 ( 
.A(n_2474),
.Y(n_2508)
);

NOR2x1_ASAP7_75t_L g2509 ( 
.A(n_2437),
.B(n_154),
.Y(n_2509)
);

NAND3xp33_ASAP7_75t_L g2510 ( 
.A(n_2438),
.B(n_154),
.C(n_155),
.Y(n_2510)
);

NAND3x1_ASAP7_75t_L g2511 ( 
.A(n_2437),
.B(n_155),
.C(n_156),
.Y(n_2511)
);

XNOR2xp5_ASAP7_75t_L g2512 ( 
.A(n_2439),
.B(n_156),
.Y(n_2512)
);

NOR2x1_ASAP7_75t_L g2513 ( 
.A(n_2437),
.B(n_157),
.Y(n_2513)
);

NAND2x1p5_ASAP7_75t_L g2514 ( 
.A(n_2447),
.B(n_2058),
.Y(n_2514)
);

HB1xp67_ASAP7_75t_L g2515 ( 
.A(n_2474),
.Y(n_2515)
);

NOR2x1_ASAP7_75t_L g2516 ( 
.A(n_2437),
.B(n_157),
.Y(n_2516)
);

NOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2437),
.B(n_158),
.Y(n_2517)
);

NOR2x1_ASAP7_75t_L g2518 ( 
.A(n_2437),
.B(n_159),
.Y(n_2518)
);

NOR2xp67_ASAP7_75t_L g2519 ( 
.A(n_2437),
.B(n_159),
.Y(n_2519)
);

NOR2x1_ASAP7_75t_L g2520 ( 
.A(n_2437),
.B(n_160),
.Y(n_2520)
);

AOI211x1_ASAP7_75t_SL g2521 ( 
.A1(n_2456),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_2521)
);

AOI221x1_ASAP7_75t_L g2522 ( 
.A1(n_2457),
.A2(n_165),
.B1(n_161),
.B2(n_163),
.C(n_166),
.Y(n_2522)
);

OAI211xp5_ASAP7_75t_SL g2523 ( 
.A1(n_2452),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_L g2524 ( 
.A(n_2443),
.B(n_167),
.C(n_168),
.Y(n_2524)
);

NAND4xp75_ASAP7_75t_L g2525 ( 
.A(n_2438),
.B(n_170),
.C(n_168),
.D(n_169),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2472),
.B(n_169),
.Y(n_2526)
);

NAND3xp33_ASAP7_75t_L g2527 ( 
.A(n_2438),
.B(n_170),
.C(n_172),
.Y(n_2527)
);

NOR3xp33_ASAP7_75t_L g2528 ( 
.A(n_2443),
.B(n_172),
.C(n_173),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2442),
.B(n_174),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2469),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2474),
.Y(n_2531)
);

NAND3xp33_ASAP7_75t_SL g2532 ( 
.A(n_2451),
.B(n_175),
.C(n_176),
.Y(n_2532)
);

AOI211x1_ASAP7_75t_L g2533 ( 
.A1(n_2439),
.A2(n_179),
.B(n_175),
.C(n_177),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2455),
.Y(n_2534)
);

NOR3xp33_ASAP7_75t_L g2535 ( 
.A(n_2443),
.B(n_179),
.C(n_180),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2442),
.B(n_180),
.Y(n_2536)
);

AOI221xp5_ASAP7_75t_L g2537 ( 
.A1(n_2533),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.C(n_184),
.Y(n_2537)
);

NAND3xp33_ASAP7_75t_SL g2538 ( 
.A(n_2521),
.B(n_182),
.C(n_183),
.Y(n_2538)
);

AOI222xp33_ASAP7_75t_L g2539 ( 
.A1(n_2512),
.A2(n_2532),
.B1(n_2498),
.B2(n_2510),
.C1(n_2527),
.C2(n_2494),
.Y(n_2539)
);

OAI211xp5_ASAP7_75t_SL g2540 ( 
.A1(n_2488),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2540)
);

NOR2x1_ASAP7_75t_L g2541 ( 
.A(n_2487),
.B(n_185),
.Y(n_2541)
);

OAI211xp5_ASAP7_75t_L g2542 ( 
.A1(n_2477),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2542)
);

AOI221xp5_ASAP7_75t_L g2543 ( 
.A1(n_2501),
.A2(n_190),
.B1(n_188),
.B2(n_189),
.C(n_192),
.Y(n_2543)
);

OAI211xp5_ASAP7_75t_L g2544 ( 
.A1(n_2506),
.A2(n_2536),
.B(n_2529),
.C(n_2493),
.Y(n_2544)
);

AOI221xp5_ASAP7_75t_L g2545 ( 
.A1(n_2499),
.A2(n_194),
.B1(n_189),
.B2(n_190),
.C(n_195),
.Y(n_2545)
);

NAND4xp25_ASAP7_75t_L g2546 ( 
.A(n_2478),
.B(n_2476),
.C(n_2528),
.D(n_2524),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_L g2547 ( 
.A(n_2523),
.B(n_196),
.Y(n_2547)
);

AOI22xp5_ASAP7_75t_SL g2548 ( 
.A1(n_2484),
.A2(n_2073),
.B1(n_2062),
.B2(n_2175),
.Y(n_2548)
);

NOR4xp25_ASAP7_75t_L g2549 ( 
.A(n_2485),
.B(n_199),
.C(n_197),
.D(n_198),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2526),
.B(n_197),
.Y(n_2550)
);

OAI211xp5_ASAP7_75t_L g2551 ( 
.A1(n_2475),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_2551)
);

AOI221xp5_ASAP7_75t_L g2552 ( 
.A1(n_2535),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_2552)
);

AOI221xp5_ASAP7_75t_SL g2553 ( 
.A1(n_2486),
.A2(n_204),
.B1(n_201),
.B2(n_202),
.C(n_205),
.Y(n_2553)
);

OAI211xp5_ASAP7_75t_L g2554 ( 
.A1(n_2509),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_2534),
.Y(n_2555)
);

AOI221xp5_ASAP7_75t_L g2556 ( 
.A1(n_2496),
.A2(n_210),
.B1(n_206),
.B2(n_207),
.C(n_211),
.Y(n_2556)
);

NOR3xp33_ASAP7_75t_L g2557 ( 
.A(n_2508),
.B(n_210),
.C(n_211),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_L g2558 ( 
.A(n_2534),
.B(n_212),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2480),
.B(n_213),
.Y(n_2559)
);

AOI31xp33_ASAP7_75t_L g2560 ( 
.A1(n_2513),
.A2(n_215),
.A3(n_213),
.B(n_214),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2519),
.B(n_215),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2516),
.Y(n_2562)
);

XNOR2xp5_ASAP7_75t_L g2563 ( 
.A(n_2489),
.B(n_216),
.Y(n_2563)
);

OAI211xp5_ASAP7_75t_SL g2564 ( 
.A1(n_2491),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_2564)
);

OAI211xp5_ASAP7_75t_L g2565 ( 
.A1(n_2517),
.A2(n_220),
.B(n_217),
.C(n_219),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2518),
.Y(n_2566)
);

OAI211xp5_ASAP7_75t_SL g2567 ( 
.A1(n_2531),
.A2(n_224),
.B(n_221),
.C(n_223),
.Y(n_2567)
);

OAI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2497),
.A2(n_221),
.B(n_223),
.Y(n_2568)
);

AOI21xp5_ASAP7_75t_L g2569 ( 
.A1(n_2530),
.A2(n_224),
.B(n_225),
.Y(n_2569)
);

AOI211xp5_ASAP7_75t_L g2570 ( 
.A1(n_2503),
.A2(n_227),
.B(n_225),
.C(n_226),
.Y(n_2570)
);

NAND3xp33_ASAP7_75t_SL g2571 ( 
.A(n_2500),
.B(n_226),
.C(n_227),
.Y(n_2571)
);

AOI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2484),
.A2(n_2179),
.B1(n_2175),
.B2(n_2073),
.Y(n_2572)
);

AOI221xp5_ASAP7_75t_L g2573 ( 
.A1(n_2534),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.C(n_231),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2502),
.A2(n_228),
.B(n_229),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2520),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2495),
.B(n_230),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2482),
.B(n_231),
.Y(n_2577)
);

NAND3xp33_ASAP7_75t_L g2578 ( 
.A(n_2522),
.B(n_232),
.C(n_233),
.Y(n_2578)
);

O2A1O1Ixp33_ASAP7_75t_L g2579 ( 
.A1(n_2492),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_2579)
);

AO22x2_ASAP7_75t_L g2580 ( 
.A1(n_2525),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_2580)
);

O2A1O1Ixp33_ASAP7_75t_L g2581 ( 
.A1(n_2481),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_2581)
);

AOI221xp5_ASAP7_75t_SL g2582 ( 
.A1(n_2483),
.A2(n_2504),
.B1(n_2505),
.B2(n_2490),
.C(n_2514),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2479),
.B(n_238),
.Y(n_2583)
);

OR2x2_ASAP7_75t_L g2584 ( 
.A(n_2515),
.B(n_238),
.Y(n_2584)
);

OAI211xp5_ASAP7_75t_SL g2585 ( 
.A1(n_2507),
.A2(n_242),
.B(n_239),
.C(n_240),
.Y(n_2585)
);

OR2x2_ASAP7_75t_L g2586 ( 
.A(n_2507),
.B(n_239),
.Y(n_2586)
);

OAI211xp5_ASAP7_75t_SL g2587 ( 
.A1(n_2511),
.A2(n_244),
.B(n_240),
.C(n_243),
.Y(n_2587)
);

OA22x2_ASAP7_75t_L g2588 ( 
.A1(n_2512),
.A2(n_2062),
.B1(n_245),
.B2(n_243),
.Y(n_2588)
);

NAND4xp75_ASAP7_75t_L g2589 ( 
.A(n_2533),
.B(n_246),
.C(n_244),
.D(n_245),
.Y(n_2589)
);

NAND3xp33_ASAP7_75t_L g2590 ( 
.A(n_2533),
.B(n_246),
.C(n_247),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2480),
.B(n_248),
.Y(n_2591)
);

OAI221xp5_ASAP7_75t_L g2592 ( 
.A1(n_2487),
.A2(n_251),
.B1(n_248),
.B2(n_250),
.C(n_252),
.Y(n_2592)
);

OAI211xp5_ASAP7_75t_L g2593 ( 
.A1(n_2533),
.A2(n_254),
.B(n_251),
.C(n_253),
.Y(n_2593)
);

NOR3xp33_ASAP7_75t_L g2594 ( 
.A(n_2477),
.B(n_254),
.C(n_255),
.Y(n_2594)
);

AOI211xp5_ASAP7_75t_L g2595 ( 
.A1(n_2487),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2493),
.Y(n_2596)
);

AOI211xp5_ASAP7_75t_L g2597 ( 
.A1(n_2487),
.A2(n_260),
.B(n_256),
.C(n_258),
.Y(n_2597)
);

NAND3xp33_ASAP7_75t_L g2598 ( 
.A(n_2533),
.B(n_260),
.C(n_261),
.Y(n_2598)
);

AOI221x1_ASAP7_75t_L g2599 ( 
.A1(n_2487),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.C(n_264),
.Y(n_2599)
);

NAND2x1p5_ASAP7_75t_L g2600 ( 
.A(n_2493),
.B(n_2179),
.Y(n_2600)
);

AOI221xp5_ASAP7_75t_L g2601 ( 
.A1(n_2533),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.C(n_265),
.Y(n_2601)
);

NAND2xp33_ASAP7_75t_SL g2602 ( 
.A(n_2495),
.B(n_265),
.Y(n_2602)
);

OAI31xp33_ASAP7_75t_L g2603 ( 
.A1(n_2510),
.A2(n_269),
.A3(n_266),
.B(n_267),
.Y(n_2603)
);

NOR3xp33_ASAP7_75t_L g2604 ( 
.A(n_2544),
.B(n_2546),
.C(n_2596),
.Y(n_2604)
);

INVx2_ASAP7_75t_SL g2605 ( 
.A(n_2555),
.Y(n_2605)
);

NAND3xp33_ASAP7_75t_L g2606 ( 
.A(n_2545),
.B(n_267),
.C(n_270),
.Y(n_2606)
);

AND3x4_ASAP7_75t_L g2607 ( 
.A(n_2541),
.B(n_270),
.C(n_271),
.Y(n_2607)
);

CKINVDCx20_ASAP7_75t_R g2608 ( 
.A(n_2602),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2580),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2549),
.B(n_272),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2580),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2550),
.B(n_272),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2572),
.B(n_273),
.Y(n_2613)
);

BUFx6f_ASAP7_75t_L g2614 ( 
.A(n_2555),
.Y(n_2614)
);

AND3x4_ASAP7_75t_L g2615 ( 
.A(n_2576),
.B(n_273),
.C(n_274),
.Y(n_2615)
);

OAI22xp5_ASAP7_75t_SL g2616 ( 
.A1(n_2563),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2616)
);

AOI21xp33_ASAP7_75t_SL g2617 ( 
.A1(n_2560),
.A2(n_275),
.B(n_276),
.Y(n_2617)
);

AND4x1_ASAP7_75t_L g2618 ( 
.A(n_2539),
.B(n_279),
.C(n_277),
.D(n_278),
.Y(n_2618)
);

AND3x4_ASAP7_75t_L g2619 ( 
.A(n_2576),
.B(n_2557),
.C(n_2594),
.Y(n_2619)
);

AND2x4_ASAP7_75t_L g2620 ( 
.A(n_2562),
.B(n_277),
.Y(n_2620)
);

NAND3xp33_ASAP7_75t_L g2621 ( 
.A(n_2552),
.B(n_278),
.C(n_280),
.Y(n_2621)
);

AOI21xp33_ASAP7_75t_L g2622 ( 
.A1(n_2555),
.A2(n_280),
.B(n_281),
.Y(n_2622)
);

INVxp67_ASAP7_75t_L g2623 ( 
.A(n_2558),
.Y(n_2623)
);

NAND4xp75_ASAP7_75t_L g2624 ( 
.A(n_2599),
.B(n_284),
.C(n_282),
.D(n_283),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2584),
.Y(n_2625)
);

NOR2x1_ASAP7_75t_L g2626 ( 
.A(n_2566),
.B(n_282),
.Y(n_2626)
);

NOR2xp67_ASAP7_75t_L g2627 ( 
.A(n_2578),
.B(n_283),
.Y(n_2627)
);

XOR2xp5_ASAP7_75t_SL g2628 ( 
.A(n_2586),
.B(n_284),
.Y(n_2628)
);

NOR2x1_ASAP7_75t_L g2629 ( 
.A(n_2575),
.B(n_285),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2583),
.B(n_286),
.Y(n_2630)
);

OAI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_2592),
.A2(n_2072),
.B1(n_2083),
.B2(n_2067),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_2559),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2547),
.B(n_286),
.Y(n_2633)
);

OAI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2590),
.A2(n_2598),
.B(n_2593),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2595),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2588),
.Y(n_2636)
);

NOR3xp33_ASAP7_75t_L g2637 ( 
.A(n_2571),
.B(n_287),
.C(n_290),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_2561),
.Y(n_2638)
);

NOR2xp67_ASAP7_75t_L g2639 ( 
.A(n_2538),
.B(n_291),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2564),
.B(n_291),
.Y(n_2640)
);

NAND4xp75_ASAP7_75t_L g2641 ( 
.A(n_2582),
.B(n_295),
.C(n_292),
.D(n_293),
.Y(n_2641)
);

NAND2xp33_ASAP7_75t_SL g2642 ( 
.A(n_2591),
.B(n_292),
.Y(n_2642)
);

NOR3xp33_ASAP7_75t_L g2643 ( 
.A(n_2577),
.B(n_293),
.C(n_295),
.Y(n_2643)
);

NOR2x1_ASAP7_75t_L g2644 ( 
.A(n_2551),
.B(n_2554),
.Y(n_2644)
);

NOR3xp33_ASAP7_75t_L g2645 ( 
.A(n_2587),
.B(n_296),
.C(n_297),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2553),
.B(n_296),
.Y(n_2646)
);

OAI221xp5_ASAP7_75t_L g2647 ( 
.A1(n_2603),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.C(n_300),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_L g2648 ( 
.A(n_2585),
.B(n_298),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2600),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2540),
.B(n_299),
.Y(n_2650)
);

NOR3xp33_ASAP7_75t_SL g2651 ( 
.A(n_2568),
.B(n_2589),
.C(n_2565),
.Y(n_2651)
);

NAND4xp75_ASAP7_75t_L g2652 ( 
.A(n_2569),
.B(n_303),
.C(n_300),
.D(n_301),
.Y(n_2652)
);

NOR3xp33_ASAP7_75t_L g2653 ( 
.A(n_2543),
.B(n_301),
.C(n_303),
.Y(n_2653)
);

NOR2x1_ASAP7_75t_L g2654 ( 
.A(n_2542),
.B(n_304),
.Y(n_2654)
);

AOI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2567),
.A2(n_2601),
.B1(n_2537),
.B2(n_2597),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2574),
.B(n_304),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_R g2657 ( 
.A(n_2570),
.B(n_2548),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2581),
.B(n_305),
.Y(n_2658)
);

NOR3x1_ASAP7_75t_L g2659 ( 
.A(n_2579),
.B(n_2556),
.C(n_2573),
.Y(n_2659)
);

NOR2x1_ASAP7_75t_L g2660 ( 
.A(n_2596),
.B(n_305),
.Y(n_2660)
);

NOR2x1_ASAP7_75t_L g2661 ( 
.A(n_2596),
.B(n_306),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2580),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2550),
.B(n_306),
.Y(n_2663)
);

NOR5xp2_ASAP7_75t_L g2664 ( 
.A(n_2544),
.B(n_307),
.C(n_309),
.D(n_310),
.E(n_311),
.Y(n_2664)
);

AOI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2602),
.A2(n_310),
.B1(n_307),
.B2(n_309),
.Y(n_2665)
);

AOI22xp5_ASAP7_75t_L g2666 ( 
.A1(n_2602),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_2666)
);

AOI211xp5_ASAP7_75t_L g2667 ( 
.A1(n_2587),
.A2(n_317),
.B(n_313),
.C(n_314),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2580),
.Y(n_2668)
);

OAI211xp5_ASAP7_75t_L g2669 ( 
.A1(n_2665),
.A2(n_2666),
.B(n_2617),
.C(n_2634),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2620),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2663),
.B(n_314),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2614),
.B(n_318),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2628),
.B(n_318),
.Y(n_2673)
);

OAI222xp33_ASAP7_75t_L g2674 ( 
.A1(n_2610),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.C1(n_322),
.C2(n_323),
.Y(n_2674)
);

XNOR2xp5_ASAP7_75t_L g2675 ( 
.A(n_2615),
.B(n_319),
.Y(n_2675)
);

AOI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2608),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_SL g2677 ( 
.A1(n_2605),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_2677)
);

NOR3xp33_ASAP7_75t_SL g2678 ( 
.A(n_2642),
.B(n_326),
.C(n_327),
.Y(n_2678)
);

NAND3xp33_ASAP7_75t_L g2679 ( 
.A(n_2643),
.B(n_327),
.C(n_328),
.Y(n_2679)
);

XNOR2xp5_ASAP7_75t_L g2680 ( 
.A(n_2607),
.B(n_329),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2626),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2614),
.B(n_329),
.Y(n_2682)
);

NAND3xp33_ASAP7_75t_SL g2683 ( 
.A(n_2604),
.B(n_330),
.C(n_331),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_2646),
.A2(n_2656),
.B(n_2639),
.Y(n_2684)
);

NOR3xp33_ASAP7_75t_L g2685 ( 
.A(n_2625),
.B(n_330),
.C(n_333),
.Y(n_2685)
);

NAND4xp25_ASAP7_75t_SL g2686 ( 
.A(n_2667),
.B(n_336),
.C(n_334),
.D(n_335),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2655),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2687)
);

NAND5xp2_ASAP7_75t_L g2688 ( 
.A(n_2651),
.B(n_337),
.C(n_338),
.D(n_339),
.E(n_340),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_SL g2689 ( 
.A1(n_2648),
.A2(n_341),
.B1(n_338),
.B2(n_339),
.Y(n_2689)
);

NOR3xp33_ASAP7_75t_L g2690 ( 
.A(n_2649),
.B(n_341),
.C(n_342),
.Y(n_2690)
);

OR2x2_ASAP7_75t_L g2691 ( 
.A(n_2630),
.B(n_342),
.Y(n_2691)
);

NOR3xp33_ASAP7_75t_L g2692 ( 
.A(n_2616),
.B(n_343),
.C(n_344),
.Y(n_2692)
);

XOR2x2_ASAP7_75t_L g2693 ( 
.A(n_2624),
.B(n_2652),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2633),
.B(n_2645),
.Y(n_2694)
);

AO22x2_ASAP7_75t_L g2695 ( 
.A1(n_2609),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_2695)
);

NAND4xp75_ASAP7_75t_L g2696 ( 
.A(n_2629),
.B(n_348),
.C(n_346),
.D(n_347),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2612),
.B(n_347),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2618),
.B(n_348),
.Y(n_2698)
);

OAI211xp5_ASAP7_75t_L g2699 ( 
.A1(n_2660),
.A2(n_351),
.B(n_349),
.C(n_350),
.Y(n_2699)
);

OAI322xp33_ASAP7_75t_L g2700 ( 
.A1(n_2611),
.A2(n_349),
.A3(n_350),
.B1(n_352),
.B2(n_353),
.C1(n_354),
.C2(n_355),
.Y(n_2700)
);

NAND3xp33_ASAP7_75t_L g2701 ( 
.A(n_2637),
.B(n_352),
.C(n_353),
.Y(n_2701)
);

OAI221xp5_ASAP7_75t_L g2702 ( 
.A1(n_2647),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.C(n_357),
.Y(n_2702)
);

O2A1O1Ixp33_ASAP7_75t_L g2703 ( 
.A1(n_2662),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_2703)
);

NAND3xp33_ASAP7_75t_SL g2704 ( 
.A(n_2664),
.B(n_358),
.C(n_359),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2661),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_SL g2706 ( 
.A1(n_2650),
.A2(n_2640),
.B1(n_2614),
.B2(n_2636),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_2668),
.Y(n_2707)
);

AOI211xp5_ASAP7_75t_L g2708 ( 
.A1(n_2635),
.A2(n_359),
.B(n_361),
.C(n_362),
.Y(n_2708)
);

AND4x1_ASAP7_75t_L g2709 ( 
.A(n_2644),
.B(n_362),
.C(n_363),
.D(n_364),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2641),
.Y(n_2710)
);

NOR3x1_ASAP7_75t_SL g2711 ( 
.A(n_2632),
.B(n_364),
.C(n_365),
.Y(n_2711)
);

NOR4xp25_ASAP7_75t_L g2712 ( 
.A(n_2623),
.B(n_2606),
.C(n_2621),
.D(n_2622),
.Y(n_2712)
);

NAND4xp25_ASAP7_75t_L g2713 ( 
.A(n_2659),
.B(n_365),
.C(n_366),
.D(n_367),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2711),
.Y(n_2714)
);

OAI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2689),
.A2(n_2627),
.B1(n_2619),
.B2(n_2654),
.Y(n_2715)
);

XOR2xp5_ASAP7_75t_L g2716 ( 
.A(n_2680),
.B(n_2638),
.Y(n_2716)
);

INVx2_ASAP7_75t_SL g2717 ( 
.A(n_2673),
.Y(n_2717)
);

OAI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2701),
.A2(n_2658),
.B1(n_2613),
.B2(n_2653),
.Y(n_2718)
);

BUFx10_ASAP7_75t_L g2719 ( 
.A(n_2681),
.Y(n_2719)
);

AOI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2686),
.A2(n_2658),
.B1(n_2620),
.B2(n_2631),
.Y(n_2720)
);

NAND3x1_ASAP7_75t_L g2721 ( 
.A(n_2692),
.B(n_2657),
.C(n_367),
.Y(n_2721)
);

AOI221xp5_ASAP7_75t_SL g2722 ( 
.A1(n_2684),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.C(n_371),
.Y(n_2722)
);

AOI22x1_ASAP7_75t_L g2723 ( 
.A1(n_2675),
.A2(n_368),
.B1(n_370),
.B2(n_371),
.Y(n_2723)
);

OAI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2698),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_2724)
);

OAI22xp5_ASAP7_75t_L g2725 ( 
.A1(n_2671),
.A2(n_2679),
.B1(n_2710),
.B2(n_2702),
.Y(n_2725)
);

AND3x2_ASAP7_75t_L g2726 ( 
.A(n_2707),
.B(n_372),
.C(n_374),
.Y(n_2726)
);

INVxp67_ASAP7_75t_L g2727 ( 
.A(n_2688),
.Y(n_2727)
);

NOR3xp33_ASAP7_75t_SL g2728 ( 
.A(n_2683),
.B(n_375),
.C(n_376),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2697),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2685),
.B(n_375),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2696),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_2705),
.B(n_376),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2690),
.B(n_377),
.Y(n_2733)
);

AOI221xp5_ASAP7_75t_L g2734 ( 
.A1(n_2704),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.C(n_381),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_SL g2735 ( 
.A(n_2674),
.B(n_378),
.Y(n_2735)
);

INVxp67_ASAP7_75t_SL g2736 ( 
.A(n_2672),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2709),
.B(n_379),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2706),
.A2(n_380),
.B1(n_381),
.B2(n_382),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2691),
.Y(n_2739)
);

XNOR2x1_ASAP7_75t_L g2740 ( 
.A(n_2693),
.B(n_383),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2682),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2695),
.Y(n_2742)
);

OR3x2_ASAP7_75t_L g2743 ( 
.A(n_2713),
.B(n_2678),
.C(n_2712),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_SL g2744 ( 
.A(n_2708),
.B(n_383),
.Y(n_2744)
);

AOI211xp5_ASAP7_75t_L g2745 ( 
.A1(n_2699),
.A2(n_384),
.B(n_386),
.C(n_387),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2670),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2695),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2694),
.Y(n_2748)
);

AND2x4_ASAP7_75t_L g2749 ( 
.A(n_2676),
.B(n_387),
.Y(n_2749)
);

NOR3x1_ASAP7_75t_L g2750 ( 
.A(n_2737),
.B(n_2669),
.C(n_2687),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2742),
.Y(n_2751)
);

AOI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2746),
.A2(n_2677),
.B1(n_2703),
.B2(n_2700),
.Y(n_2752)
);

AOI22xp5_ASAP7_75t_L g2753 ( 
.A1(n_2740),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_2753)
);

OAI22xp5_ASAP7_75t_SL g2754 ( 
.A1(n_2714),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_2754)
);

OA22x2_ASAP7_75t_L g2755 ( 
.A1(n_2720),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_2755)
);

OAI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_2727),
.A2(n_391),
.B1(n_392),
.B2(n_394),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2726),
.Y(n_2757)
);

NOR4xp25_ASAP7_75t_L g2758 ( 
.A(n_2721),
.B(n_394),
.C(n_395),
.D(n_396),
.Y(n_2758)
);

HB1xp67_ASAP7_75t_L g2759 ( 
.A(n_2747),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2728),
.B(n_397),
.Y(n_2760)
);

INVx3_ASAP7_75t_SL g2761 ( 
.A(n_2719),
.Y(n_2761)
);

OAI22x1_ASAP7_75t_L g2762 ( 
.A1(n_2723),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.Y(n_2762)
);

OR4x2_ASAP7_75t_L g2763 ( 
.A(n_2743),
.B(n_398),
.C(n_400),
.D(n_401),
.Y(n_2763)
);

OAI22x1_ASAP7_75t_L g2764 ( 
.A1(n_2731),
.A2(n_400),
.B1(n_402),
.B2(n_403),
.Y(n_2764)
);

AO22x2_ASAP7_75t_L g2765 ( 
.A1(n_2715),
.A2(n_404),
.B1(n_405),
.B2(n_407),
.Y(n_2765)
);

NOR3xp33_ASAP7_75t_SL g2766 ( 
.A(n_2725),
.B(n_405),
.C(n_408),
.Y(n_2766)
);

OAI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2745),
.A2(n_408),
.B1(n_409),
.B2(n_410),
.Y(n_2767)
);

AOI221xp5_ASAP7_75t_L g2768 ( 
.A1(n_2734),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.C(n_412),
.Y(n_2768)
);

OR4x2_ASAP7_75t_L g2769 ( 
.A(n_2735),
.B(n_411),
.C(n_412),
.D(n_413),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2724),
.Y(n_2770)
);

XOR2xp5_ASAP7_75t_L g2771 ( 
.A(n_2716),
.B(n_413),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2732),
.Y(n_2772)
);

NOR2xp33_ASAP7_75t_L g2773 ( 
.A(n_2733),
.B(n_414),
.Y(n_2773)
);

OR4x1_ASAP7_75t_L g2774 ( 
.A(n_2717),
.B(n_414),
.C(n_415),
.D(n_416),
.Y(n_2774)
);

NOR3xp33_ASAP7_75t_L g2775 ( 
.A(n_2748),
.B(n_415),
.C(n_416),
.Y(n_2775)
);

HB1xp67_ASAP7_75t_L g2776 ( 
.A(n_2738),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2769),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2751),
.A2(n_2730),
.B1(n_2736),
.B2(n_2741),
.Y(n_2778)
);

XNOR2xp5_ASAP7_75t_L g2779 ( 
.A(n_2762),
.B(n_2718),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2774),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2765),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2755),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2758),
.B(n_2722),
.Y(n_2783)
);

OAI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2761),
.A2(n_2749),
.B1(n_2739),
.B2(n_2729),
.Y(n_2784)
);

AOI22xp5_ASAP7_75t_SL g2785 ( 
.A1(n_2757),
.A2(n_2732),
.B1(n_2744),
.B2(n_420),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2771),
.Y(n_2786)
);

INVx2_ASAP7_75t_SL g2787 ( 
.A(n_2763),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2765),
.Y(n_2788)
);

INVx3_ASAP7_75t_L g2789 ( 
.A(n_2772),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_SL g2790 ( 
.A1(n_2773),
.A2(n_417),
.B1(n_418),
.B2(n_420),
.Y(n_2790)
);

AOI21xp33_ASAP7_75t_SL g2791 ( 
.A1(n_2767),
.A2(n_417),
.B(n_418),
.Y(n_2791)
);

OA21x2_ASAP7_75t_L g2792 ( 
.A1(n_2752),
.A2(n_421),
.B(n_422),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2760),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2764),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_L g2795 ( 
.A1(n_2759),
.A2(n_425),
.B1(n_426),
.B2(n_428),
.Y(n_2795)
);

OAI22xp5_ASAP7_75t_SL g2796 ( 
.A1(n_2776),
.A2(n_426),
.B1(n_428),
.B2(n_429),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2793),
.B(n_2766),
.Y(n_2797)
);

O2A1O1Ixp33_ASAP7_75t_L g2798 ( 
.A1(n_2781),
.A2(n_2770),
.B(n_2768),
.C(n_2775),
.Y(n_2798)
);

O2A1O1Ixp33_ASAP7_75t_L g2799 ( 
.A1(n_2788),
.A2(n_2756),
.B(n_2750),
.C(n_2753),
.Y(n_2799)
);

AND3x4_ASAP7_75t_L g2800 ( 
.A(n_2780),
.B(n_2754),
.C(n_430),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2792),
.Y(n_2801)
);

AOI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2783),
.A2(n_429),
.B(n_430),
.Y(n_2802)
);

AO22x2_ASAP7_75t_L g2803 ( 
.A1(n_2787),
.A2(n_2777),
.B1(n_2784),
.B2(n_2782),
.Y(n_2803)
);

AND3x4_ASAP7_75t_L g2804 ( 
.A(n_2794),
.B(n_2779),
.C(n_2785),
.Y(n_2804)
);

OA22x2_ASAP7_75t_L g2805 ( 
.A1(n_2789),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_2805)
);

AND3x4_ASAP7_75t_L g2806 ( 
.A(n_2791),
.B(n_431),
.C(n_432),
.Y(n_2806)
);

OAI222xp33_ASAP7_75t_L g2807 ( 
.A1(n_2778),
.A2(n_434),
.B1(n_435),
.B2(n_436),
.C1(n_438),
.C2(n_439),
.Y(n_2807)
);

XNOR2xp5_ASAP7_75t_L g2808 ( 
.A(n_2786),
.B(n_434),
.Y(n_2808)
);

NAND3xp33_ASAP7_75t_SL g2809 ( 
.A(n_2795),
.B(n_435),
.C(n_436),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_SL g2810 ( 
.A1(n_2800),
.A2(n_2790),
.B1(n_2796),
.B2(n_440),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2806),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2805),
.Y(n_2812)
);

OAI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2804),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_2813)
);

AO22x2_ASAP7_75t_L g2814 ( 
.A1(n_2801),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2808),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2799),
.A2(n_444),
.B(n_445),
.Y(n_2816)
);

AOI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2803),
.A2(n_2809),
.B1(n_2797),
.B2(n_2802),
.Y(n_2817)
);

HB1xp67_ASAP7_75t_L g2818 ( 
.A(n_2807),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2814),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2813),
.Y(n_2820)
);

OAI22xp33_ASAP7_75t_L g2821 ( 
.A1(n_2817),
.A2(n_2798),
.B1(n_445),
.B2(n_446),
.Y(n_2821)
);

NOR2x1p5_ASAP7_75t_L g2822 ( 
.A(n_2812),
.B(n_444),
.Y(n_2822)
);

AOI22xp5_ASAP7_75t_L g2823 ( 
.A1(n_2811),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_2823)
);

INVx4_ASAP7_75t_L g2824 ( 
.A(n_2815),
.Y(n_2824)
);

AOI21xp33_ASAP7_75t_SL g2825 ( 
.A1(n_2821),
.A2(n_2810),
.B(n_2818),
.Y(n_2825)
);

OAI211xp5_ASAP7_75t_L g2826 ( 
.A1(n_2823),
.A2(n_2816),
.B(n_449),
.C(n_450),
.Y(n_2826)
);

OAI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2820),
.A2(n_448),
.B(n_450),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2822),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2828),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2826),
.Y(n_2830)
);

XOR2xp5_ASAP7_75t_L g2831 ( 
.A(n_2827),
.B(n_2819),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_L g2832 ( 
.A1(n_2829),
.A2(n_2824),
.B1(n_2825),
.B2(n_453),
.Y(n_2832)
);

XNOR2xp5_ASAP7_75t_L g2833 ( 
.A(n_2831),
.B(n_451),
.Y(n_2833)
);

AOI31xp33_ASAP7_75t_L g2834 ( 
.A1(n_2830),
.A2(n_451),
.A3(n_452),
.B(n_454),
.Y(n_2834)
);

NAND2x1p5_ASAP7_75t_L g2835 ( 
.A(n_2830),
.B(n_455),
.Y(n_2835)
);

AND2x2_ASAP7_75t_SL g2836 ( 
.A(n_2832),
.B(n_455),
.Y(n_2836)
);

OAI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2835),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.Y(n_2837)
);

OR2x6_ASAP7_75t_L g2838 ( 
.A(n_2836),
.B(n_2833),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2838),
.A2(n_2837),
.B(n_2834),
.Y(n_2839)
);

AOI211xp5_ASAP7_75t_L g2840 ( 
.A1(n_2839),
.A2(n_456),
.B(n_458),
.C(n_459),
.Y(n_2840)
);


endmodule