module fake_netlist_6_288_n_2001 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2001);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2001;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_22),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_148),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_107),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_40),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_13),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_92),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_84),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_59),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_69),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_75),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_162),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_76),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_77),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_104),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_14),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_1),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_53),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_167),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_74),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_115),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_62),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_81),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_139),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_34),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_108),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_47),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_159),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_71),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_21),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_143),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_196),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_70),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_138),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_178),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_102),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_63),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_52),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_132),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_110),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_49),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_136),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_160),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_175),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_37),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_154),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_172),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_25),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_103),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_93),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_64),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_37),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_6),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_61),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_98),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_52),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_141),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_168),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_89),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_124),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_181),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_10),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_188),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_9),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_8),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_60),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_30),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_1),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_161),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_146),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_7),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_180),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_70),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_125),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_86),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_184),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_131),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_134),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_119),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_35),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_156),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_25),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_193),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_16),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_129),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_165),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_96),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_22),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_2),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_197),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_142),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_40),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_57),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_36),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_31),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_16),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_80),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_27),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_97),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_19),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_44),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_5),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_83),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_62),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_170),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_112),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_65),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_28),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_152),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_61),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_192),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_117),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_150),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_87),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_128),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_105),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_109),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_72),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_85),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_42),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_13),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_123),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_130),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_27),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_179),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_19),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_65),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_6),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_35),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_38),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_42),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_29),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_99),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_43),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_30),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_71),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_33),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_95),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_201),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_100),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_94),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_163),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_33),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_41),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_147),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_20),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_111),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_91),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_12),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_200),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_28),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_66),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_49),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_153),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_45),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_82),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_36),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_2),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_5),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_51),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_145),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_12),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_8),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_58),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_57),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_4),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_51),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_4),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_54),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_122),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_79),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_169),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_54),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_187),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_88),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_34),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_41),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_53),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_39),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_120),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_219),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_228),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_215),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_353),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_253),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_222),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_353),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_353),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_353),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_209),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_232),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_209),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_271),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_258),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_271),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_305),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_233),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_305),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_247),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_239),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_381),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_262),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_247),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_265),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_357),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_249),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_204),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_280),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_214),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_215),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_315),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_266),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_269),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_348),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_298),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_270),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_276),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_250),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_225),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_321),
.Y(n_453)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_217),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_279),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_280),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_227),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_281),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_229),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_230),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_284),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_244),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_255),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_327),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_291),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_259),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_345),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_217),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_264),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_274),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_283),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_293),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_246),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_287),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_310),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_297),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_236),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_290),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_302),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_236),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_304),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_306),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_392),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_311),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_300),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_246),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_318),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_322),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_241),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_308),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_323),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_342),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_346),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_309),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_365),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_368),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_290),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_313),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_319),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_278),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_278),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_371),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_325),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_380),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_382),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_386),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_404),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_431),
.A2(n_251),
.B1(n_401),
.B2(n_400),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_413),
.B(n_216),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_422),
.B(n_216),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_278),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_254),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_485),
.B(n_446),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_438),
.B(n_242),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_501),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_404),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_501),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_500),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_500),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_405),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_480),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_456),
.B(n_242),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_405),
.B(n_278),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_407),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_407),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_406),
.A2(n_326),
.B1(n_288),
.B2(n_387),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_408),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_432),
.B(n_254),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_403),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_434),
.B(n_257),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_409),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_411),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_411),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_412),
.B(n_205),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_480),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_412),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_415),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_415),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_416),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_416),
.B(n_207),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_417),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_426),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_419),
.A2(n_251),
.B1(n_401),
.B2(n_400),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_437),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

NAND2x1p5_ASAP7_75t_L g553 ( 
.A(n_452),
.B(n_328),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_486),
.B(n_237),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_441),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_418),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_444),
.B(n_263),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_439),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_466),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_457),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_478),
.B(n_208),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_487),
.B(n_388),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_418),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_448),
.B(n_211),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_420),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_449),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_459),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_450),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_420),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_421),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_455),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_421),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_458),
.B(n_202),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_459),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_473),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_423),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_461),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_423),
.B(n_278),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_465),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_472),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_460),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_410),
.A2(n_354),
.B1(n_330),
.B2(n_398),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_497),
.B(n_237),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_476),
.B(n_212),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_424),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_424),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_R g592 ( 
.A(n_555),
.B(n_440),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_510),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_571),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_508),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_535),
.B(n_479),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_553),
.A2(n_587),
.B1(n_566),
.B2(n_512),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_L g598 ( 
.A(n_509),
.B(n_489),
.C(n_351),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_508),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_511),
.B(n_481),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_519),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_555),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_563),
.B(n_482),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_578),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_553),
.B(n_490),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_533),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_532),
.B(n_494),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_553),
.B(n_443),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_533),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_563),
.B(n_498),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_563),
.B(n_503),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_563),
.B(n_213),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_537),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_562),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_576),
.B(n_454),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_534),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_519),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_568),
.B(n_468),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_557),
.B(n_477),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_523),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_586),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_537),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_538),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_582),
.B(n_499),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_539),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_523),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_538),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_544),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_583),
.B(n_489),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_513),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_527),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_544),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_547),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_547),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_574),
.B(n_505),
.Y(n_635)
);

AND3x2_ASAP7_75t_L g636 ( 
.A(n_578),
.B(n_240),
.C(n_223),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_540),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_530),
.Y(n_639)
);

INVx6_ASAP7_75t_L g640 ( 
.A(n_539),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_580),
.B(n_445),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_530),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_586),
.B(n_451),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_524),
.B(n_237),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_531),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_SL g647 ( 
.A(n_524),
.B(n_241),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_539),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_530),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_585),
.B(n_202),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_539),
.Y(n_651)
);

BUFx4f_ASAP7_75t_L g652 ( 
.A(n_545),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_564),
.B(n_429),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_572),
.Y(n_654)
);

BUFx4f_ASAP7_75t_L g655 ( 
.A(n_545),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_572),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_572),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_517),
.B(n_429),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_572),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

AO21x2_ASAP7_75t_L g661 ( 
.A1(n_545),
.A2(n_260),
.B(n_243),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_585),
.A2(n_273),
.B1(n_256),
.B2(n_261),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_554),
.A2(n_516),
.B1(n_525),
.B2(n_550),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

INVx4_ASAP7_75t_SL g665 ( 
.A(n_513),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_536),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_545),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_564),
.B(n_433),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_510),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_540),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_536),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_515),
.B(n_282),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_572),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_510),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_564),
.B(n_433),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_510),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_570),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_572),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_540),
.B(n_203),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_510),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_564),
.B(n_435),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_564),
.B(n_435),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_510),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_577),
.B(n_414),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_584),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_518),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_540),
.A2(n_453),
.B1(n_425),
.B2(n_483),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_529),
.B(n_203),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_515),
.Y(n_689)
);

AO22x2_ASAP7_75t_L g690 ( 
.A1(n_529),
.A2(n_399),
.B1(n_356),
.B2(n_210),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_584),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_521),
.B(n_295),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_541),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_521),
.B(n_296),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_541),
.Y(n_695)
);

BUFx8_ASAP7_75t_SL g696 ( 
.A(n_589),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_546),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_589),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_521),
.B(n_299),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_590),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_590),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_527),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_521),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_518),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_522),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_551),
.Y(n_707)
);

CKINVDCx6p67_ASAP7_75t_R g708 ( 
.A(n_581),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_527),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_527),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_527),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_522),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_552),
.A2(n_294),
.B1(n_292),
.B2(n_289),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_522),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_552),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_522),
.B(n_307),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_548),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_520),
.B(n_312),
.Y(n_718)
);

XOR2xp5_ASAP7_75t_SL g719 ( 
.A(n_558),
.B(n_336),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_520),
.B(n_337),
.Y(n_720)
);

BUFx6f_ASAP7_75t_SL g721 ( 
.A(n_558),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_565),
.B(n_427),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_565),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_549),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_528),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_559),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_549),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_528),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_556),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_528),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_619),
.B(n_430),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_614),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_621),
.A2(n_464),
.B1(n_436),
.B2(n_442),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_693),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_625),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_689),
.B(n_556),
.Y(n_736)
);

NAND2x1p5_ASAP7_75t_L g737 ( 
.A(n_625),
.B(n_361),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_693),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_621),
.A2(n_447),
.B1(n_467),
.B2(n_364),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_689),
.B(n_600),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_597),
.B(n_335),
.Y(n_741)
);

O2A1O1Ixp5_ASAP7_75t_L g742 ( 
.A1(n_612),
.A2(n_397),
.B(n_393),
.C(n_362),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_652),
.B(n_335),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_635),
.B(n_206),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_695),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_594),
.B(n_246),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_607),
.B(n_698),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_706),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_695),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_658),
.A2(n_384),
.B(n_366),
.C(n_488),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_604),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_604),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_698),
.B(n_556),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_723),
.B(n_556),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_596),
.B(n_603),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_697),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_652),
.B(n_335),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_653),
.B(n_369),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_700),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_700),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_610),
.B(n_218),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_701),
.B(n_268),
.C(n_267),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_637),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_707),
.B(n_462),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_723),
.B(n_567),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_643),
.B(n_567),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_717),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_660),
.B(n_567),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_611),
.B(n_218),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_661),
.A2(n_383),
.B1(n_402),
.B2(n_376),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_602),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_652),
.B(n_335),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_SL g773 ( 
.A1(n_687),
.A2(n_358),
.B1(n_330),
.B2(n_340),
.Y(n_773)
);

BUFx6f_ASAP7_75t_SL g774 ( 
.A(n_608),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_677),
.B(n_567),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_717),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_624),
.B(n_573),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_655),
.B(n_648),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_615),
.B(n_220),
.Y(n_779)
);

INVx8_ASAP7_75t_L g780 ( 
.A(n_653),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_724),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_685),
.B(n_573),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_691),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_655),
.B(n_347),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_702),
.B(n_726),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_704),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_595),
.B(n_573),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_595),
.B(n_588),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_724),
.Y(n_789)
);

NOR3xp33_ASAP7_75t_L g790 ( 
.A(n_629),
.B(n_469),
.C(n_463),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_599),
.B(n_588),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_602),
.Y(n_792)
);

BUFx6f_ASAP7_75t_SL g793 ( 
.A(n_608),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_599),
.B(n_588),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_601),
.B(n_588),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_601),
.B(n_528),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_592),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_712),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_655),
.B(n_347),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_617),
.B(n_528),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_648),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_701),
.B(n_347),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_641),
.B(n_275),
.C(n_272),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_684),
.B(n_463),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_617),
.B(n_542),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_661),
.A2(n_372),
.B1(n_370),
.B2(n_347),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_638),
.B(n_559),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_620),
.B(n_542),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_668),
.B(n_469),
.Y(n_809)
);

NOR2xp67_ASAP7_75t_L g810 ( 
.A(n_638),
.B(n_560),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_620),
.B(n_542),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_729),
.B(n_347),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_672),
.A2(n_495),
.B(n_470),
.C(n_471),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_729),
.B(n_714),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_647),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_651),
.B(n_220),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_626),
.B(n_542),
.Y(n_817)
);

INVxp33_ASAP7_75t_SL g818 ( 
.A(n_616),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_712),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_598),
.B(n_470),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_651),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_667),
.B(n_221),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_667),
.B(n_221),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_646),
.B(n_542),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_646),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_664),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_727),
.Y(n_827)
);

CKINVDCx14_ASAP7_75t_R g828 ( 
.A(n_670),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_727),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_668),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_663),
.B(n_224),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_715),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_653),
.B(n_560),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_543),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_715),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_636),
.Y(n_836)
);

NAND2xp33_ASAP7_75t_L g837 ( 
.A(n_714),
.B(n_513),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_666),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_653),
.B(n_561),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_666),
.B(n_543),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_706),
.B(n_224),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_644),
.B(n_226),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_671),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_630),
.B(n_513),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_640),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_671),
.B(n_543),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_608),
.A2(n_358),
.B1(n_373),
.B2(n_377),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_650),
.B(n_226),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_618),
.B(n_471),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_630),
.B(n_231),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_630),
.B(n_231),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_L g852 ( 
.A(n_630),
.B(n_513),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_630),
.B(n_234),
.Y(n_853)
);

AO22x2_ASAP7_75t_L g854 ( 
.A1(n_688),
.A2(n_493),
.B1(n_474),
.B2(n_475),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_640),
.B(n_543),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_593),
.B(n_575),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_593),
.B(n_575),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_606),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_605),
.B(n_234),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_662),
.B(n_235),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_654),
.B(n_235),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_722),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_647),
.B(n_238),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_606),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_722),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_679),
.B(n_238),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_593),
.B(n_575),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_675),
.B(n_245),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_609),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_675),
.A2(n_245),
.B1(n_248),
.B2(n_252),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_654),
.B(n_248),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_661),
.A2(n_690),
.B1(n_681),
.B2(n_682),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_676),
.B(n_579),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_L g874 ( 
.A(n_713),
.B(n_561),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_609),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_616),
.B(n_252),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_676),
.B(n_579),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_675),
.B(n_331),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_613),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_665),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_613),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_665),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_680),
.B(n_591),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_690),
.A2(n_581),
.B1(n_526),
.B2(n_591),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_656),
.B(n_331),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_675),
.B(n_333),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_670),
.B(n_475),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_845),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_740),
.B(n_681),
.Y(n_889)
);

AND2x4_ASAP7_75t_SL g890 ( 
.A(n_792),
.B(n_681),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_735),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_767),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_831),
.A2(n_690),
.B1(n_681),
.B2(n_682),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_L g894 ( 
.A1(n_744),
.A2(n_779),
.B(n_804),
.Y(n_894)
);

O2A1O1Ixp5_ASAP7_75t_L g895 ( 
.A1(n_741),
.A2(n_699),
.B(n_694),
.C(n_692),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_747),
.B(n_682),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_845),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_767),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_776),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_780),
.B(n_682),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_818),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_797),
.B(n_721),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_755),
.B(n_721),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_831),
.A2(n_690),
.B1(n_622),
.B2(n_623),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_776),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_781),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_880),
.B(n_631),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_771),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_781),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_764),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_789),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_785),
.B(n_721),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_746),
.B(n_484),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_766),
.B(n_680),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_789),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_777),
.B(n_665),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_880),
.Y(n_917)
);

AOI22xp33_ASAP7_75t_L g918 ( 
.A1(n_860),
.A2(n_634),
.B1(n_622),
.B2(n_623),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_735),
.A2(n_708),
.B1(n_716),
.B2(n_720),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_825),
.B(n_686),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_827),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_748),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_801),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_848),
.A2(n_491),
.B(n_492),
.C(n_493),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_826),
.B(n_686),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_827),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_780),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_828),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_815),
.B(n_696),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_863),
.B(n_859),
.C(n_769),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_829),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_829),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_843),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_843),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_786),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_849),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_787),
.A2(n_718),
.B(n_659),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_838),
.B(n_686),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_761),
.B(n_705),
.Y(n_939)
);

NOR2x1p5_ASAP7_75t_L g940 ( 
.A(n_762),
.B(n_340),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_862),
.B(n_705),
.Y(n_941)
);

NOR2x2_ASAP7_75t_L g942 ( 
.A(n_758),
.B(n_696),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_748),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_865),
.B(n_705),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_882),
.B(n_657),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_887),
.B(n_484),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_809),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_798),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_866),
.A2(n_750),
.B(n_842),
.C(n_820),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_732),
.B(n_627),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_819),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_748),
.Y(n_952)
);

OAI21xp33_ASAP7_75t_L g953 ( 
.A1(n_750),
.A2(n_349),
.B(n_343),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_734),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_801),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_738),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_751),
.B(n_725),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_821),
.A2(n_678),
.B1(n_673),
.B2(n_659),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_833),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_858),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_872),
.B(n_673),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_818),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_855),
.A2(n_645),
.B(n_669),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_SL g964 ( 
.A(n_835),
.B(n_349),
.C(n_343),
.Y(n_964)
);

AND2x6_ASAP7_75t_L g965 ( 
.A(n_833),
.B(n_678),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_745),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_780),
.B(n_491),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_763),
.B(n_628),
.Y(n_968)
);

NOR2x2_ASAP7_75t_L g969 ( 
.A(n_758),
.B(n_719),
.Y(n_969)
);

NOR2x1p5_ASAP7_75t_L g970 ( 
.A(n_803),
.B(n_350),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_752),
.B(n_277),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_745),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_780),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_SL g974 ( 
.A1(n_731),
.A2(n_373),
.B1(n_350),
.B2(n_354),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_864),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_749),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_832),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_833),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_783),
.B(n_632),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_839),
.B(n_492),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_756),
.B(n_633),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_756),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_830),
.B(n_495),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_839),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_759),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_759),
.B(n_633),
.Y(n_986)
);

BUFx2_ASAP7_75t_L g987 ( 
.A(n_876),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_839),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_760),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_875),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_760),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_874),
.B(n_634),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_737),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_758),
.Y(n_994)
);

OAI21xp33_ASAP7_75t_SL g995 ( 
.A1(n_778),
.A2(n_496),
.B(n_506),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_869),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_790),
.B(n_496),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_875),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_753),
.B(n_703),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_778),
.B(n_709),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_879),
.Y(n_1001)
);

BUFx8_ASAP7_75t_L g1002 ( 
.A(n_774),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_774),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_736),
.A2(n_674),
.B(n_669),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_881),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_881),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_788),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_739),
.B(n_285),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_791),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_758),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_854),
.B(n_709),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_856),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_854),
.B(n_754),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_807),
.B(n_810),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_794),
.B(n_710),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_L g1016 ( 
.A(n_733),
.B(n_367),
.C(n_378),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_814),
.A2(n_674),
.B(n_669),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_857),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_854),
.B(n_710),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_802),
.A2(n_730),
.B1(n_728),
.B2(n_711),
.Y(n_1020)
);

NAND2x2_ASAP7_75t_L g1021 ( 
.A(n_836),
.B(n_359),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_765),
.B(n_711),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_795),
.B(n_728),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_847),
.B(n_816),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_R g1025 ( 
.A(n_828),
.B(n_708),
.Y(n_1025)
);

CKINVDCx14_ASAP7_75t_R g1026 ( 
.A(n_773),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_SL g1027 ( 
.A1(n_774),
.A2(n_385),
.B1(n_395),
.B2(n_398),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_L g1028 ( 
.A(n_770),
.B(n_669),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_768),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_867),
.Y(n_1030)
);

AOI21xp33_ASAP7_75t_L g1031 ( 
.A1(n_868),
.A2(n_301),
.B(n_329),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_793),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_806),
.A2(n_642),
.B1(n_639),
.B2(n_649),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_775),
.B(n_639),
.Y(n_1034)
);

NOR2xp67_ASAP7_75t_L g1035 ( 
.A(n_870),
.B(n_878),
.Y(n_1035)
);

INVxp67_ASAP7_75t_L g1036 ( 
.A(n_816),
.Y(n_1036)
);

BUFx8_ASAP7_75t_SL g1037 ( 
.A(n_793),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_782),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_796),
.Y(n_1039)
);

BUFx4f_ASAP7_75t_L g1040 ( 
.A(n_793),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_886),
.B(n_649),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_800),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_805),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_808),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_811),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_873),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_877),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_822),
.A2(n_367),
.B1(n_344),
.B2(n_341),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_822),
.A2(n_378),
.B1(n_341),
.B2(n_394),
.Y(n_1049)
);

AND2x4_ASAP7_75t_SL g1050 ( 
.A(n_884),
.B(n_683),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_817),
.Y(n_1051)
);

BUFx8_ASAP7_75t_SL g1052 ( 
.A(n_824),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_834),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_823),
.B(n_683),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1024),
.A2(n_772),
.B1(n_743),
.B2(n_799),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_913),
.B(n_823),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_901),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_959),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_906),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_906),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_949),
.A2(n_841),
.B(n_885),
.C(n_871),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_931),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_894),
.B(n_841),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_946),
.B(n_861),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_910),
.B(n_936),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_1024),
.A2(n_390),
.B1(n_359),
.B2(n_377),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_910),
.B(n_861),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_936),
.B(n_947),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_988),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_917),
.B(n_840),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_959),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_917),
.B(n_846),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_949),
.A2(n_813),
.B(n_742),
.C(n_784),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_983),
.B(n_871),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_903),
.A2(n_799),
.B1(n_784),
.B2(n_757),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_988),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_959),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_933),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_927),
.B(n_885),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1036),
.B(n_883),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_908),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1036),
.B(n_850),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_896),
.B(n_850),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1008),
.A2(n_812),
.B(n_853),
.C(n_851),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_933),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_962),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1028),
.A2(n_852),
.B(n_844),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_898),
.Y(n_1088)
);

OAI22x1_ASAP7_75t_L g1089 ( 
.A1(n_1008),
.A2(n_379),
.B1(n_385),
.B2(n_389),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_907),
.A2(n_837),
.B(n_851),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_1052),
.Y(n_1091)
);

INVx6_ASAP7_75t_L g1092 ( 
.A(n_959),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1053),
.B(n_853),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_998),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_997),
.B(n_502),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1031),
.A2(n_812),
.B(n_837),
.C(n_507),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_971),
.B(n_504),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_899),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_977),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_903),
.B(n_683),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_998),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_928),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_985),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_985),
.Y(n_1104)
);

BUFx4f_ASAP7_75t_L g1105 ( 
.A(n_978),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_989),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_989),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_909),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_971),
.B(n_504),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1007),
.B(n_333),
.Y(n_1110)
);

BUFx12f_ASAP7_75t_L g1111 ( 
.A(n_1002),
.Y(n_1111)
);

NOR2x1_ASAP7_75t_R g1112 ( 
.A(n_1003),
.B(n_379),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_SL g1113 ( 
.A(n_987),
.B(n_334),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_890),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1009),
.B(n_334),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1039),
.B(n_338),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_890),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_911),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1043),
.B(n_338),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1044),
.B(n_339),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1035),
.A2(n_391),
.B(n_389),
.C(n_390),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1045),
.B(n_339),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_921),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_978),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_912),
.B(n_506),
.Y(n_1126)
);

AO32x2_ASAP7_75t_L g1127 ( 
.A1(n_919),
.A2(n_719),
.A3(n_3),
.B1(n_10),
.B2(n_11),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_984),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_912),
.A2(n_360),
.B(n_396),
.C(n_394),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_978),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_980),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1051),
.B(n_344),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_1016),
.B(n_286),
.C(n_303),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_927),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_889),
.B(n_355),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1038),
.B(n_355),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1050),
.A2(n_360),
.B1(n_363),
.B2(n_396),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_935),
.B(n_363),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_939),
.A2(n_514),
.B(n_518),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_957),
.B(n_314),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_L g1141 ( 
.A(n_1016),
.B(n_507),
.C(n_317),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_926),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_974),
.B(n_428),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_932),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_914),
.A2(n_514),
.B(n_526),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_934),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_984),
.B(n_73),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_892),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_980),
.B(n_316),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1042),
.B(n_320),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1050),
.A2(n_324),
.B1(n_395),
.B2(n_391),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_905),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_915),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1042),
.B(n_514),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_957),
.B(n_902),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_973),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_891),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_902),
.B(n_948),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1027),
.B(n_940),
.Y(n_1159)
);

OAI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_953),
.A2(n_0),
.B(n_11),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_SL g1161 ( 
.A(n_1048),
.B(n_1049),
.C(n_893),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1042),
.B(n_149),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_951),
.B(n_0),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1042),
.B(n_144),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_893),
.A2(n_199),
.B1(n_195),
.B2(n_194),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1037),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_970),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_954),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_992),
.A2(n_182),
.B1(n_177),
.B2(n_171),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_R g1170 ( 
.A(n_1026),
.B(n_166),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1026),
.A2(n_581),
.B1(n_526),
.B2(n_17),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1014),
.A2(n_526),
.B1(n_581),
.B2(n_164),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_891),
.B(n_14),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_991),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1025),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_956),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_991),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_888),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_900),
.B(n_157),
.Y(n_1179)
);

O2A1O1Ixp5_ASAP7_75t_L g1180 ( 
.A1(n_1000),
.A2(n_155),
.B(n_151),
.C(n_140),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_891),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_922),
.B(n_137),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_SL g1183 ( 
.A1(n_929),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_967),
.B(n_15),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_960),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_904),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_916),
.A2(n_133),
.B(n_127),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_973),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_922),
.B(n_943),
.Y(n_1189)
);

NOR3xp33_ASAP7_75t_L g1190 ( 
.A(n_964),
.B(n_23),
.C(n_24),
.Y(n_1190)
);

NAND2xp33_ASAP7_75t_SL g1191 ( 
.A(n_891),
.B(n_23),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_916),
.A2(n_121),
.B(n_118),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_967),
.B(n_26),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1046),
.B(n_26),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1013),
.A2(n_116),
.B1(n_113),
.B2(n_106),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_904),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.C(n_38),
.Y(n_1196)
);

O2A1O1Ixp5_ASAP7_75t_L g1197 ( 
.A1(n_1000),
.A2(n_101),
.B(n_90),
.C(n_78),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1017),
.A2(n_1004),
.B(n_963),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_967),
.B(n_32),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1047),
.B(n_39),
.Y(n_1201)
);

CKINVDCx10_ASAP7_75t_R g1202 ( 
.A(n_942),
.Y(n_1202)
);

AOI22x1_ASAP7_75t_L g1203 ( 
.A1(n_1012),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1198),
.A2(n_1015),
.B(n_937),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1186),
.A2(n_993),
.B1(n_918),
.B2(n_900),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1081),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1155),
.B(n_1018),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1061),
.A2(n_895),
.B(n_1023),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1073),
.A2(n_924),
.A3(n_1019),
.B(n_1011),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1068),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1057),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1090),
.A2(n_1034),
.B(n_1054),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1097),
.B(n_929),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1155),
.B(n_1029),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1058),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1073),
.A2(n_961),
.B(n_1015),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1200),
.B(n_1029),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1081),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1168),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1069),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1095),
.B(n_994),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_1105),
.Y(n_1222)
);

AO22x2_ASAP7_75t_L g1223 ( 
.A1(n_1161),
.A2(n_961),
.B1(n_1010),
.B2(n_994),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1080),
.B(n_1030),
.Y(n_1224)
);

AO32x2_ASAP7_75t_L g1225 ( 
.A1(n_1075),
.A2(n_1032),
.A3(n_924),
.B1(n_969),
.B2(n_1041),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1176),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1083),
.A2(n_999),
.A3(n_1022),
.B(n_982),
.Y(n_1227)
);

NAND3xp33_ASAP7_75t_L g1228 ( 
.A(n_1141),
.B(n_995),
.C(n_1010),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1088),
.Y(n_1229)
);

BUFx4f_ASAP7_75t_L g1230 ( 
.A(n_1111),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_R g1231 ( 
.A(n_1102),
.B(n_1040),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1084),
.A2(n_993),
.B(n_979),
.C(n_950),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1186),
.A2(n_918),
.B1(n_900),
.B2(n_1040),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1056),
.B(n_923),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1098),
.Y(n_1235)
);

OA21x2_ASAP7_75t_L g1236 ( 
.A1(n_1100),
.A2(n_938),
.B(n_925),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1058),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1100),
.A2(n_981),
.B(n_986),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1099),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1064),
.B(n_996),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1139),
.A2(n_920),
.B(n_952),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1109),
.B(n_955),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_SL g1243 ( 
.A1(n_1082),
.A2(n_1192),
.B(n_1187),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1083),
.B(n_1001),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1055),
.A2(n_897),
.B1(n_888),
.B2(n_923),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1055),
.A2(n_1020),
.B(n_1033),
.Y(n_1246)
);

AO21x2_ASAP7_75t_L g1247 ( 
.A1(n_1070),
.A2(n_958),
.B(n_945),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1070),
.A2(n_1072),
.B(n_1063),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1131),
.B(n_1032),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_SL g1250 ( 
.A1(n_1194),
.A2(n_944),
.B(n_941),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1096),
.A2(n_968),
.B(n_897),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1140),
.B(n_955),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1140),
.B(n_923),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1158),
.B(n_923),
.Y(n_1254)
);

AO32x2_ASAP7_75t_L g1255 ( 
.A1(n_1165),
.A2(n_1041),
.A3(n_1021),
.B1(n_966),
.B2(n_972),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1059),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1166),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1134),
.Y(n_1258)
);

CKINVDCx6p67_ASAP7_75t_R g1259 ( 
.A(n_1202),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1074),
.B(n_955),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1158),
.B(n_1065),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1126),
.B(n_976),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1058),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1189),
.A2(n_1006),
.B(n_1005),
.Y(n_1264)
);

BUFx2_ASAP7_75t_SL g1265 ( 
.A(n_1134),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1195),
.A2(n_990),
.A3(n_975),
.B(n_1041),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1180),
.A2(n_1041),
.B(n_965),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_1069),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1078),
.B(n_955),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_SL g1270 ( 
.A1(n_1135),
.A2(n_1021),
.B(n_965),
.C(n_48),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1086),
.B(n_1002),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1108),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1060),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1105),
.A2(n_965),
.B(n_47),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1143),
.B(n_965),
.Y(n_1275)
);

BUFx4_ASAP7_75t_SL g1276 ( 
.A(n_1175),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1118),
.Y(n_1277)
);

OA22x2_ASAP7_75t_L g1278 ( 
.A1(n_1183),
.A2(n_1089),
.B1(n_1066),
.B2(n_1159),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1085),
.B(n_46),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1141),
.B(n_48),
.C(n_50),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1180),
.A2(n_50),
.B(n_55),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1197),
.A2(n_55),
.B(n_56),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1134),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1197),
.A2(n_59),
.B(n_60),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1123),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1156),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1133),
.A2(n_63),
.B(n_64),
.C(n_66),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1154),
.A2(n_67),
.B(n_68),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1067),
.A2(n_67),
.B(n_69),
.C(n_1160),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1171),
.A2(n_1196),
.B1(n_1146),
.B2(n_1144),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1062),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1071),
.B(n_1058),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1113),
.B(n_1136),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1110),
.B(n_1115),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1154),
.A2(n_1182),
.B(n_1164),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1182),
.A2(n_1162),
.B(n_1164),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1149),
.B(n_1076),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1145),
.A2(n_1079),
.B(n_1150),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1201),
.A2(n_1121),
.A3(n_1129),
.B(n_1163),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1156),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1071),
.B(n_1091),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1135),
.A2(n_1142),
.B(n_1093),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1174),
.B(n_1177),
.Y(n_1303)
);

AO32x2_ASAP7_75t_L g1304 ( 
.A1(n_1127),
.A2(n_1151),
.A3(n_1169),
.B1(n_1167),
.B2(n_1137),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1148),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1116),
.B(n_1132),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1156),
.B(n_1188),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1121),
.A2(n_1190),
.B(n_1163),
.C(n_1120),
.Y(n_1308)
);

BUFx8_ASAP7_75t_SL g1309 ( 
.A(n_1156),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1152),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1153),
.B(n_1185),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1076),
.Y(n_1312)
);

NAND2x1_ASAP7_75t_L g1313 ( 
.A(n_1092),
.B(n_1178),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1119),
.B(n_1122),
.Y(n_1314)
);

OAI22x1_ASAP7_75t_L g1315 ( 
.A1(n_1203),
.A2(n_1173),
.B1(n_1079),
.B2(n_1193),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1190),
.B(n_1173),
.C(n_1191),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1188),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1171),
.A2(n_1199),
.B(n_1184),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1094),
.B(n_1104),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1128),
.B(n_1170),
.Y(n_1320)
);

OAI22x1_ASAP7_75t_L g1321 ( 
.A1(n_1128),
.A2(n_1117),
.B1(n_1114),
.B2(n_1147),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1101),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1188),
.B(n_1147),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1179),
.A2(n_1188),
.B1(n_1138),
.B2(n_1077),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1077),
.B(n_1124),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1103),
.Y(n_1326)
);

OAI31xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1127),
.A2(n_1106),
.A3(n_1107),
.B(n_1179),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1157),
.A2(n_1172),
.B(n_1124),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1077),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1157),
.B(n_1181),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1092),
.B(n_1112),
.Y(n_1331)
);

AO32x2_ASAP7_75t_L g1332 ( 
.A1(n_1127),
.A2(n_1179),
.A3(n_1092),
.B1(n_1124),
.B2(n_1125),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1077),
.B(n_1124),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1125),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1125),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1125),
.B(n_1130),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1130),
.B(n_733),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1073),
.A2(n_1075),
.A3(n_1083),
.B(n_949),
.Y(n_1338)
);

BUFx8_ASAP7_75t_L g1339 ( 
.A(n_1111),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1155),
.B(n_1200),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1168),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1155),
.B(n_733),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1069),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1059),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1155),
.B(n_1200),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1155),
.B(n_1200),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1087),
.A2(n_917),
.B(n_1028),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1087),
.A2(n_917),
.B(n_1028),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1168),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1095),
.B(n_913),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1168),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1141),
.A2(n_731),
.B1(n_624),
.B2(n_414),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1095),
.B(n_913),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1087),
.A2(n_917),
.B(n_1028),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1168),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1081),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1314),
.A2(n_1342),
.B(n_1306),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1218),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1219),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1220),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1352),
.A2(n_1213),
.B1(n_1254),
.B2(n_1253),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1340),
.A2(n_1345),
.B1(n_1346),
.B2(n_1207),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1257),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1208),
.A2(n_1282),
.B(n_1281),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1298),
.A2(n_1212),
.B(n_1208),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1252),
.B(n_1214),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1278),
.A2(n_1316),
.B1(n_1280),
.B2(n_1233),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1238),
.A2(n_1243),
.B(n_1251),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1296),
.A2(n_1315),
.B(n_1248),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1340),
.A2(n_1346),
.B1(n_1345),
.B2(n_1261),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1293),
.A2(n_1278),
.B1(n_1294),
.B2(n_1318),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1281),
.A2(n_1282),
.B(n_1284),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1256),
.Y(n_1374)
);

NOR2x1_ASAP7_75t_R g1375 ( 
.A(n_1239),
.B(n_1211),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1226),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1273),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1327),
.A2(n_1246),
.B(n_1308),
.C(n_1284),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_1206),
.B(n_1356),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1276),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1210),
.B(n_1261),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1309),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1221),
.B(n_1260),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1229),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1231),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1246),
.A2(n_1232),
.B(n_1295),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1234),
.B(n_1297),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1233),
.A2(n_1205),
.B1(n_1301),
.B2(n_1324),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1307),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1214),
.A2(n_1210),
.B1(n_1205),
.B2(n_1323),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1235),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1291),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1258),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1264),
.A2(n_1328),
.B(n_1250),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1267),
.A2(n_1288),
.B(n_1245),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1240),
.B(n_1220),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1312),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1244),
.A2(n_1228),
.B(n_1217),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1267),
.A2(n_1245),
.B(n_1216),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1289),
.A2(n_1318),
.B1(n_1287),
.B2(n_1337),
.C(n_1274),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1279),
.A2(n_1324),
.B(n_1217),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1321),
.B(n_1265),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1216),
.A2(n_1236),
.B(n_1270),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1242),
.B(n_1320),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1247),
.A2(n_1302),
.B(n_1279),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1272),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1236),
.A2(n_1303),
.B(n_1325),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1290),
.A2(n_1240),
.B1(n_1223),
.B2(n_1262),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1303),
.A2(n_1269),
.B(n_1311),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1343),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1275),
.A2(n_1301),
.B1(n_1271),
.B2(n_1331),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1262),
.A2(n_1290),
.B(n_1224),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1269),
.A2(n_1311),
.B(n_1336),
.Y(n_1413)
);

NAND2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1329),
.B(n_1222),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1224),
.A2(n_1355),
.B(n_1351),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1247),
.A2(n_1302),
.B(n_1336),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1223),
.B(n_1222),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1258),
.Y(n_1418)
);

CKINVDCx6p67_ASAP7_75t_R g1419 ( 
.A(n_1300),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1209),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1322),
.B(n_1326),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1333),
.A2(n_1319),
.B(n_1313),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1277),
.A2(n_1349),
.B1(n_1285),
.B2(n_1341),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1330),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1330),
.B(n_1305),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_SL g1426 ( 
.A1(n_1335),
.A2(n_1332),
.B(n_1327),
.C(n_1310),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1344),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1227),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1299),
.B(n_1307),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1292),
.A2(n_1263),
.B(n_1215),
.Y(n_1430)
);

AOI221xp5_ASAP7_75t_L g1431 ( 
.A1(n_1249),
.A2(n_1230),
.B1(n_1338),
.B2(n_1317),
.C(n_1299),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1237),
.B(n_1263),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1237),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1299),
.B(n_1338),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1249),
.A2(n_1329),
.B(n_1334),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1230),
.A2(n_1286),
.B1(n_1283),
.B2(n_1258),
.Y(n_1436)
);

OR2x4_ASAP7_75t_L g1437 ( 
.A(n_1283),
.B(n_1286),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1283),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1266),
.A2(n_1227),
.B(n_1209),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1286),
.B(n_1329),
.Y(n_1440)
);

AO31x2_ASAP7_75t_L g1441 ( 
.A1(n_1225),
.A2(n_1332),
.A3(n_1255),
.B(n_1209),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1329),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1332),
.Y(n_1443)
);

OAI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1304),
.A2(n_1225),
.B1(n_1255),
.B2(n_1339),
.C(n_1259),
.Y(n_1444)
);

AOI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1255),
.A2(n_1225),
.B(n_1304),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1304),
.A2(n_1348),
.B(n_1347),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1339),
.B(n_1350),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1342),
.B(n_894),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1314),
.A2(n_930),
.B(n_894),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1342),
.A2(n_894),
.B1(n_1024),
.B2(n_1278),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1219),
.Y(n_1451)
);

INVx11_ASAP7_75t_L g1452 ( 
.A(n_1339),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1309),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1219),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1222),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1260),
.B(n_1234),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1219),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1253),
.B(n_930),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1347),
.A2(n_1354),
.B(n_1348),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1208),
.A2(n_1204),
.B(n_1281),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1342),
.A2(n_894),
.B1(n_1024),
.B2(n_1278),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1276),
.Y(n_1463)
);

AO21x1_ASAP7_75t_L g1464 ( 
.A1(n_1281),
.A2(n_1284),
.B(n_1282),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1259),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1352),
.A2(n_930),
.B1(n_731),
.B2(n_1213),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1241),
.A2(n_1198),
.B(n_1347),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1469)
);

AOI22x1_ASAP7_75t_SL g1470 ( 
.A1(n_1257),
.A2(n_638),
.B1(n_616),
.B2(n_1091),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1208),
.A2(n_1204),
.B(n_1281),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1219),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1241),
.A2(n_1198),
.B(n_1347),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1241),
.A2(n_1198),
.B(n_1347),
.Y(n_1474)
);

OR2x6_ASAP7_75t_L g1475 ( 
.A(n_1274),
.B(n_1324),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1327),
.A2(n_894),
.B(n_1024),
.C(n_1246),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1314),
.A2(n_930),
.B(n_894),
.Y(n_1478)
);

INVx4_ASAP7_75t_SL g1479 ( 
.A(n_1299),
.Y(n_1479)
);

AOI221x1_ASAP7_75t_L g1480 ( 
.A1(n_1281),
.A2(n_1284),
.B1(n_1282),
.B2(n_1141),
.C(n_1161),
.Y(n_1480)
);

OAI21xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1327),
.A2(n_1186),
.B(n_1055),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1210),
.B(n_1261),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1342),
.A2(n_894),
.B1(n_1024),
.B2(n_1278),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1352),
.A2(n_930),
.B1(n_731),
.B2(n_1213),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1212),
.A2(n_1073),
.A3(n_1075),
.B(n_1248),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1268),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1241),
.A2(n_1198),
.B(n_1347),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1347),
.A2(n_1100),
.B(n_1348),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1219),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1241),
.A2(n_1198),
.B(n_1347),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1352),
.A2(n_731),
.B1(n_414),
.B2(n_425),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1241),
.A2(n_1198),
.B(n_1347),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1220),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1257),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1342),
.A2(n_894),
.B1(n_1024),
.B2(n_1278),
.Y(n_1497)
);

INVx8_ASAP7_75t_L g1498 ( 
.A(n_1329),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1219),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1260),
.B(n_1234),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1222),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1502)
);

BUFx4f_ASAP7_75t_SL g1503 ( 
.A(n_1339),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1241),
.A2(n_1198),
.B(n_1347),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1219),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1219),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1219),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1219),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1309),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1483),
.B(n_1396),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1363),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1481),
.A2(n_1378),
.B(n_1477),
.C(n_1448),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1450),
.A2(n_1462),
.B1(n_1484),
.B2(n_1497),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1378),
.A2(n_1477),
.B(n_1448),
.C(n_1478),
.Y(n_1516)
);

INVxp33_ASAP7_75t_L g1517 ( 
.A(n_1404),
.Y(n_1517)
);

A2O1A1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1449),
.A2(n_1497),
.B(n_1450),
.C(n_1484),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1416),
.Y(n_1519)
);

AOI221x1_ASAP7_75t_SL g1520 ( 
.A1(n_1467),
.A2(n_1485),
.B1(n_1361),
.B2(n_1505),
.C(n_1488),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1480),
.A2(n_1446),
.B(n_1403),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1465),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1465),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1462),
.A2(n_1367),
.B1(n_1372),
.B2(n_1493),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1416),
.Y(n_1525)
);

O2A1O1Ixp5_ASAP7_75t_L g1526 ( 
.A1(n_1464),
.A2(n_1386),
.B(n_1357),
.C(n_1458),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1373),
.A2(n_1364),
.B(n_1458),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1429),
.B(n_1456),
.Y(n_1528)
);

O2A1O1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1400),
.A2(n_1362),
.B(n_1367),
.C(n_1371),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1403),
.A2(n_1368),
.B(n_1365),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1381),
.B(n_1459),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1424),
.B(n_1366),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1373),
.A2(n_1364),
.B(n_1412),
.Y(n_1533)
);

O2A1O1Ixp5_ASAP7_75t_L g1534 ( 
.A1(n_1370),
.A2(n_1366),
.B(n_1434),
.C(n_1390),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1425),
.B(n_1456),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1369),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1466),
.B(n_1469),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1437),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1401),
.A2(n_1475),
.B(n_1360),
.C(n_1495),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1425),
.B(n_1456),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1475),
.A2(n_1360),
.B(n_1495),
.C(n_1402),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1376),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1363),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1410),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1476),
.B(n_1482),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1410),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1500),
.B(n_1358),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1388),
.A2(n_1444),
.B(n_1408),
.C(n_1431),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1500),
.B(n_1421),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1411),
.A2(n_1408),
.B1(n_1379),
.B2(n_1436),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1475),
.A2(n_1402),
.B(n_1397),
.C(n_1423),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1487),
.A2(n_1414),
.B(n_1375),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1487),
.B(n_1427),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1496),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1503),
.Y(n_1556)
);

AOI21x1_ASAP7_75t_SL g1557 ( 
.A1(n_1447),
.A2(n_1420),
.B(n_1432),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1389),
.B(n_1374),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1417),
.B(n_1432),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1377),
.B(n_1392),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1384),
.Y(n_1561)
);

O2A1O1Ixp5_ASAP7_75t_L g1562 ( 
.A1(n_1490),
.A2(n_1435),
.B(n_1428),
.C(n_1423),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1391),
.A2(n_1472),
.B(n_1509),
.C(n_1508),
.Y(n_1563)
);

O2A1O1Ixp5_ASAP7_75t_L g1564 ( 
.A1(n_1428),
.A2(n_1442),
.B(n_1445),
.C(n_1440),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1455),
.A2(n_1501),
.B1(n_1385),
.B2(n_1506),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1385),
.A2(n_1463),
.B1(n_1380),
.B2(n_1496),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1418),
.Y(n_1567)
);

O2A1O1Ixp5_ASAP7_75t_L g1568 ( 
.A1(n_1440),
.A2(n_1457),
.B(n_1454),
.C(n_1451),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1406),
.A2(n_1507),
.B(n_1499),
.C(n_1491),
.Y(n_1569)
);

AOI211xp5_ASAP7_75t_L g1570 ( 
.A1(n_1426),
.A2(n_1365),
.B(n_1394),
.C(n_1433),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1407),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1479),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1443),
.A2(n_1409),
.B(n_1413),
.C(n_1399),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1415),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_SL g1575 ( 
.A1(n_1470),
.A2(n_1437),
.B(n_1503),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1368),
.A2(n_1439),
.B(n_1399),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1398),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1498),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1468),
.A2(n_1492),
.B(n_1474),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1426),
.A2(n_1414),
.B(n_1510),
.C(n_1453),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1468),
.A2(n_1492),
.B(n_1489),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1438),
.B(n_1393),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1382),
.A2(n_1453),
.B1(n_1510),
.B2(n_1452),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1405),
.B(n_1422),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1419),
.B(n_1486),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1430),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1405),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1486),
.B(n_1479),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1473),
.A2(n_1504),
.B(n_1494),
.Y(n_1589)
);

CKINVDCx14_ASAP7_75t_R g1590 ( 
.A(n_1382),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1461),
.B(n_1471),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1471),
.B(n_1441),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1441),
.B(n_1395),
.Y(n_1593)
);

O2A1O1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1504),
.A2(n_1342),
.B(n_949),
.C(n_1449),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1460),
.A2(n_1208),
.B(n_1386),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1429),
.B(n_1456),
.Y(n_1596)
);

AND2x2_ASAP7_75t_SL g1597 ( 
.A(n_1373),
.B(n_1327),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1378),
.A2(n_1386),
.B(n_1477),
.Y(n_1598)
);

O2A1O1Ixp5_ASAP7_75t_L g1599 ( 
.A1(n_1464),
.A2(n_1378),
.B(n_1477),
.C(n_1281),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1480),
.A2(n_1446),
.B(n_1378),
.Y(n_1601)
);

O2A1O1Ixp5_ASAP7_75t_L g1602 ( 
.A1(n_1464),
.A2(n_1378),
.B(n_1477),
.C(n_1281),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1450),
.A2(n_1352),
.B1(n_1484),
.B2(n_1462),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1449),
.A2(n_1342),
.B(n_949),
.C(n_1478),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1357),
.B(n_1371),
.Y(n_1607)
);

O2A1O1Ixp5_ASAP7_75t_L g1608 ( 
.A1(n_1464),
.A2(n_1378),
.B(n_1477),
.C(n_1281),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1467),
.A2(n_731),
.B1(n_1352),
.B2(n_1485),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1449),
.A2(n_1342),
.B(n_949),
.C(n_1478),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1363),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1429),
.B(n_1456),
.Y(n_1612)
);

OA21x2_ASAP7_75t_L g1613 ( 
.A1(n_1480),
.A2(n_1446),
.B(n_1378),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1477),
.A2(n_1233),
.B(n_1378),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_SL g1616 ( 
.A(n_1475),
.B(n_1417),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1477),
.A2(n_1233),
.B(n_1378),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1378),
.A2(n_1386),
.B(n_1477),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1429),
.B(n_1456),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1416),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1359),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1622)
);

O2A1O1Ixp5_ASAP7_75t_L g1623 ( 
.A1(n_1464),
.A2(n_1378),
.B(n_1477),
.C(n_1281),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1357),
.B(n_1371),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1450),
.A2(n_1352),
.B1(n_1484),
.B2(n_1462),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1378),
.A2(n_1386),
.B(n_1477),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1450),
.A2(n_1352),
.B1(n_1484),
.B2(n_1462),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1407),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1387),
.B(n_1383),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1574),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1593),
.B(n_1592),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1607),
.B(n_1624),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1614),
.B(n_1617),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1597),
.B(n_1591),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1571),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1542),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1577),
.B(n_1588),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1561),
.Y(n_1640)
);

AND2x4_ASAP7_75t_SL g1641 ( 
.A(n_1559),
.B(n_1572),
.Y(n_1641)
);

AO21x2_ASAP7_75t_L g1642 ( 
.A1(n_1587),
.A2(n_1618),
.B(n_1598),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1559),
.B(n_1616),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1517),
.B(n_1531),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1524),
.A2(n_1628),
.B1(n_1603),
.B2(n_1625),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1573),
.A2(n_1599),
.B(n_1623),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1627),
.B(n_1533),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1621),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1512),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1609),
.A2(n_1515),
.B1(n_1551),
.B2(n_1597),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1559),
.A2(n_1517),
.B1(n_1601),
.B2(n_1613),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1630),
.A2(n_1530),
.B(n_1581),
.Y(n_1652)
);

AOI222xp33_ASAP7_75t_L g1653 ( 
.A1(n_1516),
.A2(n_1518),
.B1(n_1514),
.B2(n_1548),
.C1(n_1536),
.C2(n_1583),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1576),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1586),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1613),
.B(n_1521),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1613),
.B(n_1521),
.Y(n_1657)
);

OR2x6_ASAP7_75t_L g1658 ( 
.A(n_1527),
.B(n_1541),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1544),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1546),
.B(n_1511),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1521),
.B(n_1573),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1563),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1516),
.B(n_1532),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1602),
.A2(n_1608),
.B(n_1562),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1519),
.A2(n_1525),
.B(n_1620),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1595),
.B(n_1514),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1605),
.A2(n_1610),
.B(n_1526),
.Y(n_1667)
);

OAI31xp33_ASAP7_75t_L g1668 ( 
.A1(n_1518),
.A2(n_1548),
.A3(n_1529),
.B(n_1594),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1554),
.B(n_1520),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1569),
.Y(n_1670)
);

INVxp67_ASAP7_75t_R g1671 ( 
.A(n_1565),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1534),
.A2(n_1564),
.B(n_1568),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1584),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1585),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1539),
.A2(n_1552),
.B(n_1580),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1595),
.B(n_1530),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1579),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1570),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1560),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1528),
.A2(n_1619),
.B1(n_1612),
.B2(n_1596),
.Y(n_1680)
);

OA21x2_ASAP7_75t_L g1681 ( 
.A1(n_1535),
.A2(n_1540),
.B(n_1612),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1596),
.B(n_1612),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1547),
.B(n_1545),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1632),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1645),
.A2(n_1513),
.B1(n_1629),
.B2(n_1626),
.C(n_1622),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1632),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1643),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1677),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1639),
.B(n_1589),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1665),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1643),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1633),
.B(n_1550),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1665),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1674),
.B(n_1537),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1674),
.B(n_1558),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1633),
.B(n_1549),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_SL g1698 ( 
.A(n_1647),
.B(n_1578),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1665),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1636),
.B(n_1631),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1655),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1634),
.B(n_1615),
.Y(n_1702)
);

AO21x2_ASAP7_75t_L g1703 ( 
.A1(n_1661),
.A2(n_1553),
.B(n_1557),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1665),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1634),
.B(n_1538),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1636),
.B(n_1606),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1660),
.B(n_1681),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1660),
.B(n_1600),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1635),
.B(n_1567),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1676),
.B(n_1604),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1681),
.B(n_1582),
.Y(n_1711)
);

AO221x2_ASAP7_75t_L g1712 ( 
.A1(n_1667),
.A2(n_1575),
.B1(n_1590),
.B2(n_1523),
.C(n_1522),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1637),
.B(n_1578),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1681),
.B(n_1567),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1636),
.B(n_1590),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1681),
.B(n_1679),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1661),
.B(n_1578),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1639),
.B(n_1673),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1673),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1681),
.B(n_1578),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1661),
.B(n_1566),
.Y(n_1721)
);

AO21x1_ASAP7_75t_SL g1722 ( 
.A1(n_1720),
.A2(n_1678),
.B(n_1675),
.Y(n_1722)
);

NAND2xp33_ASAP7_75t_R g1723 ( 
.A(n_1715),
.B(n_1635),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1719),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1719),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1718),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1688),
.B(n_1682),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1712),
.A2(n_1635),
.B1(n_1653),
.B2(n_1650),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1718),
.Y(n_1729)
);

OA222x2_ASAP7_75t_L g1730 ( 
.A1(n_1688),
.A2(n_1635),
.B1(n_1647),
.B2(n_1658),
.C1(n_1670),
.C2(n_1662),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1718),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1695),
.B(n_1644),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_R g1733 ( 
.A(n_1715),
.B(n_1522),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1684),
.Y(n_1734)
);

INVx3_ASAP7_75t_SL g1735 ( 
.A(n_1713),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1689),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1684),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1684),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1686),
.A2(n_1668),
.B1(n_1667),
.B2(n_1635),
.C(n_1653),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1715),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1687),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1689),
.Y(n_1742)
);

OAI31xp33_ASAP7_75t_L g1743 ( 
.A1(n_1721),
.A2(n_1668),
.A3(n_1678),
.B(n_1666),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1705),
.B(n_1635),
.C(n_1666),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1703),
.Y(n_1745)
);

AOI222xp33_ASAP7_75t_L g1746 ( 
.A1(n_1686),
.A2(n_1666),
.B1(n_1663),
.B2(n_1675),
.C1(n_1669),
.C2(n_1662),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1705),
.A2(n_1669),
.B1(n_1663),
.B2(n_1670),
.C(n_1651),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1688),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1702),
.A2(n_1695),
.B1(n_1721),
.B2(n_1707),
.C(n_1708),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1709),
.A2(n_1647),
.B1(n_1658),
.B2(n_1683),
.C(n_1680),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1721),
.A2(n_1646),
.B(n_1664),
.C(n_1672),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1712),
.A2(n_1647),
.B1(n_1664),
.B2(n_1646),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1715),
.A2(n_1523),
.B1(n_1556),
.B2(n_1543),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1709),
.A2(n_1647),
.B(n_1658),
.Y(n_1754)
);

OAI31xp33_ASAP7_75t_L g1755 ( 
.A1(n_1721),
.A2(n_1656),
.A3(n_1657),
.B(n_1683),
.Y(n_1755)
);

OAI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1708),
.A2(n_1671),
.B1(n_1647),
.B2(n_1658),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1688),
.B(n_1682),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1685),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1702),
.A2(n_1671),
.B1(n_1658),
.B2(n_1709),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1712),
.A2(n_1664),
.B1(n_1646),
.B2(n_1642),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1707),
.A2(n_1642),
.B1(n_1648),
.B2(n_1638),
.C(n_1640),
.Y(n_1761)
);

INVx3_ASAP7_75t_SL g1762 ( 
.A(n_1713),
.Y(n_1762)
);

AND4x1_ASAP7_75t_L g1763 ( 
.A(n_1712),
.B(n_1657),
.C(n_1656),
.D(n_1659),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1692),
.B(n_1682),
.Y(n_1764)
);

NAND3xp33_ASAP7_75t_L g1765 ( 
.A(n_1714),
.B(n_1646),
.C(n_1664),
.Y(n_1765)
);

AND2x2_ASAP7_75t_SL g1766 ( 
.A(n_1716),
.B(n_1646),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1700),
.A2(n_1658),
.B1(n_1682),
.B2(n_1641),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1734),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1737),
.Y(n_1769)
);

INVx4_ASAP7_75t_SL g1770 ( 
.A(n_1735),
.Y(n_1770)
);

INVxp67_ASAP7_75t_SL g1771 ( 
.A(n_1758),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1738),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1758),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1741),
.Y(n_1774)
);

INVx4_ASAP7_75t_SL g1775 ( 
.A(n_1735),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1728),
.A2(n_1712),
.B(n_1717),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1736),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1749),
.B(n_1710),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1724),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1736),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_SL g1781 ( 
.A1(n_1739),
.A2(n_1712),
.B(n_1698),
.Y(n_1781)
);

OAI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1754),
.A2(n_1652),
.B(n_1654),
.Y(n_1782)
);

OAI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1743),
.A2(n_1720),
.B(n_1714),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1742),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1726),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1762),
.B(n_1692),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1733),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1744),
.B(n_1703),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1765),
.A2(n_1704),
.B(n_1694),
.Y(n_1789)
);

INVx4_ASAP7_75t_SL g1790 ( 
.A(n_1762),
.Y(n_1790)
);

INVx4_ASAP7_75t_SL g1791 ( 
.A(n_1748),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1729),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1731),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1725),
.Y(n_1794)
);

AO21x2_ASAP7_75t_L g1795 ( 
.A1(n_1763),
.A2(n_1694),
.B(n_1691),
.Y(n_1795)
);

INVx4_ASAP7_75t_SL g1796 ( 
.A(n_1748),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1733),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1747),
.A2(n_1717),
.B(n_1711),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1727),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1732),
.B(n_1710),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1766),
.B(n_1700),
.Y(n_1801)
);

INVxp67_ASAP7_75t_SL g1802 ( 
.A(n_1723),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1779),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1768),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1798),
.B(n_1700),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1797),
.B(n_1753),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1770),
.B(n_1722),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1770),
.B(n_1722),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1801),
.B(n_1716),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1785),
.B(n_1711),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1794),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1770),
.B(n_1727),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1768),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1787),
.Y(n_1814)
);

NOR4xp75_ASAP7_75t_L g1815 ( 
.A(n_1783),
.B(n_1759),
.C(n_1750),
.D(n_1767),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1770),
.B(n_1730),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1800),
.B(n_1706),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1555),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1769),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1794),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1785),
.B(n_1690),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1775),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1769),
.Y(n_1823)
);

NOR2xp67_ASAP7_75t_L g1824 ( 
.A(n_1799),
.B(n_1745),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1778),
.B(n_1706),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1775),
.B(n_1757),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1792),
.B(n_1690),
.Y(n_1827)
);

OAI31xp33_ASAP7_75t_L g1828 ( 
.A1(n_1776),
.A2(n_1756),
.A3(n_1751),
.B(n_1755),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1775),
.B(n_1757),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_R g1830 ( 
.A(n_1799),
.B(n_1556),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1777),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1771),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1775),
.B(n_1757),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1802),
.B(n_1555),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1773),
.B(n_1706),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1790),
.B(n_1791),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1781),
.Y(n_1837)
);

NAND2x1p5_ASAP7_75t_L g1838 ( 
.A(n_1788),
.B(n_1745),
.Y(n_1838)
);

OR2x6_ASAP7_75t_L g1839 ( 
.A(n_1781),
.B(n_1745),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1792),
.B(n_1690),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1790),
.B(n_1746),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1793),
.B(n_1693),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_L g1843 ( 
.A(n_1782),
.B(n_1761),
.C(n_1699),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1793),
.B(n_1740),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1772),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1791),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1772),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1790),
.B(n_1764),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1811),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1826),
.B(n_1790),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1836),
.B(n_1791),
.Y(n_1851)
);

OAI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1837),
.A2(n_1723),
.B1(n_1664),
.B2(n_1712),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1814),
.B(n_1696),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1825),
.B(n_1696),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1820),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1832),
.B(n_1697),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1697),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1837),
.A2(n_1672),
.B1(n_1789),
.B2(n_1701),
.Y(n_1858)
);

INVxp33_ASAP7_75t_L g1859 ( 
.A(n_1806),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1819),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1836),
.B(n_1791),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1819),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1835),
.B(n_1697),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1845),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1818),
.B(n_1543),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1845),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1804),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1842),
.B(n_1697),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1813),
.Y(n_1869)
);

NAND3xp33_ASAP7_75t_L g1870 ( 
.A(n_1841),
.B(n_1760),
.C(n_1752),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1831),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1823),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1803),
.B(n_1766),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1817),
.B(n_1799),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1807),
.B(n_1796),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1812),
.B(n_1796),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1847),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1831),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1821),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1846),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1826),
.B(n_1786),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1821),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1809),
.B(n_1774),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1827),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1827),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1880),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1880),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1875),
.B(n_1850),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1860),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1859),
.B(n_1834),
.Y(n_1890)
);

INVx3_ASAP7_75t_SL g1891 ( 
.A(n_1851),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1875),
.B(n_1816),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1851),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1851),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1881),
.B(n_1816),
.Y(n_1895)
);

AND2x4_ASAP7_75t_SL g1896 ( 
.A(n_1876),
.B(n_1807),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1859),
.B(n_1865),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1849),
.B(n_1810),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1855),
.B(n_1856),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1862),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1865),
.B(n_1861),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_SL g1902 ( 
.A(n_1876),
.B(n_1808),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1876),
.Y(n_1903)
);

CKINVDCx16_ASAP7_75t_R g1904 ( 
.A(n_1861),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1861),
.B(n_1808),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1884),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1884),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1864),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1866),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1871),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1867),
.B(n_1822),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1871),
.Y(n_1912)
);

NOR2x1p5_ASAP7_75t_L g1913 ( 
.A(n_1870),
.B(n_1812),
.Y(n_1913)
);

OAI22xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1904),
.A2(n_1839),
.B1(n_1611),
.B2(n_1838),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1897),
.B(n_1869),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1906),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1890),
.A2(n_1828),
.B(n_1858),
.Y(n_1917)
);

AOI221x1_ASAP7_75t_L g1918 ( 
.A1(n_1886),
.A2(n_1843),
.B1(n_1878),
.B2(n_1872),
.C(n_1877),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1893),
.B(n_1853),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1902),
.A2(n_1852),
.B1(n_1839),
.B2(n_1812),
.Y(n_1920)
);

NAND4xp25_ASAP7_75t_SL g1921 ( 
.A(n_1888),
.B(n_1873),
.C(n_1833),
.D(n_1829),
.Y(n_1921)
);

INVxp33_ASAP7_75t_L g1922 ( 
.A(n_1901),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1888),
.B(n_1649),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1913),
.A2(n_1839),
.B1(n_1852),
.B2(n_1838),
.Y(n_1924)
);

OAI31xp33_ASAP7_75t_L g1925 ( 
.A1(n_1896),
.A2(n_1838),
.A3(n_1858),
.B(n_1815),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1894),
.B(n_1879),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1906),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1906),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1886),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1892),
.A2(n_1839),
.B1(n_1848),
.B2(n_1833),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1891),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1887),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1891),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1892),
.A2(n_1830),
.B1(n_1752),
.B2(n_1795),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1887),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1927),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1927),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1928),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1931),
.B(n_1903),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1931),
.B(n_1903),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1933),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1933),
.B(n_1905),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1922),
.B(n_1891),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1917),
.B(n_1905),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1925),
.B(n_1896),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1928),
.Y(n_1946)
);

INVxp67_ASAP7_75t_L g1947 ( 
.A(n_1923),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1926),
.B(n_1895),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1916),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1945),
.A2(n_1921),
.B1(n_1914),
.B2(n_1923),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1944),
.A2(n_1934),
.B1(n_1930),
.B2(n_1920),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1942),
.B(n_1929),
.Y(n_1952)
);

AOI322xp5_ASAP7_75t_L g1953 ( 
.A1(n_1945),
.A2(n_1915),
.A3(n_1934),
.B1(n_1932),
.B2(n_1935),
.C1(n_1919),
.C2(n_1895),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1942),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1948),
.A2(n_1924),
.B1(n_1899),
.B2(n_1911),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1943),
.A2(n_1918),
.B(n_1907),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1941),
.B(n_1907),
.Y(n_1957)
);

OAI21xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1947),
.A2(n_1899),
.B(n_1908),
.Y(n_1958)
);

O2A1O1Ixp5_ASAP7_75t_SL g1959 ( 
.A1(n_1936),
.A2(n_1889),
.B(n_1900),
.C(n_1909),
.Y(n_1959)
);

OAI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1939),
.A2(n_1898),
.B1(n_1829),
.B2(n_1848),
.Y(n_1960)
);

AOI211xp5_ASAP7_75t_SL g1961 ( 
.A1(n_1940),
.A2(n_1912),
.B(n_1910),
.C(n_1889),
.Y(n_1961)
);

NOR2x1_ASAP7_75t_L g1962 ( 
.A(n_1937),
.B(n_1900),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1954),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1950),
.B(n_1898),
.Y(n_1964)
);

O2A1O1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1956),
.A2(n_1949),
.B(n_1946),
.C(n_1938),
.Y(n_1965)
);

AOI211xp5_ASAP7_75t_L g1966 ( 
.A1(n_1951),
.A2(n_1909),
.B(n_1910),
.C(n_1912),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1957),
.B(n_1882),
.Y(n_1967)
);

AOI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1958),
.A2(n_1885),
.B(n_1883),
.Y(n_1968)
);

A2O1A1Ixp33_ASAP7_75t_SL g1969 ( 
.A1(n_1961),
.A2(n_1885),
.B(n_1760),
.C(n_1774),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1962),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1970),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1963),
.B(n_1953),
.Y(n_1972)
);

NOR2xp67_ASAP7_75t_L g1973 ( 
.A(n_1968),
.B(n_1952),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1964),
.B(n_1960),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1967),
.B(n_1955),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1965),
.B(n_1959),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1969),
.B(n_1874),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1966),
.Y(n_1978)
);

O2A1O1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1972),
.A2(n_1824),
.B(n_1789),
.C(n_1795),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1971),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1975),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1973),
.B(n_1854),
.Y(n_1982)
);

NOR2x1_ASAP7_75t_L g1983 ( 
.A(n_1976),
.B(n_1795),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1974),
.B(n_1857),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1981),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1982),
.B(n_1978),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1983),
.Y(n_1987)
);

NOR2x1_ASAP7_75t_L g1988 ( 
.A(n_1987),
.B(n_1980),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1988),
.A2(n_1977),
.B1(n_1985),
.B2(n_1984),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1989),
.B(n_1986),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1989),
.Y(n_1991)
);

XNOR2x1_ASAP7_75t_SL g1992 ( 
.A(n_1991),
.B(n_1979),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1990),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1993),
.A2(n_1796),
.B1(n_1789),
.B2(n_1809),
.Y(n_1994)
);

CKINVDCx20_ASAP7_75t_R g1995 ( 
.A(n_1992),
.Y(n_1995)
);

NOR2x1_ASAP7_75t_L g1996 ( 
.A(n_1995),
.B(n_1844),
.Y(n_1996)
);

NOR2xp67_ASAP7_75t_L g1997 ( 
.A(n_1996),
.B(n_1994),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1997),
.B(n_1863),
.Y(n_1998)
);

AO221x2_ASAP7_75t_L g1999 ( 
.A1(n_1998),
.A2(n_1796),
.B1(n_1777),
.B2(n_1780),
.C(n_1784),
.Y(n_1999)
);

OAI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1999),
.A2(n_1840),
.B1(n_1844),
.B2(n_1810),
.Y(n_2000)
);

AOI211xp5_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1840),
.B(n_1782),
.C(n_1868),
.Y(n_2001)
);


endmodule