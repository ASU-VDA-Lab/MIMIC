module fake_jpeg_3263_n_725 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_725);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_725;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_716;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_717;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_718;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_723;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_715;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_720;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_714;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_724;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_719;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_722;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_721;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_68),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_69),
.Y(n_194)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_72),
.Y(n_216)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_73),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_75),
.Y(n_203)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_21),
.B(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_112),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_10),
.B(n_18),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_82),
.B(n_117),
.C(n_56),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_84),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_91),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_21),
.B(n_10),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_97),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_93),
.Y(n_213)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_94),
.Y(n_217)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_96),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_23),
.B(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_40),
.Y(n_136)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_99),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_100),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_33),
.Y(n_102)
);

INVx5_ASAP7_75t_SL g157 ( 
.A(n_102),
.Y(n_157)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_110),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_39),
.B(n_18),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_46),
.B(n_18),
.C(n_16),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

CKINVDCx6p67_ASAP7_75t_R g119 ( 
.A(n_48),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_132),
.C(n_133),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_124),
.B(n_128),
.Y(n_211)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_37),
.Y(n_125)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_37),
.Y(n_126)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_23),
.B(n_16),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_26),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_37),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_136),
.B(n_139),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_55),
.B1(n_57),
.B2(n_42),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_137),
.A2(n_144),
.B1(n_152),
.B2(n_187),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_40),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_51),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_143),
.B(n_146),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_70),
.A2(n_52),
.B1(n_51),
.B2(n_47),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_52),
.Y(n_146)
);

HAxp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_48),
.CON(n_147),
.SN(n_147)
);

NAND2x1_ASAP7_75t_SL g274 ( 
.A(n_147),
.B(n_0),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_76),
.A2(n_50),
.B1(n_37),
.B2(n_55),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_151),
.A2(n_185),
.B1(n_190),
.B2(n_38),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_55),
.B1(n_57),
.B2(n_42),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_50),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_154),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_101),
.B(n_47),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_158),
.B(n_162),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_161),
.B(n_177),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_71),
.B(n_39),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_27),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_99),
.B(n_50),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_178),
.B(n_180),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_50),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_65),
.A2(n_27),
.B1(n_26),
.B2(n_61),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_181),
.B(n_189),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_50),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_183),
.B(n_186),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_90),
.A2(n_50),
.B1(n_27),
.B2(n_26),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_20),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_67),
.A2(n_61),
.B1(n_25),
.B2(n_28),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_108),
.B(n_61),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_90),
.A2(n_20),
.B1(n_25),
.B2(n_53),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_109),
.B(n_20),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_196),
.B(n_214),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_197),
.B(n_14),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_111),
.A2(n_25),
.B1(n_28),
.B2(n_53),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_199),
.A2(n_209),
.B1(n_35),
.B2(n_2),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_91),
.B(n_53),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_206),
.B(n_222),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_114),
.A2(n_56),
.B1(n_54),
.B2(n_38),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_115),
.B(n_31),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_94),
.B(n_31),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_120),
.B(n_31),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_227),
.B(n_1),
.Y(n_304)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g314 ( 
.A(n_228),
.Y(n_314)
);

OA22x2_ASAP7_75t_L g362 ( 
.A1(n_230),
.A2(n_234),
.B1(n_306),
.B2(n_3),
.Y(n_362)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_145),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_231),
.Y(n_353)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_232),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_152),
.B1(n_137),
.B2(n_133),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_233),
.A2(n_216),
.B1(n_170),
.B2(n_175),
.Y(n_340)
);

AO22x2_ASAP7_75t_L g234 ( 
.A1(n_147),
.A2(n_38),
.B1(n_54),
.B2(n_56),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g235 ( 
.A1(n_154),
.A2(n_132),
.B1(n_130),
.B2(n_123),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_259),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_148),
.A2(n_28),
.B1(n_54),
.B2(n_34),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_236),
.Y(n_341)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_238),
.Y(n_370)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_240),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_135),
.A2(n_79),
.B1(n_100),
.B2(n_93),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_242),
.Y(n_364)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_245),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_246),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_166),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_247),
.Y(n_331)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_176),
.Y(n_248)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_148),
.A2(n_34),
.B1(n_69),
.B2(n_87),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_249),
.A2(n_251),
.B1(n_276),
.B2(n_280),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_164),
.A2(n_179),
.B1(n_34),
.B2(n_166),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_252),
.Y(n_342)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_150),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_172),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_258),
.Y(n_318)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_257),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_138),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

INVx6_ASAP7_75t_L g356 ( 
.A(n_260),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_185),
.A2(n_116),
.B(n_127),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_263),
.A2(n_149),
.B(n_2),
.Y(n_355)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_167),
.Y(n_264)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g265 ( 
.A1(n_153),
.A2(n_104),
.A3(n_86),
.B1(n_80),
.B2(n_74),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_265),
.A2(n_11),
.B(n_5),
.Y(n_366)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_184),
.Y(n_267)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_140),
.B(n_0),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_268),
.B(n_273),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_211),
.Y(n_269)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_270),
.Y(n_365)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_271),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_223),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_275),
.Y(n_324)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_274),
.B(n_289),
.C(n_296),
.Y(n_349)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_219),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_164),
.A2(n_72),
.B1(n_35),
.B2(n_24),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_193),
.Y(n_277)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_134),
.B(n_1),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_278),
.B(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_282),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_179),
.A2(n_35),
.B1(n_16),
.B2(n_15),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_155),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_281),
.A2(n_293),
.B1(n_297),
.B2(n_299),
.Y(n_329)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_224),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_286),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_208),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_288),
.B(n_290),
.Y(n_359)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_167),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g291 ( 
.A(n_226),
.Y(n_291)
);

CKINVDCx9p33_ASAP7_75t_R g348 ( 
.A(n_291),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_212),
.B(n_14),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_211),
.A2(n_226),
.B1(n_207),
.B2(n_203),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_294),
.B(n_295),
.Y(n_373)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_171),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_212),
.B(n_13),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_150),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_171),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_300),
.A2(n_301),
.B1(n_308),
.B2(n_193),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_201),
.Y(n_301)
);

INVx3_ASAP7_75t_SL g302 ( 
.A(n_160),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_302),
.A2(n_303),
.B1(n_216),
.B2(n_198),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_202),
.B(n_12),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_305),
.Y(n_315)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_194),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_169),
.B(n_1),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_309),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_194),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_192),
.B(n_1),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_269),
.A2(n_163),
.B1(n_200),
.B2(n_199),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_313),
.A2(n_333),
.B1(n_339),
.B2(n_268),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_250),
.A2(n_173),
.B1(n_200),
.B2(n_195),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_319),
.A2(n_368),
.B1(n_242),
.B2(n_274),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_287),
.A2(n_225),
.B1(n_213),
.B2(n_217),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_261),
.A2(n_220),
.B1(n_157),
.B2(n_201),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_337),
.A2(n_345),
.B1(n_360),
.B2(n_240),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_250),
.A2(n_151),
.B1(n_190),
.B2(n_195),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_338),
.A2(n_363),
.B1(n_366),
.B2(n_232),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_287),
.A2(n_225),
.B1(n_213),
.B2(n_217),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_340),
.A2(n_263),
.B1(n_308),
.B2(n_260),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_175),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_350),
.Y(n_376)
);

OR2x2_ASAP7_75t_SL g344 ( 
.A(n_229),
.B(n_198),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_344),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_262),
.A2(n_198),
.B1(n_165),
.B2(n_215),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_283),
.B(n_170),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_352),
.Y(n_380)
);

OAI32xp33_ASAP7_75t_L g354 ( 
.A1(n_285),
.A2(n_149),
.A3(n_160),
.B1(n_215),
.B2(n_165),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_357),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_355),
.A2(n_368),
.B(n_320),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_1),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_307),
.B(n_3),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_369),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_299),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_362),
.B(n_4),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_306),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_235),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_4),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g374 ( 
.A(n_325),
.B(n_268),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_374),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_364),
.A2(n_338),
.B1(n_325),
.B2(n_341),
.Y(n_375)
);

NOR2x1_ASAP7_75t_L g460 ( 
.A(n_375),
.B(n_404),
.Y(n_460)
);

OAI32xp33_ASAP7_75t_L g379 ( 
.A1(n_325),
.A2(n_298),
.A3(n_259),
.B1(n_241),
.B2(n_265),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_392),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_334),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_381),
.B(n_393),
.Y(n_446)
);

INVxp33_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_373),
.Y(n_383)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_384),
.A2(n_348),
.B1(n_342),
.B2(n_326),
.Y(n_457)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_324),
.Y(n_385)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_388),
.A2(n_401),
.B1(n_409),
.B2(n_413),
.Y(n_426)
);

OAI22x1_ASAP7_75t_L g389 ( 
.A1(n_319),
.A2(n_234),
.B1(n_259),
.B2(n_254),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_389),
.A2(n_404),
.B1(n_327),
.B2(n_245),
.Y(n_466)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_353),
.B(n_243),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_395),
.B(n_410),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_321),
.B(n_253),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_398),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_278),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_397),
.B(n_399),
.C(n_414),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_278),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_343),
.B(n_239),
.C(n_248),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_234),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_403),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_366),
.A2(n_305),
.B1(n_295),
.B2(n_255),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_332),
.Y(n_402)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_402),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_315),
.B(n_234),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_318),
.B(n_270),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_407),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_406),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_315),
.B(n_284),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_341),
.A2(n_257),
.B1(n_252),
.B2(n_297),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_364),
.A2(n_275),
.B1(n_271),
.B2(n_281),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_359),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_411),
.Y(n_443)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_361),
.Y(n_412)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_355),
.A2(n_300),
.B1(n_302),
.B2(n_294),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_SL g414 ( 
.A(n_347),
.B(n_238),
.C(n_277),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_415),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_328),
.B(n_247),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_369),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_372),
.Y(n_417)
);

INVx11_ASAP7_75t_L g448 ( 
.A(n_417),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_418),
.A2(n_349),
.B1(n_351),
.B2(n_328),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_372),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_421),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_420),
.A2(n_329),
.B(n_348),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_331),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_331),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_291),
.Y(n_452)
);

INVx3_ASAP7_75t_SL g424 ( 
.A(n_330),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g427 ( 
.A(n_381),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_427),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_378),
.A2(n_418),
.B1(n_375),
.B2(n_400),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_433),
.A2(n_435),
.B1(n_439),
.B2(n_389),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_378),
.A2(n_362),
.B1(n_354),
.B2(n_351),
.Y(n_435)
);

AO21x2_ASAP7_75t_L g436 ( 
.A1(n_413),
.A2(n_363),
.B(n_362),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_436),
.A2(n_438),
.B1(n_457),
.B2(n_464),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_376),
.A2(n_362),
.B1(n_351),
.B2(n_352),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_405),
.Y(n_440)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_387),
.Y(n_451)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g498 ( 
.A(n_452),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_376),
.B(n_358),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_391),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_454),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_460),
.A2(n_462),
.B(n_408),
.Y(n_502)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_380),
.A2(n_322),
.B1(n_311),
.B2(n_346),
.Y(n_464)
);

OAI22x1_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_422),
.B1(n_414),
.B2(n_424),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_460),
.A2(n_404),
.B(n_403),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_468),
.A2(n_482),
.B(n_483),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_428),
.B(n_397),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_428),
.Y(n_508)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_474),
.Y(n_511)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_475),
.Y(n_521)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_462),
.A2(n_420),
.B(n_423),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_477),
.A2(n_494),
.B(n_465),
.Y(n_541)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_434),
.Y(n_478)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_478),
.Y(n_531)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_442),
.Y(n_480)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_480),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_436),
.A2(n_404),
.B1(n_380),
.B2(n_384),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_481),
.A2(n_489),
.B1(n_491),
.B2(n_440),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_460),
.A2(n_377),
.B(n_393),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_429),
.A2(n_377),
.B(n_406),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_452),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_484),
.B(n_486),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_SL g485 ( 
.A1(n_438),
.A2(n_421),
.B1(n_385),
.B2(n_383),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_488),
.B1(n_493),
.B2(n_495),
.Y(n_507)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_451),
.Y(n_487)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_487),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_436),
.A2(n_374),
.B1(n_407),
.B2(n_379),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_454),
.C(n_455),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_505),
.C(n_430),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_436),
.A2(n_374),
.B1(n_396),
.B2(n_389),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_453),
.B(n_391),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_492),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_436),
.A2(n_401),
.B1(n_388),
.B2(n_416),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_436),
.A2(n_409),
.B1(n_422),
.B2(n_419),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_429),
.A2(n_455),
.B(n_446),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_497),
.A2(n_398),
.B(n_449),
.Y(n_544)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_499),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_464),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_501),
.B(n_443),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_SL g529 ( 
.A1(n_502),
.A2(n_456),
.B(n_458),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_439),
.A2(n_422),
.B1(n_410),
.B2(n_417),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_503),
.A2(n_495),
.B1(n_456),
.B2(n_477),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_432),
.B(n_399),
.Y(n_504)
);

CKINVDCx14_ASAP7_75t_R g520 ( 
.A(n_504),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_444),
.B(n_374),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_493),
.A2(n_425),
.B1(n_466),
.B2(n_426),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_506),
.A2(n_517),
.B1(n_540),
.B2(n_481),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_508),
.B(n_530),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_509),
.A2(n_541),
.B(n_542),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_496),
.B(n_431),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_512),
.B(n_357),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_498),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_513),
.B(n_519),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_433),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_514),
.B(n_523),
.Y(n_562)
);

AO22x1_ASAP7_75t_L g515 ( 
.A1(n_474),
.A2(n_435),
.B1(n_448),
.B2(n_446),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_SL g578 ( 
.A1(n_515),
.A2(n_447),
.B(n_441),
.C(n_365),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_470),
.B(n_425),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_L g560 ( 
.A(n_516),
.B(n_532),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_488),
.A2(n_426),
.B1(n_456),
.B2(n_445),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_518),
.B(n_528),
.C(n_471),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_497),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_432),
.Y(n_523)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_524),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_469),
.B(n_430),
.C(n_431),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_467),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_469),
.B(n_463),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_504),
.B(n_486),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_482),
.B(n_463),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_533),
.B(n_539),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_534),
.A2(n_480),
.B1(n_478),
.B2(n_476),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_503),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_535),
.B(n_472),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_492),
.B(n_392),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_475),
.A2(n_443),
.B1(n_465),
.B2(n_448),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_502),
.A2(n_448),
.B(n_450),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_544),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_537),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_545),
.B(n_550),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_546),
.A2(n_555),
.B1(n_569),
.B2(n_576),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_548),
.A2(n_571),
.B(n_580),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_544),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_552),
.B(n_577),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_471),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_553),
.B(n_557),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_507),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_554),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_506),
.A2(n_517),
.B1(n_515),
.B2(n_491),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_522),
.Y(n_556)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_556),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_537),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_511),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_558),
.B(n_570),
.Y(n_594)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_522),
.Y(n_559)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_559),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_489),
.Y(n_565)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_565),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_540),
.Y(n_566)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_566),
.Y(n_603)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_525),
.Y(n_567)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_567),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_541),
.A2(n_468),
.B(n_483),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_568),
.A2(n_572),
.B(n_575),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_515),
.A2(n_494),
.B1(n_484),
.B2(n_500),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_510),
.A2(n_479),
.B1(n_499),
.B2(n_487),
.Y(n_570)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_573),
.A2(n_543),
.B1(n_531),
.B2(n_459),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_542),
.A2(n_473),
.B(n_472),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_574),
.A2(n_579),
.B(n_526),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_520),
.A2(n_473),
.B1(n_501),
.B2(n_450),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_510),
.B(n_447),
.Y(n_577)
);

A2O1A1Ixp33_ASAP7_75t_SL g598 ( 
.A1(n_578),
.A2(n_543),
.B(n_536),
.C(n_531),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_L g579 ( 
.A(n_539),
.B(n_441),
.Y(n_579)
);

O2A1O1Ixp33_ASAP7_75t_SL g580 ( 
.A1(n_511),
.A2(n_346),
.B(n_322),
.C(n_311),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_532),
.B(n_316),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_581),
.B(n_563),
.Y(n_602)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_583),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_552),
.B(n_518),
.C(n_514),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_584),
.B(n_588),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_523),
.C(n_530),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_562),
.B(n_516),
.C(n_533),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_591),
.B(n_592),
.C(n_596),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_547),
.B(n_526),
.C(n_521),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_549),
.A2(n_534),
.B(n_521),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_595),
.A2(n_598),
.B(n_578),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_547),
.B(n_527),
.C(n_538),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_546),
.A2(n_527),
.B1(n_538),
.B2(n_536),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_597),
.A2(n_606),
.B1(n_556),
.B2(n_559),
.Y(n_617)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_599),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_560),
.B(n_415),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_601),
.B(n_610),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_SL g622 ( 
.A(n_602),
.B(n_564),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_316),
.C(n_365),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_605),
.B(n_608),
.C(n_611),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_554),
.A2(n_424),
.B1(n_459),
.B2(n_390),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_560),
.B(n_402),
.C(n_386),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_568),
.B(n_412),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_566),
.B(n_330),
.C(n_370),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_576),
.B(n_371),
.C(n_370),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_574),
.C(n_572),
.Y(n_625)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_613),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_617),
.Y(n_641)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_604),
.Y(n_618)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_618),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_600),
.B(n_551),
.Y(n_620)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_620),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_622),
.B(n_623),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_592),
.B(n_561),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_587),
.A2(n_551),
.B1(n_545),
.B2(n_573),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_624),
.A2(n_630),
.B1(n_585),
.B2(n_611),
.Y(n_646)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_625),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g626 ( 
.A(n_588),
.B(n_561),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_626),
.B(n_627),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_548),
.Y(n_627)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_609),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_629),
.B(n_632),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_590),
.A2(n_548),
.B1(n_555),
.B2(n_567),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_586),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_637),
.Y(n_652)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_582),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_584),
.B(n_569),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_633),
.B(n_635),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_577),
.C(n_558),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_634),
.B(n_639),
.C(n_612),
.Y(n_648)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_589),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_596),
.B(n_578),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_636),
.B(n_638),
.Y(n_659)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_595),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_605),
.B(n_578),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_583),
.B(n_580),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_614),
.A2(n_590),
.B1(n_603),
.B2(n_607),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g676 ( 
.A1(n_643),
.A2(n_647),
.B1(n_650),
.B2(n_356),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_613),
.A2(n_585),
.B(n_598),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_644),
.A2(n_651),
.B(n_638),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_646),
.A2(n_653),
.B1(n_615),
.B2(n_342),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_616),
.A2(n_597),
.B1(n_594),
.B2(n_610),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_648),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_639),
.A2(n_599),
.B1(n_598),
.B2(n_601),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_623),
.A2(n_598),
.B(n_606),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_SL g653 ( 
.A1(n_627),
.A2(n_608),
.B1(n_602),
.B2(n_591),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_633),
.B(n_326),
.C(n_327),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_654),
.B(n_656),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_619),
.B(n_367),
.C(n_371),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_619),
.B(n_367),
.C(n_361),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_657),
.B(n_314),
.Y(n_678)
);

BUFx24_ASAP7_75t_SL g661 ( 
.A(n_628),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_661),
.B(n_656),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_662),
.B(n_634),
.C(n_626),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_663),
.B(n_664),
.Y(n_690)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_642),
.B(n_621),
.C(n_636),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_660),
.Y(n_665)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_665),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_666),
.B(n_668),
.Y(n_694)
);

XOR2xp5_ASAP7_75t_L g667 ( 
.A(n_649),
.B(n_621),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_667),
.B(n_672),
.Y(n_691)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_642),
.B(n_625),
.C(n_615),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_658),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_669),
.B(n_670),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_645),
.B(n_622),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_671),
.B(n_673),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_652),
.Y(n_672)
);

XNOR2xp5_ASAP7_75t_L g673 ( 
.A(n_649),
.B(n_648),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_SL g682 ( 
.A1(n_674),
.A2(n_679),
.B1(n_680),
.B2(n_650),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_676),
.B(n_678),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_641),
.A2(n_310),
.B1(n_273),
.B2(n_289),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_652),
.A2(n_356),
.B(n_310),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_654),
.B(n_317),
.C(n_264),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g683 ( 
.A(n_681),
.B(n_659),
.C(n_657),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_683),
.Y(n_699)
);

MAJIxp5_ASAP7_75t_L g684 ( 
.A(n_677),
.B(n_659),
.C(n_640),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_684),
.B(n_685),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_673),
.B(n_655),
.Y(n_685)
);

NAND4xp25_ASAP7_75t_SL g686 ( 
.A(n_675),
.B(n_643),
.C(n_647),
.D(n_651),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_686),
.B(n_689),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_677),
.A2(n_674),
.B(n_644),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_687),
.A2(n_679),
.B(n_681),
.Y(n_700)
);

A2O1A1Ixp33_ASAP7_75t_SL g688 ( 
.A1(n_664),
.A2(n_653),
.B(n_323),
.C(n_314),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_688),
.B(n_323),
.Y(n_703)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_663),
.B(n_317),
.C(n_314),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_695),
.B(n_8),
.Y(n_706)
);

XOR2xp5_ASAP7_75t_L g697 ( 
.A(n_683),
.B(n_667),
.Y(n_697)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_697),
.Y(n_708)
);

XNOR2xp5_ASAP7_75t_L g698 ( 
.A(n_694),
.B(n_668),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_698),
.B(n_701),
.Y(n_711)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_700),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_692),
.A2(n_314),
.B1(n_228),
.B2(n_301),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_702),
.B(n_705),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_703),
.B(n_706),
.Y(n_713)
);

MAJIxp5_ASAP7_75t_L g705 ( 
.A(n_690),
.B(n_323),
.C(n_7),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_684),
.Y(n_707)
);

NOR2x1_ASAP7_75t_L g709 ( 
.A(n_707),
.B(n_696),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_709),
.B(n_688),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_704),
.A2(n_691),
.B(n_693),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_714),
.A2(n_699),
.B(n_697),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_712),
.B(n_707),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_L g719 ( 
.A1(n_715),
.A2(n_717),
.B(n_713),
.Y(n_719)
);

MAJIxp5_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_718),
.C(n_708),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_710),
.A2(n_686),
.B(n_688),
.Y(n_718)
);

AOI322xp5_ASAP7_75t_L g721 ( 
.A1(n_719),
.A2(n_720),
.A3(n_711),
.B1(n_713),
.B2(n_688),
.C1(n_695),
.C2(n_703),
.Y(n_721)
);

OAI21xp5_ASAP7_75t_L g722 ( 
.A1(n_721),
.A2(n_6),
.B(n_7),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_722),
.A2(n_7),
.B(n_8),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_723),
.B(n_8),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_724),
.B(n_8),
.Y(n_725)
);


endmodule