module real_aes_15720_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_1797;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1893;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1872;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_1856;
wire n_658;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1802;
wire n_397;
wire n_1056;
wire n_1083;
wire n_1592;
wire n_1605;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1584;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1842;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1631 ( .A1(n_0), .A2(n_97), .B1(n_1588), .B2(n_1591), .Y(n_1631) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_1), .A2(n_332), .B1(n_464), .B2(n_584), .Y(n_583) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_1), .Y(n_634) );
INVx1_ASAP7_75t_L g1513 ( .A(n_2), .Y(n_1513) );
INVx1_ASAP7_75t_L g843 ( .A(n_3), .Y(n_843) );
AO22x1_ASAP7_75t_L g882 ( .A1(n_3), .A2(n_241), .B1(n_516), .B2(n_771), .Y(n_882) );
INVx1_ASAP7_75t_L g392 ( .A(n_4), .Y(n_392) );
AND2x2_ASAP7_75t_L g445 ( .A(n_4), .B(n_266), .Y(n_445) );
AND2x2_ASAP7_75t_L g506 ( .A(n_4), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g880 ( .A(n_4), .B(n_402), .Y(n_880) );
INVx1_ASAP7_75t_L g855 ( .A(n_5), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_5), .A2(n_131), .B1(n_521), .B2(n_767), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g1438 ( .A1(n_6), .A2(n_46), .B1(n_464), .B2(n_487), .Y(n_1438) );
INVxp67_ASAP7_75t_SL g1463 ( .A(n_6), .Y(n_1463) );
INVx1_ASAP7_75t_L g1822 ( .A(n_7), .Y(n_1822) );
INVx1_ASAP7_75t_L g1162 ( .A(n_8), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_9), .A2(n_208), .B1(n_479), .B2(n_1521), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_9), .A2(n_193), .B1(n_706), .B2(n_1010), .Y(n_1529) );
XOR2x2_ASAP7_75t_L g1328 ( .A(n_10), .B(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1854 ( .A(n_11), .Y(n_1854) );
OAI22xp5_ASAP7_75t_L g1872 ( .A1(n_11), .A2(n_364), .B1(n_559), .B2(n_605), .Y(n_1872) );
OAI22xp5_ASAP7_75t_L g1826 ( .A1(n_12), .A2(n_156), .B1(n_394), .B2(n_1827), .Y(n_1826) );
OAI22xp5_ASAP7_75t_L g1830 ( .A1(n_12), .A2(n_156), .B1(n_1831), .B2(n_1833), .Y(n_1830) );
CKINVDCx5p33_ASAP7_75t_R g1289 ( .A(n_13), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_14), .A2(n_230), .B1(n_413), .B2(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1078 ( .A(n_15), .Y(n_1078) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_16), .A2(n_234), .B1(n_995), .B2(n_996), .Y(n_994) );
INVxp67_ASAP7_75t_SL g1025 ( .A(n_16), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g1550 ( .A1(n_17), .A2(n_323), .B1(n_524), .B2(n_769), .C(n_1551), .Y(n_1550) );
AOI22xp33_ASAP7_75t_SL g1567 ( .A1(n_17), .A2(n_345), .B1(n_470), .B2(n_590), .Y(n_1567) );
INVxp67_ASAP7_75t_SL g1086 ( .A(n_18), .Y(n_1086) );
AND4x1_ASAP7_75t_L g1134 ( .A(n_18), .B(n_1088), .C(n_1091), .D(n_1116), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_19), .A2(n_347), .B1(n_528), .B2(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g740 ( .A(n_19), .Y(n_740) );
INVx2_ASAP7_75t_L g423 ( .A(n_20), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_21), .A2(n_128), .B1(n_473), .B2(n_586), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_21), .A2(n_179), .B1(n_691), .B2(n_763), .Y(n_1313) );
INVx1_ASAP7_75t_L g1038 ( .A(n_22), .Y(n_1038) );
OAI222xp33_ASAP7_75t_L g1062 ( .A1(n_22), .A2(n_182), .B1(n_626), .B2(n_725), .C1(n_1063), .C2(n_1068), .Y(n_1062) );
INVx1_ASAP7_75t_L g1208 ( .A(n_23), .Y(n_1208) );
INVx1_ASAP7_75t_L g966 ( .A(n_24), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g1552 ( .A1(n_25), .A2(n_281), .B1(n_531), .B2(n_537), .Y(n_1552) );
AOI22xp33_ASAP7_75t_L g1569 ( .A1(n_25), .A2(n_278), .B1(n_464), .B2(n_797), .Y(n_1569) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_26), .A2(n_277), .B1(n_594), .B2(n_600), .Y(n_593) );
INVx1_ASAP7_75t_L g618 ( .A(n_26), .Y(n_618) );
INVx1_ASAP7_75t_L g1206 ( .A(n_27), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_27), .A2(n_75), .B1(n_1011), .B2(n_1225), .Y(n_1224) );
AOI22xp33_ASAP7_75t_SL g1801 ( .A1(n_28), .A2(n_176), .B1(n_531), .B2(n_1170), .Y(n_1801) );
AOI22xp33_ASAP7_75t_L g1810 ( .A1(n_28), .A2(n_218), .B1(n_590), .B2(n_850), .Y(n_1810) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_29), .A2(n_171), .B1(n_559), .B2(n_605), .Y(n_1090) );
OAI211xp5_ASAP7_75t_L g1092 ( .A1(n_29), .A2(n_608), .B(n_1093), .C(n_1096), .Y(n_1092) );
INVx1_ASAP7_75t_L g430 ( .A(n_30), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g1307 ( .A1(n_31), .A2(n_222), .B1(n_600), .B2(n_1164), .Y(n_1307) );
INVx1_ASAP7_75t_L g1315 ( .A(n_31), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_32), .A2(n_134), .B1(n_479), .B2(n_586), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_32), .A2(n_306), .B1(n_1011), .B2(n_1225), .Y(n_1498) );
AOI22xp33_ASAP7_75t_SL g1303 ( .A1(n_33), .A2(n_92), .B1(n_466), .B2(n_1298), .Y(n_1303) );
AOI22xp33_ASAP7_75t_SL g1321 ( .A1(n_33), .A2(n_252), .B1(n_1170), .B2(n_1322), .Y(n_1321) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_34), .A2(n_95), .B1(n_706), .B2(n_771), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_34), .A2(n_41), .B1(n_479), .B2(n_1124), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_35), .Y(n_387) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_35), .B(n_385), .Y(n_1582) );
OAI22xp5_ASAP7_75t_SL g933 ( .A1(n_36), .A2(n_307), .B1(n_934), .B2(n_935), .Y(n_933) );
INVxp67_ASAP7_75t_SL g970 ( .A(n_36), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g975 ( .A(n_37), .Y(n_975) );
INVx1_ASAP7_75t_L g1241 ( .A(n_38), .Y(n_1241) );
OAI211xp5_ASAP7_75t_L g1249 ( .A1(n_38), .A2(n_1015), .B(n_1061), .C(n_1250), .Y(n_1249) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_39), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g1556 ( .A1(n_40), .A2(n_345), .B1(n_537), .B2(n_720), .Y(n_1556) );
AOI22xp5_ASAP7_75t_L g1568 ( .A1(n_40), .A2(n_323), .B1(n_590), .B2(n_1045), .Y(n_1568) );
AOI221xp5_ASAP7_75t_L g1113 ( .A1(n_41), .A2(n_355), .B1(n_704), .B2(n_767), .C(n_1114), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1630 ( .A1(n_42), .A2(n_74), .B1(n_1581), .B2(n_1585), .Y(n_1630) );
INVx1_ASAP7_75t_L g1059 ( .A(n_43), .Y(n_1059) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_44), .A2(n_325), .B1(n_767), .B2(n_769), .C(n_1216), .Y(n_1263) );
INVxp67_ASAP7_75t_SL g1270 ( .A(n_44), .Y(n_1270) );
INVx1_ASAP7_75t_L g1246 ( .A(n_45), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_45), .A2(n_224), .B1(n_608), .B2(n_1265), .Y(n_1264) );
AOI221xp5_ASAP7_75t_L g1454 ( .A1(n_46), .A2(n_103), .B1(n_1223), .B2(n_1455), .C(n_1456), .Y(n_1454) );
INVx1_ASAP7_75t_L g723 ( .A(n_47), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_48), .A2(n_298), .B1(n_589), .B2(n_793), .Y(n_991) );
INVx1_ASAP7_75t_L g1018 ( .A(n_48), .Y(n_1018) );
OAI21xp5_ASAP7_75t_L g1560 ( .A1(n_49), .A2(n_657), .B(n_1561), .Y(n_1560) );
NAND5xp2_ASAP7_75t_L g758 ( .A(n_50), .B(n_759), .C(n_789), .D(n_804), .E(n_814), .Y(n_758) );
INVx1_ASAP7_75t_L g823 ( .A(n_50), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_51), .A2(n_155), .B1(n_559), .B2(n_605), .Y(n_604) );
OAI211xp5_ASAP7_75t_SL g607 ( .A1(n_51), .A2(n_608), .B(n_609), .C(n_616), .Y(n_607) );
INVx1_ASAP7_75t_L g722 ( .A(n_52), .Y(n_722) );
INVx1_ASAP7_75t_L g1058 ( .A(n_53), .Y(n_1058) );
XOR2xp5_ASAP7_75t_L g1845 ( .A(n_54), .B(n_1846), .Y(n_1845) );
AOI22xp33_ASAP7_75t_L g1859 ( .A1(n_55), .A2(n_199), .B1(n_691), .B2(n_1860), .Y(n_1859) );
AOI22xp33_ASAP7_75t_SL g1879 ( .A1(n_55), .A2(n_338), .B1(n_464), .B2(n_1122), .Y(n_1879) );
INVxp67_ASAP7_75t_SL g1262 ( .A(n_56), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_56), .A2(n_144), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
INVxp67_ASAP7_75t_L g1287 ( .A(n_57), .Y(n_1287) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_58), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g1793 ( .A1(n_59), .A2(n_218), .B1(n_1312), .B2(n_1794), .Y(n_1793) );
AOI22xp33_ASAP7_75t_L g1804 ( .A1(n_59), .A2(n_176), .B1(n_1519), .B2(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1094 ( .A(n_60), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g1118 ( .A1(n_60), .A2(n_106), .B1(n_594), .B2(n_1119), .Y(n_1118) );
AOI22xp33_ASAP7_75t_SL g1516 ( .A1(n_61), .A2(n_62), .B1(n_464), .B2(n_996), .Y(n_1516) );
INVx1_ASAP7_75t_L g1533 ( .A(n_61), .Y(n_1533) );
AOI221xp5_ASAP7_75t_L g1528 ( .A1(n_62), .A2(n_145), .B1(n_614), .B2(n_1098), .C(n_1217), .Y(n_1528) );
AOI22xp5_ASAP7_75t_L g1606 ( .A1(n_63), .A2(n_122), .B1(n_1581), .B2(n_1585), .Y(n_1606) );
AOI22xp5_ASAP7_75t_L g1596 ( .A1(n_64), .A2(n_271), .B1(n_1581), .B2(n_1585), .Y(n_1596) );
XOR2xp5_ASAP7_75t_L g574 ( .A(n_65), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g983 ( .A(n_66), .Y(n_983) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_67), .A2(n_302), .B1(n_586), .B2(n_589), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_67), .A2(n_270), .B1(n_641), .B2(n_643), .C(n_645), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g1439 ( .A1(n_68), .A2(n_279), .B1(n_479), .B2(n_1440), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_68), .A2(n_149), .B1(n_530), .B2(n_537), .Y(n_1457) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_69), .A2(n_183), .B1(n_521), .B2(n_767), .C(n_769), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_69), .A2(n_248), .B1(n_590), .B2(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g494 ( .A(n_70), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_71), .A2(n_248), .B1(n_720), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_71), .A2(n_183), .B1(n_590), .B2(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g1340 ( .A(n_72), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g1097 ( .A1(n_73), .A2(n_354), .B1(n_614), .B2(n_1098), .C(n_1100), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g1128 ( .A1(n_73), .A2(n_315), .B1(n_1043), .B2(n_1129), .Y(n_1128) );
AOI22xp5_ASAP7_75t_L g1540 ( .A1(n_74), .A2(n_1541), .B1(n_1542), .B2(n_1571), .Y(n_1540) );
INVxp67_ASAP7_75t_SL g1571 ( .A(n_74), .Y(n_1571) );
INVx1_ASAP7_75t_L g1195 ( .A(n_75), .Y(n_1195) );
INVx1_ASAP7_75t_L g1815 ( .A(n_76), .Y(n_1815) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_77), .A2(n_303), .B1(n_464), .B2(n_466), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_77), .A2(n_322), .B1(n_530), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_78), .A2(n_187), .B1(n_745), .B2(n_987), .Y(n_986) );
INVxp67_ASAP7_75t_SL g1024 ( .A(n_78), .Y(n_1024) );
INVx1_ASAP7_75t_L g1548 ( .A(n_79), .Y(n_1548) );
OAI22xp5_ASAP7_75t_L g1368 ( .A1(n_80), .A2(n_264), .B1(n_1369), .B2(n_1373), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_80), .A2(n_264), .B1(n_1407), .B2(n_1409), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_81), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_82), .A2(n_245), .B1(n_487), .B2(n_995), .Y(n_1153) );
AOI22xp33_ASAP7_75t_SL g1180 ( .A1(n_82), .A2(n_304), .B1(n_528), .B2(n_706), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1618 ( .A1(n_83), .A2(n_260), .B1(n_1581), .B2(n_1585), .Y(n_1618) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_84), .A2(n_103), .B1(n_487), .B2(n_1445), .Y(n_1444) );
INVxp67_ASAP7_75t_SL g1464 ( .A(n_84), .Y(n_1464) );
INVx1_ASAP7_75t_L g1549 ( .A(n_85), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_86), .B(n_432), .Y(n_1244) );
OAI221xp5_ASAP7_75t_L g1256 ( .A1(n_87), .A2(n_221), .B1(n_1257), .B2(n_1258), .C(n_1259), .Y(n_1256) );
OAI322xp33_ASAP7_75t_L g1268 ( .A1(n_87), .A2(n_600), .A3(n_951), .B1(n_1210), .B2(n_1269), .C1(n_1272), .C2(n_1276), .Y(n_1268) );
AOI22xp5_ASAP7_75t_L g1600 ( .A1(n_88), .A2(n_265), .B1(n_1588), .B2(n_1591), .Y(n_1600) );
AOI22xp33_ASAP7_75t_SL g1152 ( .A1(n_89), .A2(n_237), .B1(n_1149), .B2(n_1151), .Y(n_1152) );
INVx1_ASAP7_75t_L g1176 ( .A(n_89), .Y(n_1176) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_90), .A2(n_559), .B(n_568), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g938 ( .A1(n_91), .A2(n_167), .B1(n_516), .B2(n_939), .Y(n_938) );
INVxp67_ASAP7_75t_SL g962 ( .A(n_91), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g1311 ( .A1(n_92), .A2(n_337), .B1(n_525), .B2(n_767), .C(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1028 ( .A(n_93), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g1601 ( .A1(n_93), .A2(n_111), .B1(n_1581), .B2(n_1602), .Y(n_1601) );
AO22x1_ASAP7_75t_L g1624 ( .A1(n_94), .A2(n_273), .B1(n_1588), .B2(n_1591), .Y(n_1624) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_95), .A2(n_355), .B1(n_479), .B2(n_1124), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_96), .A2(n_288), .B1(n_464), .B2(n_672), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_96), .A2(n_284), .B1(n_524), .B2(n_525), .C(n_613), .Y(n_689) );
INVx1_ASAP7_75t_L g670 ( .A(n_98), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_98), .A2(n_313), .B1(n_531), .B2(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g1339 ( .A(n_99), .Y(n_1339) );
AOI22xp33_ASAP7_75t_SL g1048 ( .A1(n_100), .A2(n_342), .B1(n_464), .B2(n_672), .Y(n_1048) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_100), .Y(n_1053) );
INVx1_ASAP7_75t_L g1205 ( .A(n_101), .Y(n_1205) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_101), .A2(n_239), .B1(n_704), .B2(n_1216), .C(n_1217), .Y(n_1215) );
AOI22xp33_ASAP7_75t_SL g1802 ( .A1(n_102), .A2(n_372), .B1(n_1312), .B2(n_1794), .Y(n_1802) );
AOI22xp33_ASAP7_75t_L g1811 ( .A1(n_102), .A2(n_104), .B1(n_1043), .B2(n_1807), .Y(n_1811) );
AOI22xp33_ASAP7_75t_L g1796 ( .A1(n_104), .A2(n_339), .B1(n_531), .B2(n_1797), .Y(n_1796) );
XNOR2xp5_ASAP7_75t_L g710 ( .A(n_105), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g1095 ( .A(n_106), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_107), .A2(n_333), .B1(n_468), .B2(n_473), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g538 ( .A1(n_107), .A2(n_357), .B1(n_539), .B2(n_543), .C(n_547), .Y(n_538) );
OAI211xp5_ASAP7_75t_L g776 ( .A1(n_108), .A2(n_777), .B(n_778), .C(n_779), .Y(n_776) );
INVx1_ASAP7_75t_L g819 ( .A(n_108), .Y(n_819) );
INVx1_ASAP7_75t_L g1511 ( .A(n_109), .Y(n_1511) );
OAI221xp5_ASAP7_75t_L g1531 ( .A1(n_109), .A2(n_147), .B1(n_622), .B2(n_1258), .C(n_1532), .Y(n_1531) );
INVx1_ASAP7_75t_L g1260 ( .A(n_110), .Y(n_1260) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_112), .A2(n_246), .B1(n_516), .B2(n_693), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_112), .A2(n_272), .B1(n_487), .B2(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g1353 ( .A(n_113), .Y(n_1353) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_114), .A2(n_524), .B(n_547), .Y(n_731) );
INVx1_ASAP7_75t_L g739 ( .A(n_114), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_115), .A2(n_322), .B1(n_464), .B2(n_487), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_115), .A2(n_303), .B1(n_520), .B2(n_523), .C(n_525), .Y(n_519) );
INVx1_ASAP7_75t_L g655 ( .A(n_116), .Y(n_655) );
INVx1_ASAP7_75t_L g925 ( .A(n_117), .Y(n_925) );
INVx1_ASAP7_75t_L g1514 ( .A(n_118), .Y(n_1514) );
OAI221xp5_ASAP7_75t_L g1103 ( .A1(n_119), .A2(n_286), .B1(n_622), .B2(n_625), .C(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1133 ( .A(n_119), .Y(n_1133) );
INVx1_ASAP7_75t_L g385 ( .A(n_120), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_121), .A2(n_269), .B1(n_525), .B2(n_716), .C(n_717), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_121), .A2(n_190), .B1(n_453), .B2(n_464), .Y(n_741) );
AO221x2_ASAP7_75t_L g1691 ( .A1(n_123), .A2(n_351), .B1(n_1588), .B2(n_1591), .C(n_1692), .Y(n_1691) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_124), .A2(n_301), .B1(n_464), .B2(n_466), .Y(n_592) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_124), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_125), .A2(n_196), .B1(n_793), .B2(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1022 ( .A(n_125), .Y(n_1022) );
OAI22xp33_ASAP7_75t_L g1192 ( .A1(n_126), .A2(n_320), .B1(n_594), .B2(n_1119), .Y(n_1192) );
INVx1_ASAP7_75t_L g1227 ( .A(n_126), .Y(n_1227) );
OAI222xp33_ASAP7_75t_L g866 ( .A1(n_127), .A2(n_349), .B1(n_867), .B2(n_869), .C1(n_871), .C2(n_873), .Y(n_866) );
INVx1_ASAP7_75t_L g886 ( .A(n_127), .Y(n_886) );
AOI21xp33_ASAP7_75t_L g1320 ( .A1(n_128), .A2(n_769), .B(n_773), .Y(n_1320) );
INVx1_ASAP7_75t_L g1436 ( .A(n_129), .Y(n_1436) );
OAI221xp5_ASAP7_75t_L g1461 ( .A1(n_129), .A2(n_130), .B1(n_622), .B2(n_1258), .C(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1435 ( .A(n_130), .Y(n_1435) );
INVx1_ASAP7_75t_L g851 ( .A(n_131), .Y(n_851) );
OAI211xp5_ASAP7_75t_L g927 ( .A1(n_132), .A2(n_928), .B(n_929), .C(n_930), .Y(n_927) );
INVxp33_ASAP7_75t_SL g948 ( .A(n_132), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_133), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g1493 ( .A1(n_134), .A2(n_251), .B1(n_704), .B2(n_1216), .C(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1197 ( .A(n_135), .Y(n_1197) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_135), .A2(n_295), .B1(n_1216), .B2(n_1222), .C(n_1223), .Y(n_1221) );
INVxp67_ASAP7_75t_SL g1863 ( .A(n_136), .Y(n_1863) );
AOI22xp33_ASAP7_75t_L g1880 ( .A1(n_136), .A2(n_275), .B1(n_1046), .B2(n_1805), .Y(n_1880) );
INVx1_ASAP7_75t_L g1554 ( .A(n_137), .Y(n_1554) );
INVx1_ASAP7_75t_L g665 ( .A(n_138), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g703 ( .A1(n_138), .A2(n_524), .B(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_139), .A2(n_178), .B1(n_605), .B2(n_657), .Y(n_656) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_139), .A2(n_687), .B(n_688), .C(n_694), .Y(n_686) );
INVx1_ASAP7_75t_L g979 ( .A(n_140), .Y(n_979) );
OAI222xp33_ASAP7_75t_L g1014 ( .A1(n_140), .A2(n_219), .B1(n_625), .B2(n_1015), .C1(n_1016), .C2(n_1023), .Y(n_1014) );
INVx1_ASAP7_75t_L g1853 ( .A(n_141), .Y(n_1853) );
OAI22xp33_ASAP7_75t_L g1883 ( .A1(n_141), .A2(n_189), .B1(n_1119), .B2(n_1164), .Y(n_1883) );
XOR2x2_ASAP7_75t_L g1472 ( .A(n_142), .B(n_1473), .Y(n_1472) );
INVxp67_ASAP7_75t_SL g1857 ( .A(n_143), .Y(n_1857) );
AOI22xp33_ASAP7_75t_SL g1881 ( .A1(n_143), .A2(n_210), .B1(n_479), .B2(n_1149), .Y(n_1881) );
AOI221xp5_ASAP7_75t_L g1255 ( .A1(n_144), .A2(n_232), .B1(n_520), .B2(n_525), .C(n_767), .Y(n_1255) );
AOI22xp33_ASAP7_75t_SL g1523 ( .A1(n_145), .A2(n_150), .B1(n_466), .B2(n_1524), .Y(n_1523) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_146), .A2(n_278), .B1(n_545), .B2(n_716), .C(n_774), .Y(n_1555) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_146), .A2(n_281), .B1(n_453), .B2(n_464), .Y(n_1566) );
INVx1_ASAP7_75t_L g1510 ( .A(n_147), .Y(n_1510) );
AO22x1_ASAP7_75t_L g1587 ( .A1(n_148), .A2(n_358), .B1(n_1588), .B2(n_1591), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_149), .A2(n_186), .B1(n_479), .B2(n_1440), .Y(n_1442) );
INVxp67_ASAP7_75t_SL g1534 ( .A(n_150), .Y(n_1534) );
INVx1_ASAP7_75t_L g1142 ( .A(n_151), .Y(n_1142) );
OAI221xp5_ASAP7_75t_L g1174 ( .A1(n_151), .A2(n_152), .B1(n_626), .B2(n_725), .C(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1143 ( .A(n_152), .Y(n_1143) );
AOI22xp33_ASAP7_75t_SL g1480 ( .A1(n_153), .A2(n_180), .B1(n_466), .B2(n_1445), .Y(n_1480) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_153), .A2(n_204), .B1(n_525), .B2(n_539), .C(n_643), .Y(n_1499) );
OAI22xp33_ASAP7_75t_L g1484 ( .A1(n_154), .A2(n_316), .B1(n_600), .B2(n_1164), .Y(n_1484) );
INVx1_ASAP7_75t_L g1501 ( .A(n_154), .Y(n_1501) );
OAI22xp33_ASAP7_75t_L g1447 ( .A1(n_157), .A2(n_297), .B1(n_594), .B2(n_600), .Y(n_1447) );
INVx1_ASAP7_75t_L g1460 ( .A(n_157), .Y(n_1460) );
INVx1_ASAP7_75t_L g1544 ( .A(n_158), .Y(n_1544) );
INVx1_ASAP7_75t_L g1001 ( .A(n_159), .Y(n_1001) );
INVx1_ASAP7_75t_L g1292 ( .A(n_160), .Y(n_1292) );
OAI221xp5_ASAP7_75t_SL g1317 ( .A1(n_160), .A2(n_276), .B1(n_622), .B2(n_625), .C(n_1318), .Y(n_1317) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_161), .A2(n_361), .B1(n_626), .B2(n_725), .C(n_726), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g747 ( .A1(n_161), .A2(n_361), .B1(n_491), .B2(n_683), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g1389 ( .A1(n_162), .A2(n_169), .B1(n_1390), .B2(n_1393), .Y(n_1389) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_162), .A2(n_169), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
INVx1_ASAP7_75t_L g813 ( .A(n_163), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g1486 ( .A(n_164), .Y(n_1486) );
INVx1_ASAP7_75t_L g1821 ( .A(n_165), .Y(n_1821) );
INVx1_ASAP7_75t_L g1380 ( .A(n_166), .Y(n_1380) );
INVx1_ASAP7_75t_L g955 ( .A(n_167), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_168), .Y(n_603) );
AO22x1_ASAP7_75t_L g1622 ( .A1(n_170), .A2(n_360), .B1(n_1581), .B2(n_1623), .Y(n_1622) );
CKINVDCx16_ASAP7_75t_R g1693 ( .A(n_172), .Y(n_1693) );
INVx1_ASAP7_75t_L g1345 ( .A(n_173), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_174), .A2(n_359), .B1(n_559), .B2(n_605), .Y(n_1487) );
OAI22xp5_ASAP7_75t_L g1507 ( .A1(n_175), .A2(n_305), .B1(n_559), .B2(n_605), .Y(n_1507) );
CKINVDCx5p33_ASAP7_75t_R g932 ( .A(n_177), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_179), .A2(n_327), .B1(n_473), .B2(n_1301), .Y(n_1300) );
INVxp67_ASAP7_75t_SL g1491 ( .A(n_180), .Y(n_1491) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_181), .A2(n_202), .B1(n_559), .B2(n_605), .Y(n_1450) );
OAI211xp5_ASAP7_75t_L g1452 ( .A1(n_181), .A2(n_687), .B(n_1453), .C(n_1458), .Y(n_1452) );
INVx1_ASAP7_75t_L g1037 ( .A(n_182), .Y(n_1037) );
INVx1_ASAP7_75t_L g845 ( .A(n_184), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_184), .A2(n_280), .B1(n_720), .B2(n_771), .Y(n_903) );
INVx1_ASAP7_75t_L g573 ( .A(n_185), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g1465 ( .A1(n_186), .A2(n_279), .B1(n_704), .B2(n_1216), .C(n_1466), .Y(n_1465) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_187), .A2(n_234), .B1(n_614), .B2(n_641), .C(n_643), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_188), .Y(n_931) );
INVx1_ASAP7_75t_L g1851 ( .A(n_189), .Y(n_1851) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_190), .A2(n_331), .B1(n_516), .B2(n_537), .Y(n_732) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_191), .A2(n_687), .B(n_714), .C(n_721), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_191), .A2(n_353), .B1(n_605), .B2(n_657), .Y(n_750) );
INVx1_ASAP7_75t_L g942 ( .A(n_192), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g1517 ( .A1(n_193), .A2(n_289), .B1(n_1518), .B2(n_1519), .Y(n_1517) );
AOI22xp33_ASAP7_75t_SL g1148 ( .A1(n_194), .A2(n_310), .B1(n_1149), .B2(n_1151), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_194), .A2(n_237), .B1(n_531), .B2(n_1170), .Y(n_1169) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_195), .A2(n_761), .B(n_764), .C(n_775), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_195), .B(n_413), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_196), .A2(n_298), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
INVx1_ASAP7_75t_L g1478 ( .A(n_197), .Y(n_1478) );
OAI221xp5_ASAP7_75t_L g1489 ( .A1(n_197), .A2(n_335), .B1(n_725), .B2(n_1258), .C(n_1490), .Y(n_1489) );
INVx2_ASAP7_75t_L g1584 ( .A(n_198), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_198), .B(n_314), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_198), .B(n_1590), .Y(n_1592) );
AOI22xp33_ASAP7_75t_SL g1882 ( .A1(n_199), .A2(n_370), .B1(n_464), .B2(n_1043), .Y(n_1882) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_200), .A2(n_366), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
INVx1_ASAP7_75t_L g1066 ( .A(n_200), .Y(n_1066) );
CKINVDCx5p33_ASAP7_75t_R g1267 ( .A(n_201), .Y(n_1267) );
INVx1_ASAP7_75t_L g696 ( .A(n_203), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g1483 ( .A1(n_204), .A2(n_309), .B1(n_487), .B2(n_957), .Y(n_1483) );
INVx1_ASAP7_75t_L g508 ( .A(n_205), .Y(n_508) );
XOR2x2_ASAP7_75t_L g1430 ( .A(n_206), .B(n_1431), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_207), .A2(n_357), .B1(n_468), .B2(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_207), .A2(n_333), .B1(n_528), .B2(n_530), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g1535 ( .A1(n_208), .A2(n_289), .B1(n_767), .B2(n_769), .C(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g1306 ( .A(n_209), .Y(n_1306) );
INVxp67_ASAP7_75t_SL g1865 ( .A(n_210), .Y(n_1865) );
INVx1_ASAP7_75t_L g914 ( .A(n_211), .Y(n_914) );
NOR2xp33_ASAP7_75t_L g1867 ( .A(n_212), .B(n_725), .Y(n_1867) );
INVx1_ASAP7_75t_L g1877 ( .A(n_212), .Y(n_1877) );
INVx1_ASAP7_75t_L g1000 ( .A(n_213), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_214), .A2(n_294), .B1(n_693), .B2(n_720), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_214), .A2(n_312), .B1(n_464), .B2(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_215), .A2(n_284), .B1(n_464), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_215), .A2(n_288), .B1(n_537), .B2(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g1077 ( .A(n_216), .Y(n_1077) );
INVx1_ASAP7_75t_L g1201 ( .A(n_217), .Y(n_1201) );
INVx1_ASAP7_75t_L g980 ( .A(n_219), .Y(n_980) );
OAI211xp5_ASAP7_75t_L g1376 ( .A1(n_220), .A2(n_1364), .B(n_1377), .C(n_1379), .Y(n_1376) );
INVx1_ASAP7_75t_L g1422 ( .A(n_220), .Y(n_1422) );
INVx1_ASAP7_75t_L g1240 ( .A(n_221), .Y(n_1240) );
INVx1_ASAP7_75t_L g1316 ( .A(n_222), .Y(n_1316) );
CKINVDCx5p33_ASAP7_75t_R g848 ( .A(n_223), .Y(n_848) );
INVx1_ASAP7_75t_L g1243 ( .A(n_224), .Y(n_1243) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_225), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_226), .A2(n_369), .B1(n_600), .B2(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1172 ( .A(n_226), .Y(n_1172) );
INVx1_ASAP7_75t_L g1282 ( .A(n_227), .Y(n_1282) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_228), .Y(n_783) );
INVx2_ASAP7_75t_L g425 ( .A(n_229), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_229), .B(n_423), .Y(n_440) );
INVx1_ASAP7_75t_L g485 ( .A(n_229), .Y(n_485) );
OAI211xp5_ASAP7_75t_L g1219 ( .A1(n_230), .A2(n_687), .B(n_1220), .C(n_1226), .Y(n_1219) );
INVx1_ASAP7_75t_L g861 ( .A(n_231), .Y(n_861) );
NAND2xp33_ASAP7_75t_SL g904 ( .A(n_231), .B(n_521), .Y(n_904) );
INVx1_ASAP7_75t_L g1275 ( .A(n_232), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_233), .A2(n_334), .B1(n_676), .B2(n_990), .Y(n_1047) );
INVx1_ASAP7_75t_L g1064 ( .A(n_233), .Y(n_1064) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_235), .A2(n_262), .B1(n_464), .B2(n_1043), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g1069 ( .A(n_235), .Y(n_1069) );
INVx1_ASAP7_75t_L g1352 ( .A(n_236), .Y(n_1352) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_238), .A2(n_321), .B1(n_777), .B2(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g817 ( .A(n_238), .Y(n_817) );
INVx1_ASAP7_75t_L g1203 ( .A(n_239), .Y(n_1203) );
INVx1_ASAP7_75t_L g1254 ( .A(n_240), .Y(n_1254) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_241), .A2(n_800), .B(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g908 ( .A(n_242), .Y(n_908) );
OAI21xp5_ASAP7_75t_L g1074 ( .A1(n_243), .A2(n_657), .B(n_1075), .Y(n_1074) );
BUFx3_ASAP7_75t_L g417 ( .A(n_244), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_245), .A2(n_256), .B1(n_524), .B2(n_525), .C(n_613), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_246), .A2(n_290), .B1(n_487), .B2(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1619 ( .A1(n_247), .A2(n_253), .B1(n_1588), .B2(n_1591), .Y(n_1619) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_249), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_250), .A2(n_257), .B1(n_491), .B2(n_1190), .Y(n_1189) );
OAI221xp5_ASAP7_75t_L g1212 ( .A1(n_250), .A2(n_257), .B1(n_622), .B2(n_625), .C(n_1213), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_251), .A2(n_306), .B1(n_479), .B2(n_850), .Y(n_1482) );
AOI22xp33_ASAP7_75t_SL g1297 ( .A1(n_252), .A2(n_337), .B1(n_996), .B2(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g834 ( .A(n_254), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_254), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1820 ( .A(n_255), .Y(n_1820) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_256), .A2(n_304), .B1(n_487), .B2(n_987), .Y(n_1147) );
AOI21xp33_ASAP7_75t_L g943 ( .A1(n_258), .A2(n_524), .B(n_769), .Y(n_943) );
INVx1_ASAP7_75t_L g953 ( .A(n_258), .Y(n_953) );
INVx1_ASAP7_75t_L g502 ( .A(n_259), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_260), .A2(n_1186), .B1(n_1187), .B2(n_1234), .Y(n_1185) );
INVx1_ASAP7_75t_L g1234 ( .A(n_260), .Y(n_1234) );
XOR2x2_ASAP7_75t_L g920 ( .A(n_261), .B(n_921), .Y(n_920) );
AOI21xp33_ASAP7_75t_L g1055 ( .A1(n_262), .A2(n_644), .B(n_774), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_263), .B(n_1138), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1157 ( .A1(n_263), .A2(n_1158), .B1(n_1159), .B2(n_1181), .Y(n_1157) );
INVx1_ASAP7_75t_L g1183 ( .A(n_263), .Y(n_1183) );
BUFx3_ASAP7_75t_L g402 ( .A(n_266), .Y(n_402) );
INVx1_ASAP7_75t_L g507 ( .A(n_266), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g1695 ( .A(n_267), .Y(n_1695) );
AOI22xp5_ASAP7_75t_L g1595 ( .A1(n_268), .A2(n_283), .B1(n_1588), .B2(n_1591), .Y(n_1595) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_269), .A2(n_331), .B1(n_464), .B2(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_270), .A2(n_324), .B1(n_586), .B2(n_589), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g937 ( .A(n_272), .B(n_524), .Y(n_937) );
INVxp67_ASAP7_75t_SL g1295 ( .A(n_274), .Y(n_1295) );
OAI211xp5_ASAP7_75t_SL g1309 ( .A1(n_274), .A2(n_608), .B(n_1310), .C(n_1314), .Y(n_1309) );
AOI21xp5_ASAP7_75t_L g1861 ( .A1(n_275), .A2(n_769), .B(n_1217), .Y(n_1861) );
INVx1_ASAP7_75t_L g1293 ( .A(n_276), .Y(n_1293) );
INVx1_ASAP7_75t_L g617 ( .A(n_277), .Y(n_617) );
INVx1_ASAP7_75t_L g857 ( .A(n_280), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g1156 ( .A(n_282), .Y(n_1156) );
INVx1_ASAP7_75t_L g1251 ( .A(n_285), .Y(n_1251) );
INVx1_ASAP7_75t_L g1131 ( .A(n_286), .Y(n_1131) );
INVx1_ASAP7_75t_L g695 ( .A(n_287), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g940 ( .A(n_290), .B(n_520), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g1605 ( .A1(n_291), .A2(n_363), .B1(n_1588), .B2(n_1591), .Y(n_1605) );
XOR2x2_ASAP7_75t_L g1789 ( .A(n_291), .B(n_1790), .Y(n_1789) );
AOI22xp33_ASAP7_75t_L g1843 ( .A1(n_291), .A2(n_1844), .B1(n_1885), .B2(n_1890), .Y(n_1843) );
AO22x1_ASAP7_75t_L g1580 ( .A1(n_292), .A2(n_299), .B1(n_1581), .B2(n_1585), .Y(n_1580) );
INVx1_ASAP7_75t_L g1817 ( .A(n_293), .Y(n_1817) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_294), .A2(n_374), .B1(n_464), .B2(n_672), .Y(n_791) );
INVx1_ASAP7_75t_L g1209 ( .A(n_295), .Y(n_1209) );
INVx1_ASAP7_75t_L g420 ( .A(n_296), .Y(n_420) );
INVx1_ASAP7_75t_L g437 ( .A(n_296), .Y(n_437) );
INVx1_ASAP7_75t_L g1459 ( .A(n_297), .Y(n_1459) );
CKINVDCx5p33_ASAP7_75t_R g1506 ( .A(n_300), .Y(n_1506) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_301), .A2(n_332), .B1(n_523), .B2(n_611), .C(n_614), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_302), .A2(n_324), .B1(n_528), .B2(n_530), .Y(n_615) );
OAI211xp5_ASAP7_75t_L g1526 ( .A1(n_305), .A2(n_687), .B(n_1527), .C(n_1530), .Y(n_1526) );
OAI21xp33_ASAP7_75t_L g946 ( .A1(n_307), .A2(n_806), .B(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1040 ( .A(n_308), .Y(n_1040) );
INVxp67_ASAP7_75t_SL g1492 ( .A(n_309), .Y(n_1492) );
AOI21xp33_ASAP7_75t_L g1177 ( .A1(n_310), .A2(n_704), .B(n_1178), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_311), .Y(n_832) );
AOI221xp5_ASAP7_75t_SL g772 ( .A1(n_312), .A2(n_374), .B1(n_521), .B2(n_773), .C(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g680 ( .A(n_313), .Y(n_680) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_314), .B(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g1590 ( .A(n_314), .Y(n_1590) );
INVxp67_ASAP7_75t_SL g1112 ( .A(n_315), .Y(n_1112) );
INVx1_ASAP7_75t_L g1502 ( .A(n_316), .Y(n_1502) );
INVx1_ASAP7_75t_L g1385 ( .A(n_317), .Y(n_1385) );
OAI211xp5_ASAP7_75t_L g1415 ( .A1(n_317), .A2(n_1336), .B(n_1416), .C(n_1419), .Y(n_1415) );
OAI211xp5_ASAP7_75t_SL g1855 ( .A1(n_318), .A2(n_1258), .B(n_1856), .C(n_1862), .Y(n_1855) );
INVx1_ASAP7_75t_L g1876 ( .A(n_318), .Y(n_1876) );
INVx1_ASAP7_75t_L g1559 ( .A(n_319), .Y(n_1559) );
INVx1_ASAP7_75t_L g1228 ( .A(n_320), .Y(n_1228) );
INVx1_ASAP7_75t_L g803 ( .A(n_321), .Y(n_803) );
INVxp67_ASAP7_75t_SL g1277 ( .A(n_325), .Y(n_1277) );
INVx1_ASAP7_75t_L g1333 ( .A(n_326), .Y(n_1333) );
INVx1_ASAP7_75t_L g1319 ( .A(n_327), .Y(n_1319) );
INVx1_ASAP7_75t_L g1558 ( .A(n_328), .Y(n_1558) );
INVxp67_ASAP7_75t_SL g1145 ( .A(n_329), .Y(n_1145) );
OAI211xp5_ASAP7_75t_L g1166 ( .A1(n_329), .A2(n_687), .B(n_1167), .C(n_1171), .Y(n_1166) );
CKINVDCx16_ASAP7_75t_R g868 ( .A(n_330), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g1056 ( .A1(n_334), .A2(n_366), .B1(n_531), .B2(n_939), .Y(n_1056) );
INVx1_ASAP7_75t_L g1477 ( .A(n_335), .Y(n_1477) );
OAI21xp33_ASAP7_75t_L g998 ( .A1(n_336), .A2(n_559), .B(n_999), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1866 ( .A1(n_338), .A2(n_370), .B1(n_525), .B2(n_1100), .C(n_1312), .Y(n_1866) );
AOI22xp33_ASAP7_75t_SL g1806 ( .A1(n_339), .A2(n_372), .B1(n_1043), .B2(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g1344 ( .A(n_340), .Y(n_1344) );
INVx1_ASAP7_75t_L g1334 ( .A(n_341), .Y(n_1334) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_342), .Y(n_1072) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_343), .Y(n_449) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_344), .Y(n_1108) );
AOI22xp33_ASAP7_75t_SL g1121 ( .A1(n_344), .A2(n_354), .B1(n_957), .B2(n_1122), .Y(n_1121) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_346), .Y(n_398) );
INVx1_ASAP7_75t_L g743 ( .A(n_347), .Y(n_743) );
INVx1_ASAP7_75t_L g1871 ( .A(n_348), .Y(n_1871) );
NOR2xp33_ASAP7_75t_R g893 ( .A(n_349), .B(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g828 ( .A(n_350), .Y(n_828) );
INVx1_ASAP7_75t_L g579 ( .A(n_352), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g621 ( .A1(n_352), .A2(n_375), .B1(n_622), .B2(n_625), .C(n_630), .Y(n_621) );
INVx1_ASAP7_75t_L g749 ( .A(n_356), .Y(n_749) );
OAI211xp5_ASAP7_75t_L g1496 ( .A1(n_359), .A2(n_687), .B(n_1497), .C(n_1500), .Y(n_1496) );
XOR2x2_ASAP7_75t_L g1503 ( .A(n_360), .B(n_1504), .Y(n_1503) );
INVx1_ASAP7_75t_L g429 ( .A(n_362), .Y(n_429) );
INVx1_ASAP7_75t_L g443 ( .A(n_362), .Y(n_443) );
INVx2_ASAP7_75t_L g462 ( .A(n_362), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g1449 ( .A(n_365), .Y(n_1449) );
CKINVDCx5p33_ASAP7_75t_R g1231 ( .A(n_367), .Y(n_1231) );
OAI22xp33_ASAP7_75t_SL g682 ( .A1(n_368), .A2(n_373), .B1(n_491), .B2(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g697 ( .A1(n_368), .A2(n_373), .B1(n_622), .B2(n_626), .C(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g1173 ( .A(n_369), .Y(n_1173) );
XNOR2xp5_ASAP7_75t_L g652 ( .A(n_371), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g581 ( .A(n_375), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_403), .B(n_1572), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx4f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_388), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g1842 ( .A(n_382), .B(n_391), .Y(n_1842) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1889 ( .A(n_384), .B(n_387), .Y(n_1889) );
INVx1_ASAP7_75t_L g1893 ( .A(n_384), .Y(n_1893) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g1896 ( .A(n_387), .B(n_1893), .Y(n_1896) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g1427 ( .A(n_391), .B(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g526 ( .A(n_392), .B(n_402), .Y(n_526) );
AND2x4_ASAP7_75t_L g548 ( .A(n_392), .B(n_401), .Y(n_548) );
INVx1_ASAP7_75t_L g1402 ( .A(n_393), .Y(n_1402) );
AND2x4_ASAP7_75t_SL g1841 ( .A(n_393), .B(n_1842), .Y(n_1841) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x6_ASAP7_75t_L g394 ( .A(n_395), .B(n_400), .Y(n_394) );
INVxp67_ASAP7_75t_L g1071 ( .A(n_395), .Y(n_1071) );
OR2x6_ASAP7_75t_L g1408 ( .A(n_395), .B(n_1405), .Y(n_1408) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx4f_ASAP7_75t_L g633 ( .A(n_396), .Y(n_633) );
INVx3_ASAP7_75t_L g1107 ( .A(n_396), .Y(n_1107) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx2_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
AND2x2_ASAP7_75t_L g512 ( .A(n_398), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g518 ( .A(n_398), .Y(n_518) );
AND2x2_ASAP7_75t_L g522 ( .A(n_398), .B(n_399), .Y(n_522) );
INVx1_ASAP7_75t_L g563 ( .A(n_398), .Y(n_563) );
NAND2x1_ASAP7_75t_L g702 ( .A(n_398), .B(n_399), .Y(n_702) );
INVx1_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
INVx2_ASAP7_75t_L g513 ( .A(n_399), .Y(n_513) );
AND2x2_ASAP7_75t_L g517 ( .A(n_399), .B(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g553 ( .A(n_399), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_399), .B(n_518), .Y(n_638) );
OR2x2_ASAP7_75t_L g902 ( .A(n_399), .B(n_447), .Y(n_902) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g1418 ( .A(n_401), .Y(n_1418) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g1414 ( .A(n_402), .Y(n_1414) );
AND2x4_ASAP7_75t_L g1425 ( .A(n_402), .B(n_562), .Y(n_1425) );
XNOR2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_1080), .Y(n_403) );
AO22x2_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_1032), .B2(n_1079), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_753), .B1(n_754), .B2(n_1031), .Y(n_406) );
INVx1_ASAP7_75t_L g1031 ( .A(n_407), .Y(n_1031) );
XNOR2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_650), .Y(n_407) );
XOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_574), .Y(n_408) );
XNOR2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_573), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_499), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_430), .B1(n_431), .B2(n_449), .C(n_450), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_412), .B(n_1243), .Y(n_1242) );
AOI211xp5_ASAP7_75t_L g1562 ( .A1(n_412), .A2(n_452), .B(n_1554), .C(n_1563), .Y(n_1562) );
INVx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx5_ASAP7_75t_L g971 ( .A(n_413), .Y(n_971) );
OR2x6_ASAP7_75t_L g413 ( .A(n_414), .B(n_426), .Y(n_413) );
OR2x2_ASAP7_75t_L g605 ( .A(n_414), .B(n_426), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_415), .B(n_421), .Y(n_414) );
INVx8_ASAP7_75t_L g465 ( .A(n_415), .Y(n_465) );
BUFx3_ASAP7_75t_L g863 ( .A(n_415), .Y(n_863) );
BUFx3_ASAP7_75t_L g957 ( .A(n_415), .Y(n_957) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_415), .Y(n_964) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
AND2x4_ASAP7_75t_L g471 ( .A(n_416), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_417), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g454 ( .A(n_417), .B(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_417), .Y(n_476) );
OR2x2_ASAP7_75t_L g597 ( .A(n_417), .B(n_419), .Y(n_597) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g472 ( .A(n_420), .Y(n_472) );
AND2x4_ASAP7_75t_L g456 ( .A(n_421), .B(n_442), .Y(n_456) );
INVx1_ASAP7_75t_L g865 ( .A(n_421), .Y(n_865) );
AND2x6_ASAP7_75t_L g872 ( .A(n_421), .B(n_492), .Y(n_872) );
AND2x2_ASAP7_75t_L g874 ( .A(n_421), .B(n_498), .Y(n_874) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
NAND3x1_ASAP7_75t_L g483 ( .A(n_422), .B(n_484), .C(n_485), .Y(n_483) );
NAND2x1p5_ASAP7_75t_L g800 ( .A(n_422), .B(n_485), .Y(n_800) );
INVx1_ASAP7_75t_L g1372 ( .A(n_422), .Y(n_1372) );
OR2x6_ASAP7_75t_L g1375 ( .A(n_422), .B(n_669), .Y(n_1375) );
AND2x4_ASAP7_75t_L g1378 ( .A(n_422), .B(n_454), .Y(n_1378) );
OR2x4_ASAP7_75t_L g1392 ( .A(n_422), .B(n_597), .Y(n_1392) );
INVx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g460 ( .A(n_423), .Y(n_460) );
NAND2xp33_ASAP7_75t_SL g663 ( .A(n_423), .B(n_425), .Y(n_663) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AND3x4_ASAP7_75t_L g459 ( .A(n_425), .B(n_460), .C(n_461), .Y(n_459) );
AND2x2_ASAP7_75t_L g852 ( .A(n_425), .B(n_460), .Y(n_852) );
HB1xp67_ASAP7_75t_L g1397 ( .A(n_425), .Y(n_1397) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g560 ( .A(n_427), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g811 ( .A(n_427), .Y(n_811) );
OR2x2_ASAP7_75t_L g885 ( .A(n_427), .B(n_561), .Y(n_885) );
INVx1_ASAP7_75t_L g1428 ( .A(n_427), .Y(n_1428) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g439 ( .A(n_428), .Y(n_439) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_430), .A2(n_515), .B1(n_519), .B2(n_527), .C(n_532), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_431), .A2(n_603), .B(n_604), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_431), .A2(n_655), .B(n_656), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_431), .A2(n_749), .B(n_750), .Y(n_748) );
AOI211x1_ASAP7_75t_L g974 ( .A1(n_431), .A2(n_975), .B(n_976), .C(n_998), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_431), .B(n_1077), .Y(n_1076) );
AOI21xp33_ASAP7_75t_L g1088 ( .A1(n_431), .A2(n_1089), .B(n_1090), .Y(n_1088) );
NAND2xp33_ASAP7_75t_L g1155 ( .A(n_431), .B(n_1156), .Y(n_1155) );
AOI21xp33_ASAP7_75t_L g1230 ( .A1(n_431), .A2(n_1231), .B(n_1232), .Y(n_1230) );
AOI211x1_ASAP7_75t_L g1288 ( .A1(n_431), .A2(n_1289), .B(n_1290), .C(n_1304), .Y(n_1288) );
AOI21xp33_ASAP7_75t_SL g1448 ( .A1(n_431), .A2(n_1449), .B(n_1450), .Y(n_1448) );
AOI21xp33_ASAP7_75t_SL g1485 ( .A1(n_431), .A2(n_1486), .B(n_1487), .Y(n_1485) );
AOI21xp5_ASAP7_75t_L g1505 ( .A1(n_431), .A2(n_1506), .B(n_1507), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_431), .B(n_1544), .Y(n_1543) );
AOI21xp33_ASAP7_75t_SL g1870 ( .A1(n_431), .A2(n_1871), .B(n_1872), .Y(n_1870) );
INVx8_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_433), .B(n_441), .Y(n_432) );
INVx1_ASAP7_75t_L g818 ( .A(n_433), .Y(n_818) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_438), .Y(n_433) );
BUFx3_ASAP7_75t_L g961 ( .A(n_434), .Y(n_961) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_435), .Y(n_679) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g669 ( .A(n_436), .Y(n_669) );
INVx2_ASAP7_75t_L g455 ( .A(n_437), .Y(n_455) );
INVx1_ASAP7_75t_L g567 ( .A(n_437), .Y(n_567) );
OR2x2_ASAP7_75t_L g564 ( .A(n_438), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g571 ( .A(n_438), .Y(n_571) );
INVx1_ASAP7_75t_L g599 ( .A(n_438), .Y(n_599) );
OR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
OR2x2_ASAP7_75t_L g662 ( .A(n_439), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_SL g898 ( .A(n_439), .B(n_526), .Y(n_898) );
INVx1_ASAP7_75t_L g1350 ( .A(n_439), .Y(n_1350) );
HB1xp67_ASAP7_75t_L g1399 ( .A(n_439), .Y(n_1399) );
INVx1_ASAP7_75t_L g839 ( .A(n_440), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_441), .B(n_916), .Y(n_915) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_444), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g484 ( .A(n_443), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_443), .B(n_506), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
AND2x6_ASAP7_75t_L g532 ( .A(n_445), .B(n_521), .Y(n_532) );
AND2x2_ASAP7_75t_L g551 ( .A(n_445), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_445), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g629 ( .A(n_445), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_445), .B(n_462), .Y(n_890) );
AND2x2_ASAP7_75t_L g505 ( .A(n_446), .B(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g529 ( .A(n_446), .Y(n_529) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_446), .Y(n_693) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_447), .Y(n_782) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_457), .C(n_488), .Y(n_450) );
INVx2_ASAP7_75t_SL g601 ( .A(n_451), .Y(n_601) );
AND5x1_ASAP7_75t_L g921 ( .A(n_451), .B(n_922), .C(n_949), .D(n_965), .E(n_969), .Y(n_921) );
AND4x1_ASAP7_75t_L g1116 ( .A(n_451), .B(n_1117), .C(n_1120), .D(n_1130), .Y(n_1116) );
NAND5xp2_ASAP7_75t_L g1238 ( .A(n_451), .B(n_1239), .C(n_1242), .D(n_1244), .E(n_1245), .Y(n_1238) );
NAND4xp75_ASAP7_75t_L g1504 ( .A(n_451), .B(n_1505), .C(n_1508), .D(n_1525), .Y(n_1504) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_452), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_452), .B(n_735), .C(n_747), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_452), .A2(n_684), .B1(n_780), .B2(n_802), .C(n_803), .Y(n_801) );
INVx3_ASAP7_75t_L g984 ( .A(n_452), .Y(n_984) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
BUFx2_ASAP7_75t_L g584 ( .A(n_453), .Y(n_584) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g466 ( .A(n_454), .Y(n_466) );
BUFx3_ASAP7_75t_L g487 ( .A(n_454), .Y(n_487) );
BUFx2_ASAP7_75t_L g672 ( .A(n_454), .Y(n_672) );
INVx2_ASAP7_75t_L g746 ( .A(n_454), .Y(n_746) );
BUFx2_ASAP7_75t_L g1122 ( .A(n_454), .Y(n_1122) );
INVx1_ASAP7_75t_L g477 ( .A(n_455), .Y(n_477) );
NAND2x1_ASAP7_75t_L g491 ( .A(n_456), .B(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g495 ( .A(n_456), .B(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g580 ( .A(n_456), .B(n_492), .Y(n_580) );
AND2x4_ASAP7_75t_SL g684 ( .A(n_456), .B(n_496), .Y(n_684) );
AND2x4_ASAP7_75t_SL g802 ( .A(n_456), .B(n_492), .Y(n_802) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_456), .B(n_492), .Y(n_1132) );
AOI33xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_463), .A3(n_467), .B1(n_478), .B2(n_480), .B3(n_486), .Y(n_457) );
AOI33xp33_ASAP7_75t_L g582 ( .A1(n_458), .A2(n_480), .A3(n_583), .B1(n_585), .B2(n_591), .B3(n_592), .Y(n_582) );
AOI33xp33_ASAP7_75t_L g985 ( .A1(n_458), .A2(n_986), .A3(n_989), .B1(n_991), .B2(n_992), .B3(n_994), .Y(n_985) );
AOI33xp33_ASAP7_75t_L g1296 ( .A1(n_458), .A2(n_482), .A3(n_1297), .B1(n_1299), .B2(n_1300), .B3(n_1303), .Y(n_1296) );
AOI33xp33_ASAP7_75t_L g1515 ( .A1(n_458), .A2(n_1154), .A3(n_1516), .B1(n_1517), .B2(n_1520), .B3(n_1523), .Y(n_1515) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI33xp33_ASAP7_75t_L g790 ( .A1(n_459), .A2(n_791), .A3(n_792), .B1(n_794), .B2(n_796), .B3(n_798), .Y(n_790) );
AOI33xp33_ASAP7_75t_L g1041 ( .A1(n_459), .A2(n_1042), .A3(n_1044), .B1(n_1047), .B2(n_1048), .B3(n_1049), .Y(n_1041) );
AOI33xp33_ASAP7_75t_L g1120 ( .A1(n_459), .A2(n_1121), .A3(n_1123), .B1(n_1126), .B2(n_1127), .B3(n_1128), .Y(n_1120) );
AOI33xp33_ASAP7_75t_L g1146 ( .A1(n_459), .A2(n_1147), .A3(n_1148), .B1(n_1152), .B2(n_1153), .B3(n_1154), .Y(n_1146) );
AOI33xp33_ASAP7_75t_L g1437 ( .A1(n_459), .A2(n_1438), .A3(n_1439), .B1(n_1442), .B2(n_1443), .B3(n_1444), .Y(n_1437) );
AOI33xp33_ASAP7_75t_L g1479 ( .A1(n_459), .A2(n_1154), .A3(n_1480), .B1(n_1481), .B2(n_1482), .B3(n_1483), .Y(n_1479) );
AOI33xp33_ASAP7_75t_L g1565 ( .A1(n_459), .A2(n_1566), .A3(n_1567), .B1(n_1568), .B2(n_1569), .B3(n_1570), .Y(n_1565) );
NAND3xp33_ASAP7_75t_L g1803 ( .A(n_459), .B(n_1804), .C(n_1806), .Y(n_1803) );
AOI33xp33_ASAP7_75t_L g1878 ( .A1(n_459), .A2(n_1443), .A3(n_1879), .B1(n_1880), .B2(n_1881), .B3(n_1882), .Y(n_1878) );
INVx3_ASAP7_75t_L g1383 ( .A(n_460), .Y(n_1383) );
INVx1_ASAP7_75t_L g649 ( .A(n_461), .Y(n_649) );
OAI31xp33_ASAP7_75t_L g835 ( .A1(n_461), .A2(n_836), .A3(n_840), .B(n_866), .Y(n_835) );
INVx2_ASAP7_75t_SL g1467 ( .A(n_461), .Y(n_1467) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g557 ( .A(n_462), .Y(n_557) );
BUFx2_ASAP7_75t_L g1298 ( .A(n_464), .Y(n_1298) );
INVx8_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g570 ( .A(n_465), .Y(n_570) );
INVx3_ASAP7_75t_L g995 ( .A(n_465), .Y(n_995) );
INVx2_ASAP7_75t_L g1280 ( .A(n_465), .Y(n_1280) );
INVx1_ASAP7_75t_L g997 ( .A(n_466), .Y(n_997) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_469), .A2(n_856), .B1(n_1205), .B2(n_1206), .Y(n_1204) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
AND2x4_ASAP7_75t_L g572 ( .A(n_470), .B(n_571), .Y(n_572) );
INVx2_ASAP7_75t_SL g738 ( .A(n_470), .Y(n_738) );
INVx3_ASAP7_75t_L g1302 ( .A(n_470), .Y(n_1302) );
INVx3_ASAP7_75t_L g1441 ( .A(n_470), .Y(n_1441) );
HB1xp67_ASAP7_75t_L g1518 ( .A(n_470), .Y(n_1518) );
BUFx8_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g588 ( .A(n_471), .Y(n_588) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_471), .Y(n_676) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_471), .Y(n_850) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g990 ( .A(n_474), .Y(n_990) );
INVx2_ASAP7_75t_R g1046 ( .A(n_474), .Y(n_1046) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g479 ( .A(n_475), .Y(n_479) );
BUFx12f_ASAP7_75t_L g590 ( .A(n_475), .Y(n_590) );
AND2x4_ASAP7_75t_L g917 ( .A(n_475), .B(n_839), .Y(n_917) );
BUFx2_ASAP7_75t_L g1151 ( .A(n_475), .Y(n_1151) );
BUFx3_ASAP7_75t_L g1519 ( .A(n_475), .Y(n_1519) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx2_ASAP7_75t_L g493 ( .A(n_476), .Y(n_493) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_476), .B(n_567), .Y(n_566) );
BUFx2_ASAP7_75t_L g1384 ( .A(n_476), .Y(n_1384) );
INVx1_ASAP7_75t_L g498 ( .A(n_477), .Y(n_498) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_481), .A2(n_736), .B1(n_737), .B2(n_742), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g673 ( .A(n_482), .Y(n_673) );
INVx2_ASAP7_75t_L g958 ( .A(n_482), .Y(n_958) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx3_ASAP7_75t_L g993 ( .A(n_483), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_494), .B2(n_495), .Y(n_488) );
AOI222xp33_ASAP7_75t_L g533 ( .A1(n_489), .A2(n_494), .B1(n_534), .B2(n_536), .C1(n_538), .C2(n_549), .Y(n_533) );
AOI221x1_ASAP7_75t_L g949 ( .A1(n_490), .A2(n_495), .B1(n_925), .B2(n_931), .C(n_950), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_490), .A2(n_495), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_490), .A2(n_495), .B1(n_1435), .B2(n_1436), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1476 ( .A1(n_490), .A2(n_495), .B1(n_1477), .B2(n_1478), .Y(n_1476) );
AOI22xp33_ASAP7_75t_L g1509 ( .A1(n_490), .A2(n_495), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_495), .A2(n_579), .B1(n_580), .B2(n_581), .Y(n_578) );
AO22x1_ASAP7_75t_L g978 ( .A1(n_495), .A2(n_580), .B1(n_979), .B2(n_980), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_495), .A2(n_1131), .B1(n_1132), .B2(n_1133), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_495), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_495), .A2(n_580), .B1(n_1240), .B2(n_1241), .Y(n_1239) );
AOI22xp5_ASAP7_75t_L g1291 ( .A1(n_495), .A2(n_1132), .B1(n_1292), .B2(n_1293), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1875 ( .A1(n_495), .A2(n_1132), .B1(n_1876), .B2(n_1877), .Y(n_1875) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_554), .B(n_558), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_514), .C(n_533), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B1(n_508), .B2(n_509), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_502), .A2(n_508), .B1(n_569), .B2(n_572), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_503), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_504), .A2(n_510), .B1(n_695), .B2(n_696), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g1057 ( .A1(n_504), .A2(n_510), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_504), .A2(n_509), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_504), .A2(n_510), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
INVx1_ASAP7_75t_L g1265 ( .A(n_504), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_504), .A2(n_509), .B1(n_1315), .B2(n_1316), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_504), .A2(n_510), .B1(n_1513), .B2(n_1514), .Y(n_1530) );
AOI22xp33_ASAP7_75t_L g1557 ( .A1(n_504), .A2(n_510), .B1(n_1558), .B2(n_1559), .Y(n_1557) );
AOI22xp33_ASAP7_75t_L g1852 ( .A1(n_504), .A2(n_515), .B1(n_1853), .B2(n_1854), .Y(n_1852) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_505), .A2(n_510), .B1(n_722), .B2(n_723), .Y(n_721) );
AND2x4_ASAP7_75t_L g833 ( .A(n_505), .B(n_811), .Y(n_833) );
INVx1_ASAP7_75t_L g1006 ( .A(n_505), .Y(n_1006) );
AND2x4_ASAP7_75t_L g510 ( .A(n_506), .B(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g515 ( .A(n_506), .B(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_SL g535 ( .A(n_506), .B(n_521), .Y(n_535) );
AND2x2_ASAP7_75t_L g762 ( .A(n_506), .B(n_763), .Y(n_762) );
BUFx2_ASAP7_75t_L g785 ( .A(n_506), .Y(n_785) );
AND2x2_ASAP7_75t_L g812 ( .A(n_506), .B(n_511), .Y(n_812) );
HB1xp67_ASAP7_75t_L g1405 ( .A(n_507), .Y(n_1405) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_509), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1458 ( .A1(n_509), .A2(n_1005), .B1(n_1459), .B2(n_1460), .Y(n_1458) );
AOI22xp33_ASAP7_75t_L g1500 ( .A1(n_509), .A2(n_1005), .B1(n_1501), .B2(n_1502), .Y(n_1500) );
AOI21xp5_ASAP7_75t_L g1850 ( .A1(n_509), .A2(n_532), .B(n_1851), .Y(n_1850) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g620 ( .A(n_510), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_510), .A2(n_1000), .B1(n_1001), .B2(n_1005), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_510), .Y(n_1229) );
INVx2_ASAP7_75t_L g546 ( .A(n_511), .Y(n_546) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_511), .Y(n_644) );
INVx1_ASAP7_75t_L g718 ( .A(n_511), .Y(n_718) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx3_ASAP7_75t_L g524 ( .A(n_512), .Y(n_524) );
INVx2_ASAP7_75t_L g768 ( .A(n_512), .Y(n_768) );
AND2x4_ASAP7_75t_L g1404 ( .A(n_512), .B(n_1405), .Y(n_1404) );
INVx3_ASAP7_75t_L g608 ( .A(n_515), .Y(n_608) );
INVx2_ASAP7_75t_SL g687 ( .A(n_515), .Y(n_687) );
NAND2xp5_ASAP7_75t_R g1013 ( .A(n_515), .B(n_983), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_515), .B(n_1040), .Y(n_1060) );
INVx1_ASAP7_75t_L g1323 ( .A(n_516), .Y(n_1323) );
BUFx2_ASAP7_75t_L g1860 ( .A(n_516), .Y(n_1860) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g531 ( .A(n_517), .Y(n_531) );
INVx2_ASAP7_75t_L g707 ( .A(n_517), .Y(n_707) );
BUFx3_ASAP7_75t_L g720 ( .A(n_517), .Y(n_720) );
BUFx3_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_521), .Y(n_613) );
BUFx3_ASAP7_75t_L g716 ( .A(n_521), .Y(n_716) );
INVx1_ASAP7_75t_L g1099 ( .A(n_521), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1216 ( .A(n_521), .Y(n_1216) );
BUFx3_ASAP7_75t_L g1312 ( .A(n_521), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_521), .B(n_1418), .Y(n_1417) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g542 ( .A(n_522), .Y(n_542) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g1179 ( .A(n_524), .Y(n_1179) );
INVx1_ASAP7_75t_L g1795 ( .A(n_524), .Y(n_1795) );
HB1xp67_ASAP7_75t_SL g1223 ( .A(n_525), .Y(n_1223) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_SL g614 ( .A(n_526), .Y(n_614) );
INVx4_ASAP7_75t_L g774 ( .A(n_526), .Y(n_774) );
NAND4xp25_ASAP7_75t_L g936 ( .A(n_526), .B(n_937), .C(n_938), .D(n_940), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_526), .B(n_1349), .Y(n_1348) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_SL g537 ( .A(n_529), .Y(n_537) );
INVx2_ASAP7_75t_L g771 ( .A(n_529), .Y(n_771) );
INVx1_ASAP7_75t_L g939 ( .A(n_529), .Y(n_939) );
INVx2_ASAP7_75t_L g1010 ( .A(n_529), .Y(n_1010) );
INVx1_ASAP7_75t_L g1225 ( .A(n_529), .Y(n_1225) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_SL g1012 ( .A(n_531), .Y(n_1012) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_532), .A2(n_610), .B(n_615), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_532), .A2(n_689), .B(n_690), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_532), .A2(n_715), .B(n_719), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g1007 ( .A1(n_532), .A2(n_1008), .B(n_1009), .Y(n_1007) );
INVx1_ASAP7_75t_L g1061 ( .A(n_532), .Y(n_1061) );
AOI21xp5_ASAP7_75t_L g1096 ( .A1(n_532), .A2(n_1097), .B(n_1102), .Y(n_1096) );
AOI21xp5_ASAP7_75t_L g1167 ( .A1(n_532), .A2(n_1168), .B(n_1169), .Y(n_1167) );
AOI21xp5_ASAP7_75t_L g1220 ( .A1(n_532), .A2(n_1221), .B(n_1224), .Y(n_1220) );
AOI21xp5_ASAP7_75t_L g1310 ( .A1(n_532), .A2(n_1311), .B(n_1313), .Y(n_1310) );
AOI21xp5_ASAP7_75t_SL g1453 ( .A1(n_532), .A2(n_1454), .B(n_1457), .Y(n_1453) );
AOI21xp5_ASAP7_75t_L g1497 ( .A1(n_532), .A2(n_1498), .B(n_1499), .Y(n_1497) );
AOI21xp5_ASAP7_75t_SL g1527 ( .A1(n_532), .A2(n_1528), .B(n_1529), .Y(n_1527) );
AOI221xp5_ASAP7_75t_L g1553 ( .A1(n_532), .A2(n_762), .B1(n_1554), .B2(n_1555), .C(n_1556), .Y(n_1553) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_534), .B(n_925), .Y(n_924) );
AOI222xp33_ASAP7_75t_L g1547 ( .A1(n_534), .A2(n_551), .B1(n_1548), .B2(n_1549), .C1(n_1550), .C2(n_1552), .Y(n_1547) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g624 ( .A(n_535), .Y(n_624) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g1825 ( .A(n_541), .B(n_1418), .Y(n_1825) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g642 ( .A(n_542), .Y(n_642) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g1456 ( .A(n_545), .Y(n_1456) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g1495 ( .A(n_546), .Y(n_1495) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g645 ( .A(n_548), .Y(n_645) );
INVx2_ASAP7_75t_L g704 ( .A(n_548), .Y(n_704) );
INVx3_ASAP7_75t_L g769 ( .A(n_548), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g1016 ( .A1(n_548), .A2(n_1017), .B1(n_1018), .B2(n_1019), .C(n_1022), .Y(n_1016) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_552), .A2(n_780), .B1(n_781), .B2(n_783), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_552), .A2(n_781), .B1(n_931), .B2(n_932), .Y(n_930) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g628 ( .A(n_553), .Y(n_628) );
INVx1_ASAP7_75t_L g892 ( .A(n_553), .Y(n_892) );
AND2x4_ASAP7_75t_L g1421 ( .A(n_553), .B(n_1414), .Y(n_1421) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_554), .A2(n_686), .B(n_697), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g1002 ( .A1(n_554), .A2(n_1003), .B(n_1014), .Y(n_1002) );
OAI21xp5_ASAP7_75t_L g1165 ( .A1(n_554), .A2(n_1166), .B(n_1174), .Y(n_1165) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g1324 ( .A(n_555), .Y(n_1324) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_556), .B(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g1115 ( .A(n_556), .Y(n_1115) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x6_ASAP7_75t_L g799 ( .A(n_557), .B(n_800), .Y(n_799) );
AND2x4_ASAP7_75t_L g879 ( .A(n_557), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g1161 ( .A(n_559), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_559), .Y(n_1233) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
AND2x4_ASAP7_75t_L g657 ( .A(n_560), .B(n_564), .Y(n_657) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g815 ( .A(n_564), .Y(n_815) );
INVx3_ASAP7_75t_L g860 ( .A(n_565), .Y(n_860) );
BUFx6f_ASAP7_75t_L g1360 ( .A(n_565), .Y(n_1360) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g847 ( .A(n_566), .Y(n_847) );
BUFx3_ASAP7_75t_L g1365 ( .A(n_566), .Y(n_1365) );
BUFx2_ASAP7_75t_L g1388 ( .A(n_567), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_569), .A2(n_572), .B1(n_695), .B2(n_696), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_569), .A2(n_572), .B1(n_722), .B2(n_723), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_569), .A2(n_572), .B1(n_1000), .B2(n_1001), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1245 ( .A(n_569), .B(n_1246), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_569), .A2(n_807), .B1(n_1558), .B2(n_1559), .Y(n_1561) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x4_ASAP7_75t_L g816 ( .A(n_570), .B(n_571), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_570), .A2(n_797), .B1(n_832), .B2(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g600 ( .A(n_572), .Y(n_600) );
INVx2_ASAP7_75t_L g1119 ( .A(n_572), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1512 ( .A1(n_572), .A2(n_816), .B1(n_1513), .B2(n_1514), .Y(n_1512) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_602), .C(n_606), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_593), .C(n_601), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_582), .Y(n_577) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_588), .A2(n_665), .B1(n_666), .B2(n_670), .C(n_671), .Y(n_664) );
INVx3_ASAP7_75t_L g808 ( .A(n_588), .Y(n_808) );
OR2x6_ASAP7_75t_SL g837 ( .A(n_588), .B(n_838), .Y(n_837) );
BUFx2_ASAP7_75t_L g1522 ( .A(n_588), .Y(n_1522) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_594), .B(n_968), .Y(n_967) );
OR2x6_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_595), .B(n_598), .Y(n_1164) );
INVx2_ASAP7_75t_SL g1200 ( .A(n_595), .Y(n_1200) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx4f_ASAP7_75t_L g842 ( .A(n_597), .Y(n_842) );
OR2x4_ASAP7_75t_L g1371 ( .A(n_597), .B(n_1372), .Y(n_1371) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g807 ( .A(n_599), .B(n_808), .Y(n_807) );
NOR4xp25_ASAP7_75t_L g1188 ( .A(n_601), .B(n_1189), .C(n_1192), .D(n_1193), .Y(n_1188) );
NOR3xp33_ASAP7_75t_L g1432 ( .A(n_601), .B(n_1433), .C(n_1447), .Y(n_1432) );
NOR3xp33_ASAP7_75t_L g1474 ( .A(n_601), .B(n_1475), .C(n_1484), .Y(n_1474) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_605), .B(n_910), .Y(n_909) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_621), .B(n_646), .Y(n_606) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g1455 ( .A(n_613), .Y(n_1455) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g725 ( .A(n_623), .Y(n_725) );
INVx1_ASAP7_75t_L g1015 ( .A(n_623), .Y(n_1015) );
INVx4_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g1258 ( .A(n_627), .Y(n_1258) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g784 ( .A(n_629), .Y(n_784) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B1(n_635), .B2(n_639), .C(n_640), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_631), .A2(n_1024), .B1(n_1025), .B2(n_1026), .Y(n_1023) );
OAI221xp5_ASAP7_75t_L g1462 ( .A1(n_631), .A2(n_1110), .B1(n_1463), .B2(n_1464), .C(n_1465), .Y(n_1462) );
OAI221xp5_ASAP7_75t_L g1490 ( .A1(n_631), .A2(n_1026), .B1(n_1491), .B2(n_1492), .C(n_1493), .Y(n_1490) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g777 ( .A(n_633), .Y(n_777) );
INVx4_ASAP7_75t_L g928 ( .A(n_633), .Y(n_928) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx4_ASAP7_75t_L g935 ( .A(n_636), .Y(n_935) );
BUFx6f_ASAP7_75t_L g1027 ( .A(n_636), .Y(n_1027) );
INVx2_ASAP7_75t_L g1073 ( .A(n_636), .Y(n_1073) );
INVx2_ASAP7_75t_L g1111 ( .A(n_636), .Y(n_1111) );
INVx2_ASAP7_75t_SL g1253 ( .A(n_636), .Y(n_1253) );
INVx8_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g1261 ( .A(n_637), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1413 ( .A(n_637), .B(n_1414), .Y(n_1413) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g1551 ( .A(n_642), .Y(n_1551) );
BUFx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g1211 ( .A1(n_646), .A2(n_1212), .B(n_1219), .Y(n_1211) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_648), .Y(n_945) );
INVx1_ASAP7_75t_L g1869 ( .A(n_648), .Y(n_1869) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx2_ASAP7_75t_L g733 ( .A(n_649), .Y(n_733) );
AOI21x1_ASAP7_75t_L g759 ( .A1(n_649), .A2(n_760), .B(n_788), .Y(n_759) );
HB1xp67_ASAP7_75t_L g1537 ( .A(n_649), .Y(n_1537) );
BUFx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AO22x2_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_709), .B1(n_710), .B2(n_752), .Y(n_651) );
INVx1_ASAP7_75t_L g752 ( .A(n_652), .Y(n_752) );
AND4x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_658), .C(n_685), .D(n_708), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .C(n_682), .Y(n_658) );
OAI22xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_664), .B1(n_673), .B2(n_674), .Y(n_660) );
BUFx3_ASAP7_75t_L g1355 ( .A(n_661), .Y(n_1355) );
BUFx4f_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx8_ASAP7_75t_L g736 ( .A(n_662), .Y(n_736) );
BUFx2_ASAP7_75t_L g951 ( .A(n_662), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_666), .A2(n_738), .B1(n_739), .B2(n_740), .C(n_741), .Y(n_737) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx3_ASAP7_75t_L g1278 ( .A(n_669), .Y(n_1278) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B1(n_678), .B2(n_680), .C(n_681), .Y(n_674) );
INVx1_ASAP7_75t_L g1045 ( .A(n_675), .Y(n_1045) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_676), .Y(n_793) );
BUFx6f_ASAP7_75t_L g795 ( .A(n_676), .Y(n_795) );
INVx2_ASAP7_75t_L g1125 ( .A(n_676), .Y(n_1125) );
INVx2_ASAP7_75t_L g1271 ( .A(n_676), .Y(n_1271) );
AND2x4_ASAP7_75t_L g1394 ( .A(n_676), .B(n_1372), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1834 ( .A(n_676), .B(n_1372), .Y(n_1834) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_677), .A2(n_699), .B(n_703), .C(n_705), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_678), .A2(n_727), .B1(n_738), .B2(n_743), .C(n_744), .Y(n_742) );
CKINVDCx8_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
INVx3_ASAP7_75t_L g844 ( .A(n_679), .Y(n_844) );
INVx3_ASAP7_75t_L g856 ( .A(n_679), .Y(n_856) );
INVx3_ASAP7_75t_L g954 ( .A(n_679), .Y(n_954) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_684), .A2(n_802), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_684), .A2(n_802), .B1(n_1548), .B2(n_1549), .Y(n_1564) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g1797 ( .A(n_692), .Y(n_1797) );
INVx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx6f_ASAP7_75t_L g1170 ( .A(n_693), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_693), .B(n_1414), .Y(n_1816) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g778 ( .A(n_700), .Y(n_778) );
INVx2_ASAP7_75t_L g929 ( .A(n_700), .Y(n_929) );
INVx4_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx4f_ASAP7_75t_L g787 ( .A(n_701), .Y(n_787) );
OR2x6_ASAP7_75t_L g905 ( .A(n_701), .B(n_906), .Y(n_905) );
BUFx4f_ASAP7_75t_L g1017 ( .A(n_701), .Y(n_1017) );
BUFx4f_ASAP7_75t_L g1054 ( .A(n_701), .Y(n_1054) );
BUFx6f_ASAP7_75t_L g1336 ( .A(n_701), .Y(n_1336) );
BUFx4f_ASAP7_75t_L g1858 ( .A(n_701), .Y(n_1858) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
BUFx3_ASAP7_75t_L g730 ( .A(n_702), .Y(n_730) );
INVx1_ASAP7_75t_L g1067 ( .A(n_704), .Y(n_1067) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g763 ( .A(n_707), .Y(n_763) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND4x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_734), .C(n_748), .D(n_751), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_724), .B(n_733), .Y(n_712) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B(n_731), .C(n_732), .Y(n_726) );
OAI211xp5_ASAP7_75t_L g941 ( .A1(n_728), .A2(n_942), .B(n_943), .C(n_944), .Y(n_941) );
OAI211xp5_ASAP7_75t_L g1318 ( .A1(n_728), .A2(n_1319), .B(n_1320), .C(n_1321), .Y(n_1318) );
INVx5_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g894 ( .A(n_730), .B(n_895), .Y(n_894) );
O2A1O1Ixp5_ASAP7_75t_SL g1050 ( .A1(n_733), .A2(n_1051), .B(n_1062), .C(n_1074), .Y(n_1050) );
OAI33xp33_ASAP7_75t_L g1193 ( .A1(n_736), .A2(n_1194), .A3(n_1198), .B1(n_1204), .B2(n_1207), .B3(n_1210), .Y(n_1193) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g797 ( .A(n_746), .Y(n_797) );
INVx1_ASAP7_75t_L g1043 ( .A(n_746), .Y(n_1043) );
INVx1_ASAP7_75t_L g1281 ( .A(n_746), .Y(n_1281) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AO22x2_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_972), .B1(n_1029), .B2(n_1030), .Y(n_754) );
INVx1_ASAP7_75t_L g1029 ( .A(n_755), .Y(n_1029) );
XNOR2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_920), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_827), .B1(n_918), .B2(n_919), .Y(n_756) );
INVx1_ASAP7_75t_L g919 ( .A(n_757), .Y(n_919) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_820), .C(n_824), .Y(n_757) );
INVx1_ASAP7_75t_L g821 ( .A(n_759), .Y(n_821) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g911 ( .A(n_763), .B(n_912), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_770), .B2(n_772), .Y(n_764) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g773 ( .A(n_768), .Y(n_773) );
INVx1_ASAP7_75t_L g1101 ( .A(n_773), .Y(n_1101) );
INVx2_ASAP7_75t_L g1218 ( .A(n_773), .Y(n_1218) );
HB1xp67_ASAP7_75t_L g1222 ( .A(n_773), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_775) );
OAI211xp5_ASAP7_75t_L g1175 ( .A1(n_778), .A2(n_1176), .B(n_1177), .C(n_1180), .Y(n_1175) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AOI222xp33_ASAP7_75t_L g814 ( .A1(n_783), .A2(n_815), .B1(n_816), .B2(n_817), .C1(n_818), .C2(n_819), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g926 ( .A1(n_784), .A2(n_785), .B1(n_927), .B2(n_933), .Y(n_926) );
INVx1_ASAP7_75t_L g822 ( .A(n_789), .Y(n_822) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_801), .Y(n_789) );
INVx1_ASAP7_75t_L g1363 ( .A(n_795), .Y(n_1363) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1049 ( .A(n_799), .Y(n_1049) );
INVx1_ASAP7_75t_SL g1570 ( .A(n_799), .Y(n_1570) );
INVx1_ASAP7_75t_L g826 ( .A(n_804), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_813), .Y(n_804) );
NAND2x1_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .Y(n_805) );
INVx2_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_807), .A2(n_816), .B1(n_1058), .B2(n_1059), .Y(n_1075) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_810), .A2(n_832), .B1(n_833), .B2(n_834), .Y(n_831) );
AND2x4_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
INVx1_ASAP7_75t_L g825 ( .A(n_814), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_815), .A2(n_818), .B1(n_932), .B2(n_948), .Y(n_947) );
OAI21xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B(n_823), .Y(n_820) );
OAI21xp33_ASAP7_75t_L g824 ( .A1(n_823), .A2(n_825), .B(n_826), .Y(n_824) );
INVx1_ASAP7_75t_L g918 ( .A(n_827), .Y(n_918) );
XNOR2xp5_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
NOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_875), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_835), .Y(n_830) );
INVx3_ASAP7_75t_L g968 ( .A(n_833), .Y(n_968) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_839), .Y(n_870) );
OAI221xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_846), .B1(n_853), .B2(n_858), .C(n_864), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_844), .B2(n_845), .Y(n_841) );
INVx1_ASAP7_75t_L g1274 ( .A(n_842), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_842), .Y(n_1357) );
OAI221xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .B1(n_849), .B2(n_851), .C(n_852), .Y(n_846) );
OR2x6_ASAP7_75t_L g864 ( .A(n_847), .B(n_865), .Y(n_864) );
OAI211xp5_ASAP7_75t_L g899 ( .A1(n_848), .A2(n_900), .B(n_903), .C(n_904), .Y(n_899) );
INVx3_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_SL g854 ( .A(n_850), .Y(n_854) );
INVx5_ASAP7_75t_L g960 ( .A(n_850), .Y(n_960) );
INVx2_ASAP7_75t_SL g1150 ( .A(n_850), .Y(n_1150) );
HB1xp67_ASAP7_75t_L g1805 ( .A(n_850), .Y(n_1805) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_856), .B2(n_857), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_854), .A2(n_953), .B1(n_954), .B2(n_955), .C(n_956), .Y(n_952) );
OAI22xp33_ASAP7_75t_L g1194 ( .A1(n_856), .A2(n_1195), .B1(n_1196), .B2(n_1197), .Y(n_1194) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_856), .A2(n_1125), .B1(n_1333), .B2(n_1344), .Y(n_1361) );
OAI21xp5_ASAP7_75t_SL g858 ( .A1(n_859), .A2(n_861), .B(n_862), .Y(n_858) );
INVx3_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g1196 ( .A(n_860), .Y(n_1196) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_863), .Y(n_1129) );
INVx1_ASAP7_75t_L g1808 ( .A(n_863), .Y(n_1808) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_868), .A2(n_884), .B1(n_886), .B2(n_887), .Y(n_883) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx4_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NAND3xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_907), .C(n_913), .Y(n_875) );
NOR3xp33_ASAP7_75t_SL g876 ( .A(n_877), .B(n_893), .C(n_896), .Y(n_876) );
OAI21xp5_ASAP7_75t_SL g877 ( .A1(n_878), .A2(n_882), .B(n_883), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_881), .Y(n_878) );
INVx2_ASAP7_75t_L g1337 ( .A(n_879), .Y(n_1337) );
INVx4_ASAP7_75t_L g1799 ( .A(n_879), .Y(n_1799) );
INVx1_ASAP7_75t_SL g884 ( .A(n_885), .Y(n_884) );
INVx2_ASAP7_75t_SL g887 ( .A(n_888), .Y(n_887) );
NAND2x2_ASAP7_75t_L g888 ( .A(n_889), .B(n_891), .Y(n_888) );
INVx1_ASAP7_75t_L g906 ( .A(n_889), .Y(n_906) );
INVx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_SL g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g912 ( .A(n_895), .Y(n_912) );
OAI21xp5_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_899), .B(n_905), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NAND3xp33_ASAP7_75t_L g1800 ( .A(n_898), .B(n_1801), .C(n_1802), .Y(n_1800) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
BUFx2_ASAP7_75t_L g934 ( .A(n_902), .Y(n_934) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_902), .Y(n_1021) );
BUFx3_ASAP7_75t_L g1065 ( .A(n_902), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_945), .B(n_946), .Y(n_922) );
NAND4xp25_ASAP7_75t_L g923 ( .A(n_924), .B(n_926), .C(n_936), .D(n_941), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_929), .A2(n_1064), .B1(n_1065), .B2(n_1066), .C(n_1067), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_934), .A2(n_1333), .B1(n_1334), .B2(n_1335), .Y(n_1332) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_934), .A2(n_1341), .B1(n_1352), .B2(n_1353), .Y(n_1351) );
INVx2_ASAP7_75t_L g1342 ( .A(n_935), .Y(n_1342) );
OAI221xp5_ASAP7_75t_L g959 ( .A1(n_942), .A2(n_960), .B1(n_961), .B2(n_962), .C(n_963), .Y(n_959) );
OAI22xp5_ASAP7_75t_SL g950 ( .A1(n_951), .A2(n_952), .B1(n_958), .B2(n_959), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_954), .A2(n_1251), .B1(n_1270), .B2(n_1271), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_954), .A2(n_1273), .B1(n_1340), .B2(n_1353), .Y(n_1366) );
INVx2_ASAP7_75t_SL g988 ( .A(n_957), .Y(n_988) );
INVx1_ASAP7_75t_L g1446 ( .A(n_957), .Y(n_1446) );
BUFx3_ASAP7_75t_L g1524 ( .A(n_957), .Y(n_1524) );
BUFx3_ASAP7_75t_L g1202 ( .A(n_960), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_967), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_971), .B(n_983), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_971), .B(n_1040), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_971), .B(n_1145), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_971), .B(n_1295), .Y(n_1294) );
INVx2_ASAP7_75t_L g1030 ( .A(n_972), .Y(n_1030) );
XOR2x2_ASAP7_75t_L g972 ( .A(n_973), .B(n_1028), .Y(n_972) );
NAND2xp5_ASAP7_75t_SL g973 ( .A(n_974), .B(n_1002), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_977), .B(n_985), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_978), .B(n_981), .Y(n_977) );
NAND2xp5_ASAP7_75t_SL g981 ( .A(n_982), .B(n_984), .Y(n_981) );
AND4x1_ASAP7_75t_L g1035 ( .A(n_984), .B(n_1036), .C(n_1039), .D(n_1041), .Y(n_1035) );
NAND4xp25_ASAP7_75t_SL g1140 ( .A(n_984), .B(n_1141), .C(n_1144), .D(n_1146), .Y(n_1140) );
NAND4xp25_ASAP7_75t_SL g1290 ( .A(n_984), .B(n_1291), .C(n_1294), .D(n_1296), .Y(n_1290) );
INVx1_ASAP7_75t_L g1884 ( .A(n_984), .Y(n_1884) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
BUFx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
BUFx2_ASAP7_75t_L g1127 ( .A(n_993), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_993), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1443 ( .A(n_993), .Y(n_1443) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
NAND3xp33_ASAP7_75t_SL g1003 ( .A(n_1004), .B(n_1007), .C(n_1013), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_1005), .A2(n_1227), .B1(n_1228), .B2(n_1229), .Y(n_1226) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_SL g1011 ( .A(n_1012), .Y(n_1011) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx4_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx5_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1032), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
XOR2xp5_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1078), .Y(n_1033) );
NAND3xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1050), .C(n_1076), .Y(n_1034) );
NAND4xp25_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1057), .C(n_1060), .D(n_1061), .Y(n_1051) );
OAI211xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1054), .B(n_1055), .C(n_1056), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .B1(n_1072), .B2(n_1073), .Y(n_1068) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
XNOR2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1283), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
XNOR2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1235), .Y(n_1082) );
XNOR2x1_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1185), .Y(n_1083) );
OAI22x1_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1135), .B1(n_1136), .B2(n_1184), .Y(n_1084) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1085), .Y(n_1184) );
AO21x2_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1087), .B(n_1134), .Y(n_1085) );
NAND3xp33_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1091), .C(n_1116), .Y(n_1087) );
OAI21xp5_ASAP7_75t_L g1091 ( .A1(n_1092), .A2(n_1103), .B(n_1115), .Y(n_1091) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1099), .Y(n_1114) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1099), .Y(n_1536) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1108), .B1(n_1109), .B2(n_1112), .C(n_1113), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_1105), .A2(n_1339), .B1(n_1340), .B2(n_1341), .Y(n_1338) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_1105), .A2(n_1336), .B1(n_1344), .B2(n_1345), .Y(n_1343) );
INVx2_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_1107), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g1214 ( .A(n_1107), .Y(n_1214) );
OAI221xp5_ASAP7_75t_SL g1213 ( .A1(n_1109), .A2(n_1201), .B1(n_1208), .B2(n_1214), .C(n_1215), .Y(n_1213) );
BUFx2_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1532 ( .A1(n_1110), .A2(n_1214), .B1(n_1533), .B2(n_1534), .C(n_1535), .Y(n_1532) );
BUFx6f_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
OAI31xp33_ASAP7_75t_L g1248 ( .A1(n_1115), .A2(n_1249), .A3(n_1256), .B(n_1264), .Y(n_1248) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
AOI222xp33_ASAP7_75t_L g1836 ( .A1(n_1122), .A2(n_1387), .B1(n_1820), .B2(n_1821), .C1(n_1822), .C2(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1127), .Y(n_1210) );
NAND3xp33_ASAP7_75t_L g1809 ( .A(n_1127), .B(n_1810), .C(n_1811), .Y(n_1809) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
NAND2x1p5_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1157), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1155), .Y(n_1138) );
INVxp67_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NOR2xp33_ASAP7_75t_SL g1181 ( .A(n_1140), .B(n_1182), .Y(n_1181) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1155), .B(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1165), .Y(n_1159) );
AOI21xp5_ASAP7_75t_L g1160 ( .A1(n_1161), .A2(n_1162), .B(n_1163), .Y(n_1160) );
AOI21xp5_ASAP7_75t_SL g1266 ( .A1(n_1161), .A2(n_1267), .B(n_1268), .Y(n_1266) );
AOI21xp5_ASAP7_75t_L g1305 ( .A1(n_1161), .A2(n_1306), .B(n_1307), .Y(n_1305) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
AND3x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1211), .C(n_1230), .Y(n_1187) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
OAI22xp33_ASAP7_75t_L g1207 ( .A1(n_1196), .A2(n_1199), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
OAI22xp33_ASAP7_75t_L g1272 ( .A1(n_1196), .A2(n_1260), .B1(n_1273), .B2(n_1275), .Y(n_1272) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
OAI221xp5_ASAP7_75t_L g1276 ( .A1(n_1202), .A2(n_1254), .B1(n_1277), .B2(n_1278), .C(n_1279), .Y(n_1276) );
OAI33xp33_ASAP7_75t_L g1354 ( .A1(n_1210), .A2(n_1355), .A3(n_1356), .B1(n_1361), .B2(n_1362), .B3(n_1366), .Y(n_1354) );
OAI221xp5_ASAP7_75t_L g1250 ( .A1(n_1214), .A2(n_1251), .B1(n_1252), .B2(n_1254), .C(n_1255), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1259 ( .A1(n_1214), .A2(n_1260), .B1(n_1261), .B2(n_1262), .C(n_1263), .Y(n_1259) );
OAI221xp5_ASAP7_75t_L g1862 ( .A1(n_1214), .A2(n_1863), .B1(n_1864), .B2(n_1865), .C(n_1866), .Y(n_1862) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx2_ASAP7_75t_L g1466 ( .A(n_1218), .Y(n_1466) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
XNOR2x1_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1282), .Y(n_1236) );
NOR2x1_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1247), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1266), .Y(n_1247) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
HB1xp67_ASAP7_75t_L g1864 ( .A(n_1253), .Y(n_1864) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_1284), .A2(n_1285), .B1(n_1325), .B2(n_1326), .Y(n_1283) );
INVx1_ASAP7_75t_SL g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
XNOR2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1308), .Y(n_1304) );
OAI21xp33_ASAP7_75t_L g1308 ( .A1(n_1309), .A2(n_1317), .B(n_1324), .Y(n_1308) );
AOI222xp33_ASAP7_75t_L g1819 ( .A1(n_1312), .A2(n_1421), .B1(n_1820), .B2(n_1821), .C1(n_1822), .C2(n_1823), .Y(n_1819) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
AOI21xp5_ASAP7_75t_L g1545 ( .A1(n_1324), .A2(n_1546), .B(n_1560), .Y(n_1545) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
XNOR2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1469), .Y(n_1326) );
OA22x2_ASAP7_75t_L g1327 ( .A1(n_1328), .A2(n_1429), .B1(n_1430), .B2(n_1468), .Y(n_1327) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1328), .Y(n_1468) );
NAND3xp33_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1367), .C(n_1400), .Y(n_1329) );
NOR2xp33_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1354), .Y(n_1330) );
OAI33xp33_ASAP7_75t_L g1331 ( .A1(n_1332), .A2(n_1337), .A3(n_1338), .B1(n_1343), .B2(n_1346), .B3(n_1351), .Y(n_1331) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_1334), .A2(n_1345), .B1(n_1363), .B2(n_1364), .Y(n_1362) );
HB1xp67_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
OAI22xp33_ASAP7_75t_L g1356 ( .A1(n_1339), .A2(n_1352), .B1(n_1357), .B2(n_1358), .Y(n_1356) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
INVx2_ASAP7_75t_SL g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
BUFx6f_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
OAI31xp33_ASAP7_75t_L g1367 ( .A1(n_1368), .A2(n_1376), .A3(n_1389), .B(n_1395), .Y(n_1367) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1838 ( .A1(n_1370), .A2(n_1374), .B1(n_1815), .B2(n_1817), .Y(n_1838) );
INVx2_ASAP7_75t_SL g1370 ( .A(n_1371), .Y(n_1370) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx2_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
NAND3xp33_ASAP7_75t_L g1835 ( .A(n_1377), .B(n_1836), .C(n_1838), .Y(n_1835) );
CKINVDCx8_ASAP7_75t_R g1377 ( .A(n_1378), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1381), .B1(n_1385), .B2(n_1386), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_1380), .A2(n_1420), .B1(n_1422), .B2(n_1423), .Y(n_1419) );
BUFx3_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
BUFx3_ASAP7_75t_L g1837 ( .A(n_1382), .Y(n_1837) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1384), .Y(n_1382) );
AND2x4_ASAP7_75t_L g1387 ( .A(n_1383), .B(n_1388), .Y(n_1387) );
BUFx6f_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx2_ASAP7_75t_SL g1832 ( .A(n_1392), .Y(n_1832) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
AND2x2_ASAP7_75t_SL g1395 ( .A(n_1396), .B(n_1398), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1839 ( .A(n_1396), .B(n_1398), .Y(n_1839) );
INVx1_ASAP7_75t_SL g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
OAI31xp33_ASAP7_75t_SL g1400 ( .A1(n_1401), .A2(n_1406), .A3(n_1415), .B(n_1426), .Y(n_1400) );
INVx3_ASAP7_75t_SL g1403 ( .A(n_1404), .Y(n_1403) );
CKINVDCx16_ASAP7_75t_R g1827 ( .A(n_1404), .Y(n_1827) );
HB1xp67_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
INVx2_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
INVx2_ASAP7_75t_L g1818 ( .A(n_1413), .Y(n_1818) );
INVx3_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
BUFx3_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
INVx2_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
INVx2_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
BUFx3_ASAP7_75t_L g1823 ( .A(n_1425), .Y(n_1823) );
BUFx3_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
BUFx2_ASAP7_75t_SL g1828 ( .A(n_1427), .Y(n_1828) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
NAND3xp33_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1448), .C(n_1451), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1437), .Y(n_1433) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
OAI21xp5_ASAP7_75t_L g1451 ( .A1(n_1452), .A2(n_1461), .B(n_1467), .Y(n_1451) );
OAI21xp5_ASAP7_75t_L g1488 ( .A1(n_1467), .A2(n_1489), .B(n_1496), .Y(n_1488) );
AOI22xp5_ASAP7_75t_L g1469 ( .A1(n_1470), .A2(n_1471), .B1(n_1538), .B2(n_1539), .Y(n_1469) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
XNOR2x1_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1503), .Y(n_1471) );
NAND3xp33_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1485), .C(n_1488), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1479), .Y(n_1475) );
BUFx2_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
AND3x1_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1512), .C(n_1515), .Y(n_1508) );
INVx2_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
OAI21xp5_ASAP7_75t_L g1525 ( .A1(n_1526), .A2(n_1531), .B(n_1537), .Y(n_1525) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
HB1xp67_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
NAND3xp33_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1545), .C(n_1562), .Y(n_1542) );
NAND3xp33_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1553), .C(n_1557), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
OAI221xp5_ASAP7_75t_L g1572 ( .A1(n_1573), .A2(n_1786), .B1(n_1789), .B2(n_1840), .C(n_1843), .Y(n_1572) );
AOI21xp5_ASAP7_75t_L g1573 ( .A1(n_1574), .A2(n_1697), .B(n_1756), .Y(n_1573) );
NAND5xp2_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1640), .C(n_1660), .D(n_1673), .E(n_1683), .Y(n_1574) );
O2A1O1Ixp33_ASAP7_75t_L g1575 ( .A1(n_1576), .A2(n_1607), .B(n_1614), .C(n_1625), .Y(n_1575) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1576), .Y(n_1644) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1577), .B(n_1597), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1577), .B(n_1604), .Y(n_1633) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1577), .B(n_1599), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1577), .B(n_1598), .Y(n_1701) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1577), .B(n_1710), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1745 ( .A(n_1577), .B(n_1611), .Y(n_1745) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1577), .Y(n_1768) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1593), .Y(n_1577) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1578), .B(n_1639), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1578), .B(n_1598), .Y(n_1651) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1578), .B(n_1594), .Y(n_1659) );
AND3x1_ASAP7_75t_L g1733 ( .A(n_1578), .B(n_1594), .C(n_1598), .Y(n_1733) );
OR2x2_ASAP7_75t_L g1774 ( .A(n_1578), .B(n_1639), .Y(n_1774) );
INVx2_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1579), .B(n_1593), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_1579), .B(n_1594), .Y(n_1664) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1587), .Y(n_1579) );
INVx2_ASAP7_75t_L g1694 ( .A(n_1581), .Y(n_1694) );
AND2x6_ASAP7_75t_L g1581 ( .A(n_1582), .B(n_1583), .Y(n_1581) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1582), .B(n_1586), .Y(n_1585) );
AND2x4_ASAP7_75t_L g1588 ( .A(n_1582), .B(n_1589), .Y(n_1588) );
AND2x6_ASAP7_75t_L g1591 ( .A(n_1582), .B(n_1592), .Y(n_1591) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1582), .B(n_1586), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1623 ( .A(n_1582), .B(n_1586), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1788 ( .A(n_1582), .B(n_1589), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1589 ( .A(n_1584), .B(n_1590), .Y(n_1589) );
INVxp67_ASAP7_75t_L g1696 ( .A(n_1585), .Y(n_1696) );
HB1xp67_ASAP7_75t_L g1894 ( .A(n_1589), .Y(n_1894) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1593), .B(n_1639), .Y(n_1736) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
OR2x2_ASAP7_75t_L g1669 ( .A(n_1594), .B(n_1639), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1594), .B(n_1639), .Y(n_1730) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_1595), .B(n_1596), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1597), .B(n_1659), .Y(n_1658) );
NAND2xp5_ASAP7_75t_L g1744 ( .A(n_1597), .B(n_1664), .Y(n_1744) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1597), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1603), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1598), .B(n_1613), .Y(n_1679) );
OR2x2_ASAP7_75t_L g1681 ( .A(n_1598), .B(n_1682), .Y(n_1681) );
INVx2_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1599), .B(n_1613), .Y(n_1612) );
OAI322xp33_ASAP7_75t_L g1625 ( .A1(n_1599), .A2(n_1621), .A3(n_1626), .B1(n_1632), .B2(n_1634), .C1(n_1636), .C2(n_1637), .Y(n_1625) );
BUFx2_ASAP7_75t_L g1639 ( .A(n_1599), .Y(n_1639) );
OR2x2_ASAP7_75t_L g1662 ( .A(n_1599), .B(n_1663), .Y(n_1662) );
AOI321xp33_ASAP7_75t_L g1683 ( .A1(n_1599), .A2(n_1684), .A3(n_1685), .B1(n_1686), .B2(n_1688), .C(n_1690), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1599), .B(n_1664), .Y(n_1721) );
OR2x2_ASAP7_75t_L g1782 ( .A(n_1599), .B(n_1716), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1601), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_1603), .B(n_1615), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_1603), .B(n_1664), .Y(n_1682) );
NOR2xp33_ASAP7_75t_L g1688 ( .A(n_1603), .B(n_1689), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1603), .B(n_1655), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1755 ( .A(n_1603), .B(n_1613), .Y(n_1755) );
OAI21xp33_ASAP7_75t_L g1776 ( .A1(n_1603), .A2(n_1755), .B(n_1777), .Y(n_1776) );
INVx2_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1604), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1604), .B(n_1617), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1604), .B(n_1621), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1604), .B(n_1639), .Y(n_1708) );
NAND2xp5_ASAP7_75t_L g1716 ( .A(n_1604), .B(n_1664), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1604), .B(n_1629), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1606), .Y(n_1604) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1612), .Y(n_1608) );
NAND2xp5_ASAP7_75t_L g1738 ( .A(n_1609), .B(n_1674), .Y(n_1738) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1626 ( .A(n_1610), .B(n_1627), .Y(n_1626) );
NOR2xp33_ASAP7_75t_L g1668 ( .A(n_1610), .B(n_1669), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1700 ( .A(n_1610), .B(n_1701), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1610), .B(n_1733), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1610), .B(n_1679), .Y(n_1740) );
INVx2_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1710 ( .A(n_1611), .B(n_1627), .Y(n_1710) );
O2A1O1Ixp33_ASAP7_75t_L g1784 ( .A1(n_1611), .A2(n_1753), .B(n_1754), .C(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1612), .Y(n_1785) );
OR2x2_ASAP7_75t_L g1684 ( .A(n_1613), .B(n_1659), .Y(n_1684) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1613), .Y(n_1754) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1620), .Y(n_1614) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1615), .B(n_1621), .Y(n_1687) );
INVx2_ASAP7_75t_L g1705 ( .A(n_1615), .Y(n_1705) );
A2O1A1O1Ixp25_ASAP7_75t_L g1750 ( .A1(n_1615), .A2(n_1629), .B(n_1707), .C(n_1751), .D(n_1752), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1765 ( .A(n_1615), .B(n_1766), .Y(n_1765) );
INVx2_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1616), .B(n_1620), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1616), .B(n_1629), .Y(n_1643) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
OR2x2_ASAP7_75t_L g1628 ( .A(n_1617), .B(n_1629), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1617), .B(n_1656), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1617), .B(n_1629), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1618), .B(n_1619), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1620), .B(n_1627), .Y(n_1636) );
NOR2xp33_ASAP7_75t_L g1667 ( .A(n_1620), .B(n_1628), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1620), .B(n_1655), .Y(n_1702) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1620), .B(n_1629), .Y(n_1712) );
OR2x2_ASAP7_75t_L g1723 ( .A(n_1620), .B(n_1629), .Y(n_1723) );
CKINVDCx6p67_ASAP7_75t_R g1620 ( .A(n_1621), .Y(n_1620) );
OR2x2_ASAP7_75t_L g1666 ( .A(n_1621), .B(n_1629), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1621), .B(n_1629), .Y(n_1674) );
NAND2xp5_ASAP7_75t_L g1747 ( .A(n_1621), .B(n_1748), .Y(n_1747) );
CKINVDCx5p33_ASAP7_75t_R g1769 ( .A(n_1621), .Y(n_1769) );
OR2x2_ASAP7_75t_L g1772 ( .A(n_1621), .B(n_1642), .Y(n_1772) );
OR2x6_ASAP7_75t_L g1621 ( .A(n_1622), .B(n_1624), .Y(n_1621) );
OR2x2_ASAP7_75t_L g1725 ( .A(n_1622), .B(n_1624), .Y(n_1725) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1626), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1652 ( .A(n_1627), .B(n_1633), .Y(n_1652) );
INVx2_ASAP7_75t_L g1627 ( .A(n_1628), .Y(n_1627) );
INVx3_ASAP7_75t_L g1647 ( .A(n_1629), .Y(n_1647) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1629), .Y(n_1656) );
AOI22xp5_ASAP7_75t_L g1673 ( .A1(n_1629), .A2(n_1674), .B1(n_1675), .B2(n_1680), .Y(n_1673) );
AND2x4_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1631), .Y(n_1629) );
INVxp67_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1671 ( .A(n_1635), .B(n_1672), .Y(n_1671) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1636), .Y(n_1783) );
CKINVDCx14_ASAP7_75t_R g1637 ( .A(n_1638), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1639), .B(n_1659), .Y(n_1713) );
NOR2xp33_ASAP7_75t_L g1640 ( .A(n_1641), .B(n_1653), .Y(n_1640) );
OAI211xp5_ASAP7_75t_L g1641 ( .A1(n_1642), .A2(n_1644), .B(n_1645), .C(n_1652), .Y(n_1641) );
AOI21xp33_ASAP7_75t_L g1714 ( .A1(n_1642), .A2(n_1715), .B(n_1716), .Y(n_1714) );
CKINVDCx6p67_ASAP7_75t_R g1642 ( .A(n_1643), .Y(n_1642) );
AOI21xp33_ASAP7_75t_L g1778 ( .A1(n_1644), .A2(n_1719), .B(n_1779), .Y(n_1778) );
NAND2xp5_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1648), .Y(n_1645) );
CKINVDCx14_ASAP7_75t_R g1646 ( .A(n_1647), .Y(n_1646) );
AOI221xp5_ASAP7_75t_L g1780 ( .A1(n_1648), .A2(n_1674), .B1(n_1781), .B2(n_1783), .C(n_1784), .Y(n_1780) );
NOR2xp33_ASAP7_75t_L g1648 ( .A(n_1649), .B(n_1651), .Y(n_1648) );
CKINVDCx14_ASAP7_75t_R g1649 ( .A(n_1650), .Y(n_1649) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1651), .Y(n_1748) );
NOR2xp33_ASAP7_75t_L g1653 ( .A(n_1654), .B(n_1657), .Y(n_1653) );
AOI21xp5_ASAP7_75t_L g1759 ( .A1(n_1654), .A2(n_1760), .B(n_1761), .Y(n_1759) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1659), .Y(n_1689) );
AOI221xp5_ASAP7_75t_L g1660 ( .A1(n_1661), .A2(n_1665), .B1(n_1667), .B2(n_1668), .C(n_1670), .Y(n_1660) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1662), .B(n_1735), .Y(n_1734) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1664), .B(n_1708), .Y(n_1707) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1666), .B(n_1672), .Y(n_1715) );
OAI221xp5_ASAP7_75t_L g1752 ( .A1(n_1666), .A2(n_1690), .B1(n_1753), .B2(n_1754), .C(n_1755), .Y(n_1752) );
AOI221xp5_ASAP7_75t_L g1762 ( .A1(n_1667), .A2(n_1701), .B1(n_1763), .B2(n_1769), .C(n_1770), .Y(n_1762) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
AOI222xp33_ASAP7_75t_L g1726 ( .A1(n_1674), .A2(n_1727), .B1(n_1731), .B2(n_1732), .C1(n_1734), .C2(n_1737), .Y(n_1726) );
NAND2xp5_ASAP7_75t_L g1753 ( .A(n_1674), .B(n_1705), .Y(n_1753) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
NOR2xp33_ASAP7_75t_L g1724 ( .A(n_1676), .B(n_1725), .Y(n_1724) );
NAND2xp5_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1679), .Y(n_1676) );
OAI21xp33_ASAP7_75t_L g1711 ( .A1(n_1677), .A2(n_1712), .B(n_1713), .Y(n_1711) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1679), .Y(n_1728) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
AOI211xp5_ASAP7_75t_SL g1770 ( .A1(n_1682), .A2(n_1771), .B(n_1772), .C(n_1773), .Y(n_1770) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
OAI22xp5_ASAP7_75t_L g1741 ( .A1(n_1687), .A2(n_1742), .B1(n_1744), .B2(n_1745), .Y(n_1741) );
INVx2_ASAP7_75t_SL g1690 ( .A(n_1691), .Y(n_1690) );
OAI22xp5_ASAP7_75t_SL g1692 ( .A1(n_1693), .A2(n_1694), .B1(n_1695), .B2(n_1696), .Y(n_1692) );
NAND5xp2_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1717), .C(n_1726), .D(n_1739), .E(n_1750), .Y(n_1697) );
AOI211xp5_ASAP7_75t_L g1698 ( .A1(n_1699), .A2(n_1702), .B(n_1703), .C(n_1714), .Y(n_1698) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
AOI221xp5_ASAP7_75t_L g1775 ( .A1(n_1702), .A2(n_1732), .B1(n_1743), .B2(n_1776), .C(n_1778), .Y(n_1775) );
OAI211xp5_ASAP7_75t_L g1703 ( .A1(n_1704), .A2(n_1706), .B(n_1709), .C(n_1711), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1719 ( .A(n_1704), .B(n_1720), .Y(n_1719) );
INVx2_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1708), .Y(n_1767) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1710), .Y(n_1749) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1712), .Y(n_1779) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1713), .Y(n_1777) );
INVxp67_ASAP7_75t_SL g1751 ( .A(n_1715), .Y(n_1751) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1716), .Y(n_1720) );
O2A1O1Ixp33_ASAP7_75t_SL g1717 ( .A1(n_1718), .A2(n_1721), .B(n_1722), .C(n_1724), .Y(n_1717) );
INVxp67_ASAP7_75t_SL g1718 ( .A(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1721), .Y(n_1761) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
AOI211xp5_ASAP7_75t_L g1739 ( .A1(n_1725), .A2(n_1740), .B(n_1741), .C(n_1746), .Y(n_1739) );
A2O1A1Ixp33_ASAP7_75t_L g1757 ( .A1(n_1725), .A2(n_1730), .B(n_1758), .C(n_1759), .Y(n_1757) );
NAND2xp5_ASAP7_75t_SL g1727 ( .A(n_1728), .B(n_1729), .Y(n_1727) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
AOI21xp33_ASAP7_75t_L g1746 ( .A1(n_1735), .A2(n_1747), .B(n_1749), .Y(n_1746) );
OAI21xp33_ASAP7_75t_L g1763 ( .A1(n_1735), .A2(n_1764), .B(n_1765), .Y(n_1763) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVxp67_ASAP7_75t_SL g1737 ( .A(n_1738), .Y(n_1737) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1740), .Y(n_1760) );
INVx2_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
NAND4xp25_ASAP7_75t_L g1756 ( .A(n_1757), .B(n_1762), .C(n_1775), .D(n_1780), .Y(n_1756) );
OR2x2_ASAP7_75t_L g1766 ( .A(n_1767), .B(n_1768), .Y(n_1766) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1774), .Y(n_1773) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
CKINVDCx20_ASAP7_75t_R g1786 ( .A(n_1787), .Y(n_1786) );
CKINVDCx5p33_ASAP7_75t_R g1787 ( .A(n_1788), .Y(n_1787) );
NAND3xp33_ASAP7_75t_L g1790 ( .A(n_1791), .B(n_1812), .C(n_1829), .Y(n_1790) );
AND4x1_ASAP7_75t_L g1791 ( .A(n_1792), .B(n_1800), .C(n_1803), .D(n_1809), .Y(n_1791) );
NAND3xp33_ASAP7_75t_L g1792 ( .A(n_1793), .B(n_1796), .C(n_1798), .Y(n_1792) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
INVx2_ASAP7_75t_SL g1798 ( .A(n_1799), .Y(n_1798) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
OAI21xp5_ASAP7_75t_L g1812 ( .A1(n_1813), .A2(n_1826), .B(n_1828), .Y(n_1812) );
NAND3xp33_ASAP7_75t_L g1813 ( .A(n_1814), .B(n_1819), .C(n_1824), .Y(n_1813) );
AOI22xp33_ASAP7_75t_L g1814 ( .A1(n_1815), .A2(n_1816), .B1(n_1817), .B2(n_1818), .Y(n_1814) );
INVx2_ASAP7_75t_L g1824 ( .A(n_1825), .Y(n_1824) );
OAI21xp5_ASAP7_75t_L g1829 ( .A1(n_1830), .A2(n_1835), .B(n_1839), .Y(n_1829) );
INVx2_ASAP7_75t_SL g1831 ( .A(n_1832), .Y(n_1831) );
INVx2_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
CKINVDCx5p33_ASAP7_75t_R g1840 ( .A(n_1841), .Y(n_1840) );
INVxp33_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
HB1xp67_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
NAND3xp33_ASAP7_75t_L g1847 ( .A(n_1848), .B(n_1870), .C(n_1873), .Y(n_1847) );
OAI31xp33_ASAP7_75t_L g1848 ( .A1(n_1849), .A2(n_1855), .A3(n_1867), .B(n_1868), .Y(n_1848) );
NAND2xp5_ASAP7_75t_L g1849 ( .A(n_1850), .B(n_1852), .Y(n_1849) );
OAI211xp5_ASAP7_75t_L g1856 ( .A1(n_1857), .A2(n_1858), .B(n_1859), .C(n_1861), .Y(n_1856) );
INVx1_ASAP7_75t_L g1868 ( .A(n_1869), .Y(n_1868) );
NOR3xp33_ASAP7_75t_L g1873 ( .A(n_1874), .B(n_1883), .C(n_1884), .Y(n_1873) );
NAND2xp5_ASAP7_75t_L g1874 ( .A(n_1875), .B(n_1878), .Y(n_1874) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1886), .Y(n_1885) );
INVx1_ASAP7_75t_L g1886 ( .A(n_1887), .Y(n_1886) );
HB1xp67_ASAP7_75t_L g1887 ( .A(n_1888), .Y(n_1887) );
BUFx3_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
HB1xp67_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
HB1xp67_ASAP7_75t_L g1891 ( .A(n_1892), .Y(n_1891) );
OAI21xp5_ASAP7_75t_L g1892 ( .A1(n_1893), .A2(n_1894), .B(n_1895), .Y(n_1892) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1896), .Y(n_1895) );
endmodule