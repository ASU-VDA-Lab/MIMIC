module fake_netlist_1_643_n_1185 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1185);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1185;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1174;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1078;
wire n_1097;
wire n_572;
wire n_1125;
wire n_324;
wire n_1016;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_1132;
wire n_1155;
wire n_1101;
wire n_1159;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_1160;
wire n_1184;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_729;
wire n_519;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1017;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_1178;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_1157;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_1110;
wire n_327;
wire n_944;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_58), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_123), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_159), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_202), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_104), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_211), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_169), .B(n_204), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_111), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_103), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_270), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_15), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_21), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_229), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_44), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_212), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_42), .Y(n_293) );
CKINVDCx16_ASAP7_75t_R g294 ( .A(n_225), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_248), .Y(n_295) );
CKINVDCx16_ASAP7_75t_R g296 ( .A(n_40), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_98), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_28), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_183), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_266), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_104), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_210), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_186), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_209), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_61), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_236), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_222), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_219), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_0), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_124), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_44), .B(n_240), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_237), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_217), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_245), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_99), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_78), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_140), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_172), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_71), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_150), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_168), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_26), .B(n_190), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_132), .Y(n_323) );
INVxp33_ASAP7_75t_SL g324 ( .A(n_139), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_167), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_189), .Y(n_326) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_249), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_61), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_114), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_36), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_19), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_93), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_21), .Y(n_333) );
INVxp33_ASAP7_75t_L g334 ( .A(n_160), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_235), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_164), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_263), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_22), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_181), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_208), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_52), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_256), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_257), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_109), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_110), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_118), .B(n_180), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_221), .Y(n_347) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_214), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_259), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_262), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_51), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_233), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_275), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_241), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_82), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_226), .Y(n_356) );
CKINVDCx16_ASAP7_75t_R g357 ( .A(n_246), .Y(n_357) );
NOR2xp67_ASAP7_75t_L g358 ( .A(n_265), .B(n_3), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_51), .Y(n_359) );
BUFx10_ASAP7_75t_L g360 ( .A(n_14), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_254), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_195), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_112), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_231), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_220), .B(n_46), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_15), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_234), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_207), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_232), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_117), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_134), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_244), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_192), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_170), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_37), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_126), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_193), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_53), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_196), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g380 ( .A(n_97), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_267), .Y(n_381) );
CKINVDCx14_ASAP7_75t_R g382 ( .A(n_90), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_121), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_264), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_1), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_218), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_260), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_3), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_251), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_131), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_108), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_2), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_216), .B(n_162), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_129), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_75), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_105), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_47), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_96), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_153), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_125), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_178), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_191), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_261), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_80), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_17), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_185), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_252), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_66), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_98), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_27), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_239), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_64), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_188), .B(n_227), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_305), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_305), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_362), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_328), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_303), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_408), .B(n_0), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_328), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_285), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_376), .B(n_2), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_290), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_378), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_290), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_323), .B(n_4), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_290), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_394), .B(n_4), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_334), .B(n_5), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_333), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_290), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_340), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_405), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_333), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_340), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_338), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_338), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_296), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_340), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_340), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_351), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_378), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_319), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_279), .Y(n_447) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_284), .B(n_277), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_280), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_319), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_403), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_303), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_403), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_447), .B(n_300), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_448), .A2(n_288), .B1(n_289), .B2(n_282), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_428), .Y(n_457) );
BUFx10_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_447), .B(n_450), .Y(n_459) );
AND2x6_ASAP7_75t_L g460 ( .A(n_432), .B(n_393), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_424), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_415), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_419), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_415), .Y(n_466) );
INVx3_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_436), .B(n_380), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_417), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_419), .Y(n_471) );
INVx5_ASAP7_75t_L g472 ( .A(n_428), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_450), .B(n_300), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_417), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_426), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_422), .B(n_310), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_427), .B(n_304), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_427), .B(n_304), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_422), .B(n_402), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_426), .B(n_294), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_448), .A2(n_293), .B1(n_301), .B2(n_298), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_428), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_446), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_422), .B(n_348), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_430), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_436), .B(n_357), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_430), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_430), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_453), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_432), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_430), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_445), .B(n_308), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_430), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_432), .B(n_407), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_448), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_494), .B(n_429), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_498), .B(n_441), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_464), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_498), .B(n_453), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_499), .A2(n_297), .B1(n_309), .B2(n_278), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_464), .Y(n_506) );
AND2x6_ASAP7_75t_SL g507 ( .A(n_476), .B(n_420), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_461), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_459), .B(n_431), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_459), .B(n_420), .Y(n_510) );
INVx5_ASAP7_75t_L g511 ( .A(n_460), .Y(n_511) );
NAND2xp33_ASAP7_75t_L g512 ( .A(n_460), .B(n_283), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_465), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_476), .B(n_324), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_499), .B(n_295), .Y(n_515) );
AND3x1_ASAP7_75t_L g516 ( .A(n_456), .B(n_441), .C(n_316), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_499), .A2(n_416), .B1(n_418), .B2(n_414), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_482), .B(n_324), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_475), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_499), .B(n_299), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_465), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_466), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_458), .B(n_302), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_458), .B(n_306), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_458), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_458), .B(n_313), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_471), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_471), .B(n_317), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_487), .B(n_281), .Y(n_529) );
AO22x1_ASAP7_75t_L g530 ( .A1(n_460), .A2(n_392), .B1(n_331), .B2(n_291), .Y(n_530) );
OR2x6_ASAP7_75t_L g531 ( .A(n_468), .B(n_423), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_482), .B(n_414), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_479), .B(n_416), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_469), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_469), .Y(n_535) );
NOR2x2_ASAP7_75t_L g536 ( .A(n_489), .B(n_278), .Y(n_536) );
INVx4_ASAP7_75t_L g537 ( .A(n_460), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_489), .B(n_360), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_471), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_489), .B(n_468), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_470), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_491), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_481), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_481), .B(n_421), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_468), .B(n_360), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_470), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_483), .B(n_307), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_460), .B(n_421), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_491), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_484), .A2(n_437), .B1(n_439), .B2(n_433), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_493), .A2(n_413), .B(n_312), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_460), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_484), .A2(n_349), .B1(n_374), .B2(n_314), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_455), .B(n_437), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_455), .B(n_314), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_473), .B(n_439), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_493), .B(n_440), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_467), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_467), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_467), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_496), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_493), .B(n_318), .Y(n_564) );
BUFx2_ASAP7_75t_L g565 ( .A(n_486), .Y(n_565) );
AND2x6_ASAP7_75t_SL g566 ( .A(n_477), .B(n_315), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_486), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_477), .B(n_320), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_478), .B(n_444), .Y(n_569) );
NOR2xp33_ASAP7_75t_R g570 ( .A(n_472), .B(n_349), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_472), .B(n_325), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_472), .B(n_392), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_525), .B(n_374), .Y(n_573) );
AND2x6_ASAP7_75t_L g574 ( .A(n_563), .B(n_390), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_540), .B(n_297), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_515), .A2(n_365), .B(n_327), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_520), .A2(n_381), .B(n_364), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_511), .B(n_396), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_516), .A2(n_396), .B1(n_406), .B2(n_401), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_521), .Y(n_580) );
BUFx3_ASAP7_75t_L g581 ( .A(n_508), .Y(n_581) );
AOI21x1_ASAP7_75t_L g582 ( .A1(n_520), .A2(n_462), .B(n_457), .Y(n_582) );
AOI21x1_ASAP7_75t_L g583 ( .A1(n_564), .A2(n_462), .B(n_457), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_510), .B(n_286), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_509), .A2(n_411), .B(n_386), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_501), .A2(n_406), .B1(n_330), .B2(n_332), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_504), .A2(n_336), .B(n_329), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_500), .B(n_341), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_533), .B(n_355), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_570), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_519), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_544), .B(n_359), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_538), .B(n_388), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_537), .A2(n_404), .B1(n_409), .B2(n_398), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_521), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_523), .A2(n_343), .B(n_342), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_557), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_531), .B(n_404), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_511), .Y(n_599) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_558), .Y(n_601) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_549), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_524), .A2(n_347), .B(n_345), .Y(n_603) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_549), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_545), .B(n_507), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_524), .A2(n_352), .B(n_350), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_557), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_555), .B(n_366), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_530), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_511), .B(n_287), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_526), .A2(n_356), .B(n_353), .Y(n_611) );
CKINVDCx6p67_ASAP7_75t_R g612 ( .A(n_531), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_553), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_526), .A2(n_367), .B(n_363), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_554), .B(n_375), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_564), .A2(n_369), .B(n_368), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_503), .Y(n_617) );
AOI21x1_ASAP7_75t_L g618 ( .A1(n_571), .A2(n_485), .B(n_480), .Y(n_618) );
BUFx12f_ASAP7_75t_L g619 ( .A(n_566), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_553), .B(n_292), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_532), .A2(n_371), .B(n_370), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_572), .B(n_321), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_569), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_517), .B(n_514), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_518), .B(n_397), .Y(n_625) );
INVx4_ASAP7_75t_L g626 ( .A(n_560), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_548), .A2(n_410), .B(n_412), .C(n_395), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_560), .Y(n_628) );
NOR2xp33_ASAP7_75t_SL g629 ( .A(n_547), .B(n_335), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_502), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_550), .B(n_337), .Y(n_631) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_529), .B(n_8), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_565), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_506), .B(n_339), .Y(n_634) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_568), .B(n_372), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_522), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_534), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_535), .A2(n_546), .B(n_556), .C(n_541), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_559), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_512), .B(n_385), .C(n_319), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_567), .B(n_344), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_513), .A2(n_539), .B(n_527), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_505), .A2(n_358), .B1(n_379), .B2(n_373), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_542), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_561), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_562), .Y(n_646) );
INVx4_ASAP7_75t_L g647 ( .A(n_551), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_568), .B(n_9), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_528), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_528), .Y(n_650) );
AOI22x1_ASAP7_75t_L g651 ( .A1(n_571), .A2(n_434), .B1(n_438), .B2(n_425), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_543), .B(n_311), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_515), .A2(n_384), .B(n_383), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_540), .B(n_385), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_543), .B(n_311), .Y(n_655) );
AO21x2_ASAP7_75t_L g656 ( .A1(n_552), .A2(n_389), .B(n_387), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_563), .A2(n_322), .B(n_400), .C(n_399), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_540), .B(n_10), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_563), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_521), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_563), .A2(n_312), .B(n_326), .C(n_308), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_537), .Y(n_662) );
INVx11_ASAP7_75t_L g663 ( .A(n_536), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_563), .Y(n_664) );
INVx3_ASAP7_75t_L g665 ( .A(n_537), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_525), .B(n_377), .Y(n_666) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_600), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_624), .A2(n_497), .B(n_485), .Y(n_668) );
AO21x1_ASAP7_75t_L g669 ( .A1(n_642), .A2(n_346), .B(n_425), .Y(n_669) );
OAI21x1_ASAP7_75t_L g670 ( .A1(n_583), .A2(n_361), .B(n_354), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_575), .B(n_11), .Y(n_671) );
OAI21x1_ASAP7_75t_L g672 ( .A1(n_618), .A2(n_361), .B(n_354), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_638), .A2(n_497), .B(n_490), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_659), .B(n_391), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_591), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g676 ( .A(n_663), .Y(n_676) );
INVx4_ASAP7_75t_L g677 ( .A(n_626), .Y(n_677) );
AO32x2_ASAP7_75t_L g678 ( .A1(n_643), .A2(n_449), .A3(n_443), .B1(n_435), .B2(n_434), .Y(n_678) );
AO32x2_ASAP7_75t_L g679 ( .A1(n_643), .A2(n_435), .A3(n_449), .B1(n_443), .B2(n_442), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_623), .A2(n_490), .B(n_488), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_594), .B(n_12), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_664), .Y(n_682) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_600), .Y(n_683) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_597), .A2(n_451), .B1(n_438), .B2(n_442), .C(n_425), .Y(n_684) );
O2A1O1Ixp5_ASAP7_75t_L g685 ( .A1(n_631), .A2(n_488), .B(n_495), .C(n_492), .Y(n_685) );
NOR2xp33_ASAP7_75t_SL g686 ( .A(n_594), .B(n_452), .Y(n_686) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_600), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_630), .Y(n_688) );
OAI21x1_ASAP7_75t_L g689 ( .A1(n_582), .A2(n_495), .B(n_492), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_636), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_639), .A2(n_454), .B1(n_443), .B2(n_449), .Y(n_691) );
AO31x2_ASAP7_75t_L g692 ( .A1(n_661), .A2(n_443), .A3(n_449), .B(n_435), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_637), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_658), .B(n_13), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_628), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_645), .Y(n_696) );
BUFx3_ASAP7_75t_L g697 ( .A(n_612), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_584), .A2(n_463), .B(n_472), .Y(n_698) );
NOR2xp33_ASAP7_75t_SL g699 ( .A(n_629), .B(n_435), .Y(n_699) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_602), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_654), .Y(n_701) );
AO32x2_ASAP7_75t_L g702 ( .A1(n_579), .A2(n_16), .A3(n_17), .B1(n_18), .B2(n_19), .Y(n_702) );
AO31x2_ASAP7_75t_L g703 ( .A1(n_657), .A2(n_463), .A3(n_23), .B(n_18), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_607), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_626), .Y(n_705) );
AO31x2_ASAP7_75t_L g706 ( .A1(n_621), .A2(n_463), .A3(n_25), .B(n_20), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_648), .Y(n_707) );
AO22x2_ASAP7_75t_L g708 ( .A1(n_578), .A2(n_25), .B1(n_20), .B2(n_24), .Y(n_708) );
AND2x2_ASAP7_75t_SL g709 ( .A(n_609), .B(n_24), .Y(n_709) );
AO31x2_ASAP7_75t_L g710 ( .A1(n_580), .A2(n_463), .A3(n_30), .B(n_26), .Y(n_710) );
AO21x2_ASAP7_75t_L g711 ( .A1(n_656), .A2(n_463), .B(n_107), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_617), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_652), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_574), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_627), .A2(n_472), .B(n_463), .C(n_31), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_653), .A2(n_472), .B(n_463), .C(n_31), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_646), .Y(n_717) );
INVx5_ASAP7_75t_L g718 ( .A(n_574), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_644), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_625), .A2(n_608), .B(n_622), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_615), .B(n_29), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_586), .B(n_32), .Y(n_722) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_633), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_585), .A2(n_113), .B(n_106), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_655), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_650), .A2(n_116), .B(n_115), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_589), .A2(n_120), .B(n_119), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_593), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_605), .B(n_35), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_592), .A2(n_127), .B(n_122), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_649), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_590), .A2(n_40), .B1(n_38), .B2(n_39), .Y(n_732) );
BUFx6f_ASAP7_75t_L g733 ( .A(n_602), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_595), .A2(n_130), .B(n_128), .Y(n_734) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_632), .A2(n_43), .B1(n_41), .B2(n_42), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_598), .A2(n_45), .B1(n_41), .B2(n_43), .Y(n_736) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_596), .A2(n_135), .B(n_133), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_660), .Y(n_738) );
O2A1O1Ixp33_ASAP7_75t_SL g739 ( .A1(n_610), .A2(n_137), .B(n_138), .C(n_136), .Y(n_739) );
BUFx10_ASAP7_75t_L g740 ( .A(n_574), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_588), .A2(n_142), .B(n_141), .Y(n_741) );
OAI21x1_ASAP7_75t_SL g742 ( .A1(n_587), .A2(n_576), .B(n_603), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_606), .A2(n_144), .B(n_143), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_611), .A2(n_146), .B(n_145), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_SL g745 ( .A1(n_640), .A2(n_184), .B(n_276), .C(n_274), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_614), .A2(n_148), .B(n_147), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_613), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_SL g748 ( .A1(n_599), .A2(n_187), .B(n_273), .C(n_272), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_651), .A2(n_151), .B(n_149), .Y(n_749) );
OAI21x1_ASAP7_75t_L g750 ( .A1(n_635), .A2(n_154), .B(n_152), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_656), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_620), .A2(n_156), .B(n_155), .Y(n_752) );
OAI22x1_ASAP7_75t_L g753 ( .A1(n_573), .A2(n_48), .B1(n_49), .B2(n_50), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_666), .A2(n_158), .B(n_157), .Y(n_754) );
INVx3_ASAP7_75t_L g755 ( .A(n_662), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_662), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_756) );
AND2x4_ASAP7_75t_L g757 ( .A(n_665), .B(n_54), .Y(n_757) );
OAI21x1_ASAP7_75t_L g758 ( .A1(n_616), .A2(n_163), .B(n_161), .Y(n_758) );
OAI21x1_ASAP7_75t_L g759 ( .A1(n_577), .A2(n_166), .B(n_165), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_634), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_SL g761 ( .A1(n_599), .A2(n_194), .B(n_271), .C(n_269), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_641), .A2(n_173), .B(n_171), .Y(n_762) );
AOI221x1_ASAP7_75t_L g763 ( .A1(n_604), .A2(n_55), .B1(n_56), .B2(n_57), .C(n_58), .Y(n_763) );
OAI21x1_ASAP7_75t_L g764 ( .A1(n_647), .A2(n_175), .B(n_174), .Y(n_764) );
AO31x2_ASAP7_75t_L g765 ( .A1(n_647), .A2(n_59), .A3(n_60), .B(n_62), .Y(n_765) );
INVx2_ASAP7_75t_SL g766 ( .A(n_581), .Y(n_766) );
BUFx12f_ASAP7_75t_L g767 ( .A(n_619), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_663), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_624), .A2(n_177), .B(n_176), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_626), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_638), .A2(n_182), .B(n_179), .Y(n_771) );
AO31x2_ASAP7_75t_L g772 ( .A1(n_661), .A2(n_63), .A3(n_64), .B(n_65), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_659), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_638), .A2(n_203), .B(n_268), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_591), .Y(n_775) );
AO31x2_ASAP7_75t_L g776 ( .A1(n_669), .A2(n_67), .A3(n_68), .B(n_69), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_713), .B(n_67), .Y(n_777) );
AO31x2_ASAP7_75t_L g778 ( .A1(n_751), .A2(n_68), .A3(n_69), .B(n_70), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_725), .B(n_70), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_682), .Y(n_780) );
AO31x2_ASAP7_75t_L g781 ( .A1(n_751), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_709), .B(n_72), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_675), .Y(n_783) );
AND2x4_ASAP7_75t_L g784 ( .A(n_677), .B(n_75), .Y(n_784) );
INVx2_ASAP7_75t_SL g785 ( .A(n_775), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_721), .B(n_76), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_671), .B(n_77), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_773), .Y(n_788) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_729), .A2(n_79), .B1(n_81), .B2(n_82), .C(n_83), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_688), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_747), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_690), .Y(n_792) );
BUFx8_ASAP7_75t_L g793 ( .A(n_767), .Y(n_793) );
INVx1_ASAP7_75t_SL g794 ( .A(n_723), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_693), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_686), .A2(n_84), .B1(n_85), .B2(n_86), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_677), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_705), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_705), .B(n_87), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_695), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_696), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_696), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_717), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_717), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_707), .B(n_88), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_715), .A2(n_89), .B(n_91), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_699), .A2(n_213), .B(n_258), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_681), .A2(n_92), .B1(n_94), .B2(n_95), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_704), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_757), .A2(n_92), .B1(n_94), .B2(n_95), .Y(n_810) );
AND2x2_ASAP7_75t_L g811 ( .A(n_722), .B(n_100), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_716), .A2(n_101), .B(n_102), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_708), .Y(n_813) );
OAI222xp33_ASAP7_75t_L g814 ( .A1(n_736), .A2(n_197), .B1(n_198), .B2(n_199), .C1(n_200), .C2(n_201), .Y(n_814) );
AO21x2_ASAP7_75t_L g815 ( .A1(n_711), .A2(n_205), .B(n_206), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_712), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_719), .Y(n_817) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_667), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_708), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_731), .B(n_215), .Y(n_820) );
INVx2_ASAP7_75t_L g821 ( .A(n_701), .Y(n_821) );
INVx1_ASAP7_75t_SL g822 ( .A(n_770), .Y(n_822) );
INVx1_ASAP7_75t_SL g823 ( .A(n_770), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_692), .Y(n_824) );
OA21x2_ASAP7_75t_L g825 ( .A1(n_771), .A2(n_223), .B(n_224), .Y(n_825) );
OA21x2_ASAP7_75t_L g826 ( .A1(n_774), .A2(n_228), .B(n_230), .Y(n_826) );
INVx4_ASAP7_75t_L g827 ( .A(n_718), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_753), .Y(n_828) );
INVx4_ASAP7_75t_SL g829 ( .A(n_765), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_692), .Y(n_830) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_667), .Y(n_831) );
INVx3_ASAP7_75t_L g832 ( .A(n_740), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_676), .Y(n_833) );
INVx4_ASAP7_75t_L g834 ( .A(n_718), .Y(n_834) );
BUFx3_ASAP7_75t_L g835 ( .A(n_766), .Y(n_835) );
AOI322xp5_ASAP7_75t_L g836 ( .A1(n_728), .A2(n_238), .A3(n_242), .B1(n_243), .B2(n_247), .C1(n_250), .C2(n_253), .Y(n_836) );
NAND2xp5_ASAP7_75t_SL g837 ( .A(n_718), .B(n_255), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_694), .B(n_760), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_673), .A2(n_742), .B(n_685), .Y(n_839) );
OAI21x1_ASAP7_75t_L g840 ( .A1(n_749), .A2(n_764), .B(n_750), .Y(n_840) );
AND2x4_ASAP7_75t_L g841 ( .A(n_697), .B(n_714), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_674), .B(n_755), .Y(n_842) );
INVxp67_ASAP7_75t_SL g843 ( .A(n_667), .Y(n_843) );
INVx3_ASAP7_75t_L g844 ( .A(n_683), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_735), .A2(n_756), .B1(n_674), .B2(n_732), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_765), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_765), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_683), .A2(n_733), .B1(n_700), .B2(n_687), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_702), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_680), .A2(n_769), .B(n_730), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_706), .Y(n_851) );
OA21x2_ASAP7_75t_L g852 ( .A1(n_759), .A2(n_763), .B(n_737), .Y(n_852) );
BUFx2_ASAP7_75t_R g853 ( .A(n_768), .Y(n_853) );
AO21x2_ASAP7_75t_L g854 ( .A1(n_727), .A2(n_761), .B(n_748), .Y(n_854) );
AOI21xp5_ASAP7_75t_L g855 ( .A1(n_741), .A2(n_724), .B(n_745), .Y(n_855) );
OAI21x1_ASAP7_75t_SL g856 ( .A1(n_754), .A2(n_762), .B(n_752), .Y(n_856) );
BUFx8_ASAP7_75t_L g857 ( .A(n_702), .Y(n_857) );
A2O1A1Ixp33_ASAP7_75t_L g858 ( .A1(n_743), .A2(n_744), .B(n_746), .C(n_726), .Y(n_858) );
A2O1A1Ixp33_ASAP7_75t_L g859 ( .A1(n_684), .A2(n_758), .B(n_734), .C(n_738), .Y(n_859) );
INVx4_ASAP7_75t_SL g860 ( .A(n_710), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_706), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_702), .Y(n_862) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_706), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_772), .B(n_703), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_772), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_772), .B(n_700), .Y(n_866) );
BUFx4f_ASAP7_75t_SL g867 ( .A(n_683), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_703), .Y(n_868) );
INVx2_ASAP7_75t_L g869 ( .A(n_703), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_687), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_687), .A2(n_700), .B1(n_733), .B2(n_691), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_710), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_710), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_678), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_739), .A2(n_733), .B(n_678), .Y(n_875) );
INVx3_ASAP7_75t_L g876 ( .A(n_678), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_679), .Y(n_877) );
OAI21x1_ASAP7_75t_L g878 ( .A1(n_672), .A2(n_670), .B(n_689), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_677), .B(n_601), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_681), .A2(n_499), .B1(n_456), .B2(n_484), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_688), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_688), .Y(n_882) );
CKINVDCx6p67_ASAP7_75t_R g883 ( .A(n_767), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_682), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_682), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_720), .A2(n_668), .B(n_698), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_682), .B(n_659), .Y(n_887) );
AND2x4_ASAP7_75t_L g888 ( .A(n_803), .B(n_804), .Y(n_888) );
BUFx4f_ASAP7_75t_L g889 ( .A(n_879), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_881), .B(n_882), .Y(n_890) );
BUFx3_ASAP7_75t_L g891 ( .A(n_867), .Y(n_891) );
OA21x2_ASAP7_75t_L g892 ( .A1(n_868), .A2(n_869), .B(n_872), .Y(n_892) );
AO21x2_ASAP7_75t_L g893 ( .A1(n_839), .A2(n_866), .B(n_875), .Y(n_893) );
OA21x2_ASAP7_75t_L g894 ( .A1(n_873), .A2(n_861), .B(n_851), .Y(n_894) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_866), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_863), .Y(n_896) );
AO21x2_ASAP7_75t_L g897 ( .A1(n_846), .A2(n_847), .B(n_874), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_780), .Y(n_898) );
AND2x2_ASAP7_75t_L g899 ( .A(n_790), .B(n_792), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_795), .B(n_816), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_880), .A2(n_828), .B1(n_808), .B2(n_813), .Y(n_901) );
AO21x2_ASAP7_75t_L g902 ( .A1(n_877), .A2(n_830), .B(n_824), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_879), .B(n_811), .Y(n_903) );
INVx2_ASAP7_75t_L g904 ( .A(n_876), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_788), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_884), .Y(n_906) );
OA21x2_ASAP7_75t_L g907 ( .A1(n_865), .A2(n_864), .B(n_886), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_885), .Y(n_908) );
OAI222xp33_ASAP7_75t_L g909 ( .A1(n_810), .A2(n_808), .B1(n_782), .B2(n_796), .C1(n_845), .C2(n_789), .Y(n_909) );
AND2x4_ASAP7_75t_L g910 ( .A(n_797), .B(n_844), .Y(n_910) );
INVx2_ASAP7_75t_L g911 ( .A(n_876), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_887), .B(n_809), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_800), .Y(n_913) );
AOI21xp5_ASAP7_75t_SL g914 ( .A1(n_825), .A2(n_826), .B(n_810), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_817), .B(n_821), .Y(n_915) );
OA21x2_ASAP7_75t_L g916 ( .A1(n_840), .A2(n_862), .B(n_849), .Y(n_916) );
INVx2_ASAP7_75t_SL g917 ( .A(n_797), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_805), .Y(n_918) );
OA21x2_ASAP7_75t_L g919 ( .A1(n_878), .A2(n_819), .B(n_855), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_805), .Y(n_920) );
HB1xp67_ASAP7_75t_L g921 ( .A(n_822), .Y(n_921) );
OA21x2_ASAP7_75t_L g922 ( .A1(n_850), .A2(n_806), .B(n_812), .Y(n_922) );
AOI22x1_ASAP7_75t_L g923 ( .A1(n_784), .A2(n_834), .B1(n_827), .B2(n_812), .Y(n_923) );
AO21x2_ASAP7_75t_L g924 ( .A1(n_815), .A2(n_859), .B(n_854), .Y(n_924) );
OR2x6_ASAP7_75t_L g925 ( .A(n_799), .B(n_784), .Y(n_925) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_818), .Y(n_926) );
OR2x2_ASAP7_75t_L g927 ( .A(n_786), .B(n_783), .Y(n_927) );
AO21x2_ASAP7_75t_L g928 ( .A1(n_815), .A2(n_854), .B(n_858), .Y(n_928) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_822), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_777), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_779), .Y(n_931) );
AO21x2_ASAP7_75t_L g932 ( .A1(n_856), .A2(n_848), .B(n_820), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_778), .Y(n_933) );
AND2x4_ASAP7_75t_L g934 ( .A(n_844), .B(n_798), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_778), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_778), .Y(n_936) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_823), .Y(n_937) );
HB1xp67_ASAP7_75t_L g938 ( .A(n_823), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_781), .Y(n_939) );
OR2x2_ASAP7_75t_L g940 ( .A(n_785), .B(n_787), .Y(n_940) );
INVx3_ASAP7_75t_L g941 ( .A(n_827), .Y(n_941) );
INVx3_ASAP7_75t_L g942 ( .A(n_834), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_818), .Y(n_943) );
INVx3_ASAP7_75t_L g944 ( .A(n_818), .Y(n_944) );
BUFx2_ASAP7_75t_L g945 ( .A(n_835), .Y(n_945) );
OR2x2_ASAP7_75t_L g946 ( .A(n_838), .B(n_842), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_831), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_829), .Y(n_948) );
INVx4_ASAP7_75t_L g949 ( .A(n_841), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_776), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_776), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_776), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_798), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_829), .B(n_870), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_829), .Y(n_955) );
OA21x2_ASAP7_75t_L g956 ( .A1(n_814), .A2(n_807), .B(n_871), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_860), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_836), .B(n_843), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_860), .Y(n_959) );
OR2x6_ASAP7_75t_L g960 ( .A(n_832), .B(n_837), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_836), .B(n_860), .Y(n_961) );
BUFx8_ASAP7_75t_SL g962 ( .A(n_833), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_852), .B(n_825), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_826), .B(n_857), .Y(n_964) );
AO21x2_ASAP7_75t_L g965 ( .A1(n_853), .A2(n_883), .B(n_793), .Y(n_965) );
OR2x6_ASAP7_75t_L g966 ( .A(n_799), .B(n_784), .Y(n_966) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_866), .Y(n_967) );
OR2x2_ASAP7_75t_L g968 ( .A(n_794), .B(n_791), .Y(n_968) );
OR2x6_ASAP7_75t_L g969 ( .A(n_799), .B(n_784), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_801), .B(n_802), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_780), .Y(n_971) );
INVx3_ASAP7_75t_L g972 ( .A(n_879), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_801), .B(n_802), .Y(n_973) );
INVx2_ASAP7_75t_L g974 ( .A(n_801), .Y(n_974) );
INVx3_ASAP7_75t_L g975 ( .A(n_879), .Y(n_975) );
INVxp67_ASAP7_75t_L g976 ( .A(n_791), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_933), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_916), .Y(n_978) );
INVx4_ASAP7_75t_L g979 ( .A(n_925), .Y(n_979) );
NAND2x1_ASAP7_75t_L g980 ( .A(n_925), .B(n_966), .Y(n_980) );
INVx5_ASAP7_75t_L g981 ( .A(n_925), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_970), .B(n_973), .Y(n_982) );
AND2x4_ASAP7_75t_SL g983 ( .A(n_925), .B(n_966), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_970), .B(n_973), .Y(n_984) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_962), .Y(n_985) );
INVx4_ASAP7_75t_L g986 ( .A(n_966), .Y(n_986) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_968), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_935), .Y(n_988) );
INVx5_ASAP7_75t_SL g989 ( .A(n_966), .Y(n_989) );
AND2x4_ASAP7_75t_L g990 ( .A(n_955), .B(n_957), .Y(n_990) );
OR2x2_ASAP7_75t_L g991 ( .A(n_969), .B(n_895), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_898), .Y(n_992) );
BUFx2_ASAP7_75t_L g993 ( .A(n_969), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_905), .Y(n_994) );
NOR2x1_ASAP7_75t_SL g995 ( .A(n_969), .B(n_960), .Y(n_995) );
BUFx2_ASAP7_75t_L g996 ( .A(n_969), .Y(n_996) );
NOR2x1_ASAP7_75t_SL g997 ( .A(n_960), .B(n_949), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_906), .Y(n_998) );
BUFx3_ASAP7_75t_L g999 ( .A(n_889), .Y(n_999) );
INVx1_ASAP7_75t_SL g1000 ( .A(n_945), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_915), .B(n_899), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_908), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_936), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_895), .B(n_967), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_889), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_939), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_892), .Y(n_1007) );
AND2x4_ASAP7_75t_L g1008 ( .A(n_957), .B(n_959), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_891), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_976), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_961), .A2(n_901), .B1(n_923), .B2(n_958), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_974), .B(n_888), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_888), .B(n_890), .Y(n_1013) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_948), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_888), .B(n_890), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_897), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_897), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_900), .B(n_950), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_921), .B(n_929), .Y(n_1019) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_954), .B(n_948), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_904), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_971), .Y(n_1022) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_921), .Y(n_1023) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_896), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_929), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_937), .B(n_938), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_951), .B(n_952), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_964), .B(n_904), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_964), .Y(n_1029) );
INVx4_ASAP7_75t_L g1030 ( .A(n_949), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_903), .A2(n_930), .B1(n_931), .B2(n_918), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_913), .B(n_911), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_907), .B(n_922), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_907), .B(n_922), .Y(n_1034) );
INVx4_ASAP7_75t_L g1035 ( .A(n_949), .Y(n_1035) );
INVxp67_ASAP7_75t_L g1036 ( .A(n_940), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_912), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_907), .B(n_922), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_946), .B(n_920), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_927), .B(n_975), .Y(n_1040) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_926), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_972), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1018), .B(n_894), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_992), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1018), .B(n_894), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_982), .B(n_919), .Y(n_1046) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_1004), .B(n_902), .Y(n_1047) );
BUFx2_ASAP7_75t_L g1048 ( .A(n_1014), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_982), .B(n_919), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_1028), .B(n_893), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_977), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_994), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_988), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_984), .B(n_953), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_998), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1013), .B(n_919), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_1039), .B(n_917), .Y(n_1057) );
NOR2xp33_ASAP7_75t_L g1058 ( .A(n_1009), .B(n_1000), .Y(n_1058) );
INVx2_ASAP7_75t_SL g1059 ( .A(n_1014), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_1013), .B(n_893), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1002), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1015), .B(n_963), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1063 ( .A(n_1036), .B(n_965), .Y(n_1063) );
OR2x2_ASAP7_75t_L g1064 ( .A(n_1024), .B(n_928), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1015), .B(n_963), .Y(n_1065) );
INVx4_ASAP7_75t_L g1066 ( .A(n_1030), .Y(n_1066) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_1020), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1022), .Y(n_1068) );
NAND2xp5_ASAP7_75t_SL g1069 ( .A(n_1030), .B(n_942), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1037), .B(n_910), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1003), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1006), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1012), .B(n_932), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1001), .B(n_934), .Y(n_1074) );
NOR2xp33_ASAP7_75t_L g1075 ( .A(n_987), .B(n_891), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1028), .B(n_924), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_1019), .B(n_941), .Y(n_1077) );
INVx2_ASAP7_75t_L g1078 ( .A(n_978), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1031), .B(n_934), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_1023), .Y(n_1080) );
OR2x2_ASAP7_75t_L g1081 ( .A(n_1019), .B(n_941), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1006), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1010), .B(n_934), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1029), .B(n_947), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1029), .B(n_947), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_1027), .B(n_943), .Y(n_1086) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_1026), .B(n_942), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1060), .B(n_1033), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1044), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1052), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_1078), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1092 ( .A(n_1050), .B(n_990), .Y(n_1092) );
NOR2xp33_ASAP7_75t_L g1093 ( .A(n_1063), .B(n_909), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1056), .B(n_1034), .Y(n_1094) );
NOR2xp67_ASAP7_75t_SL g1095 ( .A(n_1066), .B(n_999), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1055), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1046), .B(n_1038), .Y(n_1097) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1061), .Y(n_1098) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1050), .B(n_1008), .Y(n_1099) );
AND2x4_ASAP7_75t_L g1100 ( .A(n_1050), .B(n_1008), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_1080), .B(n_1011), .Y(n_1101) );
NOR2xp33_ASAP7_75t_L g1102 ( .A(n_1083), .B(n_1040), .Y(n_1102) );
NOR2xp33_ASAP7_75t_SL g1103 ( .A(n_1066), .B(n_985), .Y(n_1103) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1043), .B(n_1008), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1049), .B(n_1062), .Y(n_1105) );
INVx1_ASAP7_75t_SL g1106 ( .A(n_1058), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1068), .B(n_1025), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1049), .B(n_1062), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1054), .B(n_1032), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1065), .B(n_1027), .Y(n_1110) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_1067), .Y(n_1111) );
NOR2xp33_ASAP7_75t_L g1112 ( .A(n_1079), .B(n_1040), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1047), .B(n_991), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_1047), .B(n_1021), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1045), .B(n_1007), .Y(n_1115) );
INVx2_ASAP7_75t_L g1116 ( .A(n_1091), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1117 ( .A1(n_1103), .A2(n_1069), .B(n_997), .Y(n_1117) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_1093), .B(n_1075), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1089), .Y(n_1119) );
AOI21xp33_ASAP7_75t_L g1120 ( .A1(n_1101), .A2(n_980), .B(n_1064), .Y(n_1120) );
INVxp67_ASAP7_75t_L g1121 ( .A(n_1111), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1105), .B(n_1084), .Y(n_1122) );
CKINVDCx16_ASAP7_75t_R g1123 ( .A(n_1106), .Y(n_1123) );
AND2x4_ASAP7_75t_L g1124 ( .A(n_1092), .B(n_1048), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1108), .B(n_1084), .Y(n_1125) );
NAND2xp33_ASAP7_75t_SL g1126 ( .A(n_1095), .B(n_980), .Y(n_1126) );
OAI222xp33_ASAP7_75t_L g1127 ( .A1(n_1110), .A2(n_979), .B1(n_986), .B2(n_996), .C1(n_993), .C2(n_1059), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1090), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1108), .B(n_1085), .Y(n_1129) );
AOI21xp33_ASAP7_75t_L g1130 ( .A1(n_1107), .A2(n_1064), .B(n_1077), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1088), .B(n_1086), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1088), .B(n_1086), .Y(n_1132) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1091), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1096), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1098), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_1097), .B(n_1077), .Y(n_1136) );
INVxp67_ASAP7_75t_SL g1137 ( .A(n_1121), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1116), .Y(n_1138) );
HB1xp67_ASAP7_75t_L g1139 ( .A(n_1121), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1116), .Y(n_1140) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_1123), .A2(n_983), .B1(n_995), .B2(n_997), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1119), .Y(n_1142) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1128), .Y(n_1143) );
AO21x1_ASAP7_75t_L g1144 ( .A1(n_1126), .A2(n_979), .B(n_986), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1134), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1135), .Y(n_1146) );
AOI222xp33_ASAP7_75t_L g1147 ( .A1(n_1118), .A2(n_1112), .B1(n_1102), .B2(n_1057), .C1(n_1070), .C2(n_1094), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1136), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1133), .Y(n_1149) );
AOI21xp5_ASAP7_75t_L g1150 ( .A1(n_1144), .A2(n_1117), .B(n_1127), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1142), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1143), .Y(n_1152) );
AOI322xp5_ASAP7_75t_L g1153 ( .A1(n_1148), .A2(n_1132), .A3(n_1131), .B1(n_1125), .B2(n_1122), .C1(n_1129), .C2(n_1094), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1154 ( .A1(n_1141), .A2(n_1124), .B1(n_979), .B2(n_1104), .Y(n_1154) );
AOI22x1_ASAP7_75t_L g1155 ( .A1(n_1139), .A2(n_1035), .B1(n_1005), .B2(n_1104), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1145), .Y(n_1156) );
OAI31xp33_ASAP7_75t_L g1157 ( .A1(n_1139), .A2(n_1120), .A3(n_1130), .B(n_1092), .Y(n_1157) );
INVxp67_ASAP7_75t_L g1158 ( .A(n_1137), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1146), .Y(n_1159) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_1147), .A2(n_1102), .B1(n_1115), .B2(n_1100), .Y(n_1160) );
NAND3xp33_ASAP7_75t_SL g1161 ( .A(n_1150), .B(n_1035), .C(n_1081), .Y(n_1161) );
AOI211xp5_ASAP7_75t_SL g1162 ( .A1(n_1154), .A2(n_914), .B(n_941), .C(n_1087), .Y(n_1162) );
AOI221xp5_ASAP7_75t_L g1163 ( .A1(n_1158), .A2(n_1138), .B1(n_1140), .B2(n_1149), .C(n_1109), .Y(n_1163) );
AND3x1_ASAP7_75t_L g1164 ( .A(n_1157), .B(n_1005), .C(n_1140), .Y(n_1164) );
NOR3xp33_ASAP7_75t_L g1165 ( .A(n_1151), .B(n_1035), .C(n_944), .Y(n_1165) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_1153), .B(n_1016), .C(n_1017), .Y(n_1166) );
OAI221xp5_ASAP7_75t_L g1167 ( .A1(n_1164), .A2(n_1160), .B1(n_1155), .B2(n_1156), .C(n_1159), .Y(n_1167) );
NOR2x1_ASAP7_75t_L g1168 ( .A(n_1161), .B(n_1152), .Y(n_1168) );
OAI211xp5_ASAP7_75t_SL g1169 ( .A1(n_1162), .A2(n_1113), .B(n_1081), .C(n_1074), .Y(n_1169) );
NAND5xp2_ASAP7_75t_L g1170 ( .A(n_1165), .B(n_1073), .C(n_1076), .D(n_989), .E(n_1085), .Y(n_1170) );
NOR3xp33_ASAP7_75t_L g1171 ( .A(n_1167), .B(n_1166), .C(n_1163), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1168), .Y(n_1172) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1169), .Y(n_1173) );
NOR4xp25_ASAP7_75t_L g1174 ( .A(n_1170), .B(n_1051), .C(n_1071), .D(n_1072), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1175 ( .A(n_1172), .Y(n_1175) );
INVx4_ASAP7_75t_L g1176 ( .A(n_1173), .Y(n_1176) );
AO22x2_ASAP7_75t_L g1177 ( .A1(n_1176), .A2(n_1171), .B1(n_1174), .B2(n_1100), .Y(n_1177) );
OAI22x1_ASAP7_75t_L g1178 ( .A1(n_1175), .A2(n_981), .B1(n_956), .B2(n_1099), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1177), .Y(n_1179) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1178), .Y(n_1180) );
OAI22xp5_ASAP7_75t_L g1181 ( .A1(n_1179), .A2(n_989), .B1(n_1114), .B2(n_1042), .Y(n_1181) );
OAI22xp33_ASAP7_75t_L g1182 ( .A1(n_1180), .A2(n_960), .B1(n_956), .B2(n_1041), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1181), .B(n_1182), .Y(n_1183) );
AO21x2_ASAP7_75t_L g1184 ( .A1(n_1183), .A2(n_1072), .B(n_1071), .Y(n_1184) );
AOI21xp5_ASAP7_75t_L g1185 ( .A1(n_1184), .A2(n_1053), .B(n_1082), .Y(n_1185) );
endmodule