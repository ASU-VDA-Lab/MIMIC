module fake_jpeg_2726_n_150 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_29),
.Y(n_59)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_45),
.Y(n_64)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_11),
.B1(n_17),
.B2(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_2),
.C(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_50),
.Y(n_65)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_16),
.B(n_26),
.Y(n_50)
);

CKINVDCx9p33_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_55),
.B(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_11),
.B1(n_17),
.B2(n_21),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_35),
.B1(n_42),
.B2(n_29),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_27),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_14),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_31),
.A2(n_23),
.B1(n_14),
.B2(n_6),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_63),
.B1(n_70),
.B2(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_41),
.B(n_6),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_29),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_89),
.B1(n_63),
.B2(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_95),
.Y(n_104)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_74),
.B(n_66),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_67),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_105),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_90),
.B1(n_92),
.B2(n_84),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_76),
.C(n_59),
.Y(n_110)
);

OR2x4_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_70),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_83),
.B(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_54),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_54),
.B1(n_66),
.B2(n_74),
.Y(n_115)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_83),
.B(n_86),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_118),
.C(n_122),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_98),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_124),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_104),
.B(n_111),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_129),
.C(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_130),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_108),
.B(n_105),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_106),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_108),
.B(n_125),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_132),
.B(n_109),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_113),
.B1(n_117),
.B2(n_122),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_132),
.B1(n_107),
.B2(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_115),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_125),
.B1(n_106),
.B2(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_141),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_142),
.B(n_138),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_103),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_140),
.B(n_107),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_147),
.B1(n_144),
.B2(n_103),
.Y(n_148)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_81),
.B(n_94),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_54),
.Y(n_150)
);


endmodule