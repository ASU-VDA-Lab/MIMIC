module fake_jpeg_10722_n_628 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_628);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_628;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_30),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_61),
.B(n_62),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_7),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_19),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_68),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_30),
.B(n_11),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_74),
.B(n_78),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_76),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_36),
.B(n_37),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_82),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_84),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_87),
.Y(n_144)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_11),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_89),
.B(n_94),
.Y(n_209)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_15),
.C(n_14),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_16),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_97),
.B(n_13),
.Y(n_167)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_123),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_20),
.Y(n_112)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_20),
.Y(n_115)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_25),
.Y(n_118)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_48),
.Y(n_120)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_121),
.Y(n_132)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_21),
.B(n_15),
.Y(n_123)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_25),
.Y(n_124)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_25),
.Y(n_126)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_79),
.A2(n_51),
.B1(n_56),
.B2(n_38),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_131),
.A2(n_178),
.B1(n_197),
.B2(n_47),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_89),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_135),
.B(n_151),
.Y(n_271)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_146),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_126),
.B1(n_125),
.B2(n_82),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_148),
.A2(n_179),
.B1(n_46),
.B2(n_42),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_100),
.B(n_41),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_157),
.Y(n_240)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_162),
.Y(n_251)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_164),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_167),
.B(n_180),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_62),
.B(n_52),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_22),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_65),
.A2(n_38),
.B1(n_56),
.B2(n_43),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_174),
.A2(n_41),
.B1(n_39),
.B2(n_22),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_79),
.A2(n_51),
.B1(n_56),
.B2(n_38),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_67),
.A2(n_43),
.B1(n_57),
.B2(n_42),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_94),
.B(n_23),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_70),
.B(n_23),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_185),
.B(n_0),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_72),
.A2(n_43),
.B1(n_58),
.B2(n_40),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_73),
.Y(n_199)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_75),
.Y(n_201)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_201),
.Y(n_278)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_77),
.Y(n_206)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_210),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_211),
.B(n_222),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_174),
.B1(n_154),
.B2(n_209),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_212),
.A2(n_220),
.B1(n_235),
.B2(n_237),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_138),
.B(n_58),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_214),
.B(n_224),
.Y(n_325)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_127),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_215),
.Y(n_334)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_216),
.Y(n_320)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_217),
.Y(n_326)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_218),
.Y(n_311)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_186),
.A2(n_81),
.B1(n_117),
.B2(n_111),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_154),
.B(n_173),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_221),
.B(n_247),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_128),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_129),
.B(n_55),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_145),
.Y(n_226)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_226),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_179),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_227),
.B(n_236),
.Y(n_295)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_228),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_140),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_145),
.Y(n_231)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_233),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_83),
.B1(n_87),
.B2(n_91),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_234),
.A2(n_244),
.B1(n_245),
.B2(n_203),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_131),
.A2(n_107),
.B1(n_101),
.B2(n_118),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_196),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_178),
.A2(n_68),
.B1(n_24),
.B2(n_40),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_149),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g323 ( 
.A(n_238),
.Y(n_323)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_243),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_152),
.A2(n_166),
.B1(n_184),
.B2(n_195),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_246),
.B(n_248),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_84),
.B(n_24),
.C(n_55),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_148),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_197),
.A2(n_200),
.B(n_160),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_249),
.A2(n_189),
.B(n_136),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_143),
.A2(n_57),
.B1(n_46),
.B2(n_35),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_250),
.A2(n_279),
.B1(n_278),
.B2(n_270),
.Y(n_336)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_159),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_252),
.B(n_254),
.Y(n_319)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_133),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_153),
.Y(n_255)
);

INVx4_ASAP7_75t_SL g288 ( 
.A(n_255),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_156),
.A2(n_35),
.B1(n_47),
.B2(n_39),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g309 ( 
.A1(n_256),
.A2(n_277),
.B1(n_137),
.B2(n_181),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_258),
.B(n_266),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_263),
.Y(n_328)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_155),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_260),
.B(n_261),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_193),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_172),
.Y(n_262)
);

INVx5_ASAP7_75t_SL g324 ( 
.A(n_262),
.Y(n_324)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_265),
.A2(n_273),
.B1(n_275),
.B2(n_1),
.Y(n_310)
);

AOI32xp33_ASAP7_75t_L g266 ( 
.A1(n_132),
.A2(n_47),
.A3(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_193),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_268),
.Y(n_298)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_177),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_269),
.Y(n_297)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_187),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_272),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_134),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_274),
.Y(n_333)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_194),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_132),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_276),
.Y(n_301)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_208),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_163),
.B(n_12),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_3),
.C(n_4),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_141),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_280),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_130),
.B(n_0),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_170),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_282),
.A2(n_144),
.B1(n_192),
.B2(n_190),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_283),
.A2(n_237),
.B1(n_249),
.B2(n_265),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_188),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_285),
.B(n_287),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_191),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_290),
.B(n_316),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_192),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_294),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_220),
.B(n_190),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_244),
.A2(n_189),
.B1(n_176),
.B2(n_163),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_299),
.A2(n_331),
.B1(n_232),
.B2(n_280),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_304),
.A2(n_275),
.B(n_239),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_309),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_171),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_308),
.B(n_322),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g361 ( 
.A1(n_310),
.A2(n_336),
.B1(n_243),
.B2(n_238),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_245),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_SL g318 ( 
.A(n_281),
.B(n_5),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_318),
.A2(n_274),
.B(n_230),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_273),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_229),
.B(n_1),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_225),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_214),
.A2(n_221),
.B1(n_256),
.B2(n_235),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_250),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_337),
.B(n_340),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_267),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_302),
.Y(n_341)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_361),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_337),
.A2(n_234),
.B1(n_233),
.B2(n_215),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_345),
.A2(n_370),
.B1(n_381),
.B2(n_342),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_335),
.A2(n_285),
.B1(n_293),
.B2(n_294),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_346),
.A2(n_351),
.B1(n_382),
.B2(n_344),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_289),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_356),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_293),
.B(n_322),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_350),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_335),
.A2(n_277),
.B1(n_210),
.B2(n_282),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_353),
.A2(n_384),
.B(n_297),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_354),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_319),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_291),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_365),
.Y(n_395)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_328),
.B(n_271),
.Y(n_362)
);

O2A1O1Ixp33_ASAP7_75t_SL g365 ( 
.A1(n_290),
.A2(n_277),
.B(n_213),
.C(n_218),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_338),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_369),
.Y(n_416)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_320),
.Y(n_368)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_295),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_303),
.A2(n_253),
.B1(n_226),
.B2(n_231),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_371),
.B(n_377),
.Y(n_410)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_328),
.B(n_301),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_373),
.B(n_379),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_304),
.B(n_251),
.C(n_257),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_383),
.C(n_385),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_324),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_376),
.Y(n_420)
);

AND2x2_ASAP7_75t_SL g377 ( 
.A(n_308),
.B(n_262),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_316),
.A2(n_272),
.B1(n_255),
.B2(n_3),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_324),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_328),
.A2(n_283),
.B1(n_317),
.B2(n_309),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_317),
.A2(n_309),
.B1(n_325),
.B2(n_301),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_306),
.B(n_292),
.C(n_297),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_318),
.A2(n_298),
.B(n_340),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g385 ( 
.A(n_327),
.B(n_309),
.C(n_306),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_358),
.B(n_292),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_390),
.B(n_393),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_373),
.B(n_307),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_364),
.B(n_348),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_418),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_397),
.A2(n_411),
.B1(n_414),
.B2(n_419),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_400),
.A2(n_377),
.B1(n_365),
.B2(n_355),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_353),
.A2(n_284),
.B(n_312),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_401),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_344),
.A2(n_296),
.B1(n_330),
.B2(n_286),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_404),
.A2(n_370),
.B1(n_345),
.B2(n_360),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_346),
.A2(n_296),
.B1(n_334),
.B2(n_330),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_352),
.A2(n_334),
.B1(n_312),
.B2(n_286),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_412),
.A2(n_421),
.B1(n_379),
.B2(n_376),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_344),
.A2(n_315),
.B1(n_311),
.B2(n_332),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_415),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_363),
.A2(n_311),
.B(n_323),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_352),
.A2(n_315),
.B1(n_313),
.B2(n_329),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_381),
.A2(n_339),
.B1(n_313),
.B2(n_329),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_363),
.A2(n_314),
.B(n_284),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_401),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_369),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_429),
.C(n_456),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_426),
.A2(n_427),
.B1(n_441),
.B2(n_457),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_382),
.B1(n_348),
.B2(n_364),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_349),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_428),
.B(n_434),
.C(n_438),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_347),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_386),
.Y(n_430)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_430),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_416),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_447),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_432),
.A2(n_445),
.B1(n_450),
.B2(n_451),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_371),
.C(n_383),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_448),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_385),
.C(n_374),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_366),
.Y(n_439)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_406),
.B(n_367),
.Y(n_442)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_442),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_397),
.A2(n_385),
.B1(n_362),
.B2(n_365),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_446),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_416),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_388),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_375),
.C(n_377),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_390),
.C(n_388),
.Y(n_464)
);

OAI22x1_ASAP7_75t_SL g450 ( 
.A1(n_404),
.A2(n_377),
.B1(n_384),
.B2(n_343),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_395),
.A2(n_375),
.B1(n_359),
.B2(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_398),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_350),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_454),
.Y(n_458)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_402),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_403),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_389),
.B(n_380),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_395),
.A2(n_354),
.B1(n_372),
.B2(n_368),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_438),
.B(n_410),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_459),
.B(n_457),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_410),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_462),
.B(n_485),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_464),
.B(n_477),
.C(n_451),
.Y(n_502)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_424),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_465),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_425),
.A2(n_392),
.B(n_387),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_467),
.A2(n_482),
.B(n_450),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_429),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_479),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_427),
.A2(n_411),
.B1(n_414),
.B2(n_399),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_472),
.A2(n_478),
.B1(n_488),
.B2(n_444),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_449),
.C(n_431),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_441),
.A2(n_399),
.B1(n_389),
.B2(n_419),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_454),
.Y(n_479)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_481),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_433),
.A2(n_405),
.B(n_418),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_447),
.Y(n_483)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_393),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_442),
.A2(n_413),
.B1(n_417),
.B2(n_422),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_486),
.A2(n_487),
.B1(n_448),
.B2(n_435),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_439),
.A2(n_422),
.B1(n_403),
.B2(n_415),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_426),
.A2(n_405),
.B1(n_421),
.B2(n_412),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_490),
.A2(n_513),
.B1(n_432),
.B2(n_476),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_473),
.A2(n_437),
.B(n_435),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_491),
.A2(n_517),
.B(n_518),
.Y(n_539)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_475),
.Y(n_493)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_493),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_477),
.B(n_456),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_494),
.B(n_501),
.Y(n_544)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_475),
.Y(n_495)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_495),
.Y(n_529)
);

INVx13_ASAP7_75t_L g496 ( 
.A(n_466),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_471),
.B(n_470),
.Y(n_497)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_498),
.A2(n_458),
.B1(n_479),
.B2(n_482),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_473),
.Y(n_500)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_500),
.Y(n_542)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_480),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_502),
.B(n_510),
.C(n_467),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_461),
.B(n_443),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_511),
.Y(n_538)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_480),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_505),
.A2(n_506),
.B1(n_515),
.B2(n_489),
.Y(n_525)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_460),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_464),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_509),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_474),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_458),
.B(n_423),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_459),
.B(n_450),
.C(n_444),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g511 ( 
.A(n_469),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_512),
.A2(n_402),
.B(n_408),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_474),
.A2(n_443),
.B1(n_405),
.B2(n_455),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_460),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_462),
.B(n_405),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_516),
.B(n_423),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_485),
.B(n_453),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_478),
.B(n_452),
.Y(n_518)
);

XOR2x2_ASAP7_75t_L g546 ( 
.A(n_521),
.B(n_540),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_522),
.A2(n_530),
.B1(n_495),
.B2(n_493),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_526),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_525),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_463),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_498),
.A2(n_470),
.B1(n_483),
.B2(n_484),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_528),
.B(n_530),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_500),
.A2(n_483),
.B1(n_472),
.B2(n_488),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_489),
.C(n_484),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_531),
.B(n_537),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_532),
.A2(n_501),
.B1(n_505),
.B2(n_499),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_514),
.B(n_476),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_533),
.B(n_534),
.C(n_516),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_468),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_513),
.A2(n_468),
.B1(n_446),
.B2(n_440),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_536),
.A2(n_515),
.B1(n_506),
.B2(n_503),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_502),
.B(n_436),
.C(n_430),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_541),
.A2(n_499),
.B(n_509),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_508),
.B(n_409),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_492),
.Y(n_563)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_535),
.Y(n_545)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_545),
.Y(n_571)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_542),
.Y(n_547)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_547),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_548),
.A2(n_562),
.B1(n_521),
.B2(n_520),
.Y(n_580)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_550),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_541),
.A2(n_512),
.B(n_491),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_551),
.A2(n_555),
.B(n_549),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_538),
.B(n_497),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_553),
.A2(n_531),
.B1(n_539),
.B2(n_529),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_558),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_555),
.B(n_556),
.Y(n_582)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_536),
.Y(n_556)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_544),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_557),
.B(n_523),
.Y(n_566)
);

CKINVDCx12_ASAP7_75t_R g560 ( 
.A(n_524),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_560),
.Y(n_575)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_527),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_561),
.B(n_520),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_563),
.B(n_523),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_537),
.B(n_492),
.C(n_519),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_564),
.B(n_519),
.C(n_540),
.Y(n_574)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_565),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_566),
.B(n_408),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g567 ( 
.A1(n_548),
.A2(n_522),
.B(n_532),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_567),
.B(n_576),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_569),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_572),
.A2(n_561),
.B(n_409),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_534),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_573),
.B(n_574),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_SL g576 ( 
.A(n_554),
.B(n_543),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_559),
.B(n_526),
.C(n_533),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_579),
.B(n_581),
.C(n_552),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_580),
.B(n_562),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_552),
.B(n_546),
.C(n_556),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_583),
.B(n_587),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_581),
.A2(n_551),
.B(n_545),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_585),
.A2(n_589),
.B(n_496),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_575),
.B(n_570),
.C(n_574),
.Y(n_587)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_588),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_582),
.A2(n_550),
.B(n_549),
.Y(n_589)
);

AOI21x1_ASAP7_75t_L g590 ( 
.A1(n_573),
.A2(n_553),
.B(n_547),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_590),
.A2(n_593),
.B(n_589),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_568),
.B(n_546),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_591),
.B(n_594),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_578),
.A2(n_571),
.B1(n_577),
.B2(n_567),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_SL g606 ( 
.A(n_596),
.B(n_407),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_570),
.C(n_579),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_597),
.A2(n_602),
.B(n_591),
.Y(n_611)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_599),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_584),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_588),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_576),
.C(n_580),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_595),
.B(n_567),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_603),
.B(n_605),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_604),
.A2(n_593),
.B(n_592),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_586),
.Y(n_605)
);

XNOR2x1_ASAP7_75t_L g614 ( 
.A(n_606),
.B(n_288),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_609),
.B(n_610),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_611),
.A2(n_613),
.B(n_607),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_601),
.A2(n_586),
.B(n_407),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_612),
.B(n_614),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_598),
.A2(n_600),
.B(n_605),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_617),
.B(n_618),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_608),
.A2(n_333),
.B1(n_314),
.B2(n_288),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_615),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_619),
.B(n_326),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_622),
.B(n_620),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_623),
.B(n_621),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_624),
.B(n_616),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_625),
.A2(n_618),
.B(n_339),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_SL g627 ( 
.A1(n_626),
.A2(n_288),
.B(n_323),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_627),
.A2(n_323),
.B(n_424),
.Y(n_628)
);


endmodule