module fake_jpeg_22500_n_136 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_29),
.Y(n_30)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_17),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_12),
.B1(n_16),
.B2(n_18),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_12),
.B1(n_25),
.B2(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_45),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_46),
.B1(n_25),
.B2(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_16),
.B1(n_12),
.B2(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_51),
.B1(n_48),
.B2(n_45),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_28),
.B1(n_33),
.B2(n_39),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_60),
.B1(n_64),
.B2(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_30),
.Y(n_56)
);

BUFx24_ASAP7_75t_SL g69 ( 
.A(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_71),
.Y(n_83)
);

OA21x2_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_35),
.B(n_31),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_75),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_24),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_47),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_80),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_54),
.B(n_57),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_85),
.B(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_82),
.A2(n_87),
.B(n_18),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_88),
.C(n_74),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_19),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_22),
.C(n_63),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_77),
.C(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_76),
.B1(n_66),
.B2(n_22),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_94),
.B1(n_99),
.B2(n_88),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_69),
.B1(n_27),
.B2(n_19),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_15),
.B(n_14),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_98),
.B(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_27),
.B1(n_18),
.B2(n_15),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_107),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_84),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_105),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_96),
.B(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_95),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_93),
.B1(n_97),
.B2(n_77),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_92),
.B1(n_96),
.B2(n_99),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_104),
.B(n_15),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_94),
.Y(n_113)
);

OAI31xp33_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_105),
.A3(n_106),
.B(n_107),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_115),
.B(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_20),
.Y(n_121)
);

OAI321xp33_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_13),
.B1(n_20),
.B2(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_4),
.Y(n_127)
);

NAND4xp25_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_8),
.C(n_9),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_118),
.B(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_7),
.C(n_8),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_129),
.C(n_133),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_9),
.B(n_10),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_SL g136 ( 
.A(n_134),
.B(n_135),
.Y(n_136)
);


endmodule