module fake_jpeg_3491_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_SL g51 ( 
.A(n_49),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_79),
.Y(n_94)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_71),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_76),
.Y(n_87)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_0),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_65),
.B1(n_61),
.B2(n_70),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_80),
.B1(n_77),
.B2(n_60),
.Y(n_100)
);

FAx1_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_70),
.CI(n_61),
.CON(n_82),
.SN(n_82)
);

NAND2x1p5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_78),
.Y(n_103)
);

CKINVDCx9p33_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_61),
.B1(n_60),
.B2(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_76),
.B1(n_63),
.B2(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_87),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_105),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_108),
.B1(n_81),
.B2(n_84),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_67),
.B1(n_62),
.B2(n_56),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_106),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_58),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_68),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_54),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_90),
.B1(n_92),
.B2(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_64),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_110),
.B(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_103),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_35),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_123),
.B1(n_127),
.B2(n_129),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_2),
.Y(n_151)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_88),
.B1(n_59),
.B2(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_108),
.A2(n_59),
.B1(n_55),
.B2(n_57),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_133),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_112),
.C(n_21),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_136),
.C(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_20),
.C(n_44),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_0),
.B(n_1),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_11),
.B(n_12),
.Y(n_173)
);

INVx5_ASAP7_75t_SL g138 ( 
.A(n_121),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_22),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_26),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_145),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_46),
.B1(n_43),
.B2(n_42),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_148),
.B(n_10),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_37),
.C(n_36),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_115),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_154),
.B1(n_5),
.B2(n_7),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_34),
.C(n_32),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_4),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_159),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_136),
.C(n_140),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_162),
.C(n_165),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_123),
.B(n_30),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_172),
.B(n_173),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_29),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_164),
.B1(n_13),
.B2(n_14),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_28),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_170),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_171),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_11),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_18),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_24),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_15),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_176),
.B(n_179),
.Y(n_197)
);

AO22x1_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_138),
.B1(n_144),
.B2(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_169),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_23),
.C(n_17),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_185),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_184),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_168),
.C(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_196),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_183),
.C(n_182),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_201),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_190),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_203),
.B(n_194),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_195),
.C(n_183),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_202),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_197),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_205),
.B1(n_180),
.B2(n_188),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_168),
.Y(n_213)
);


endmodule