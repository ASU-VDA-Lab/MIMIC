module fake_netlist_6_2589_n_4357 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_464, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4357);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_464;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4357;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_700;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3301;
wire n_3089;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_873;
wire n_1285;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_544;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_4308;
wire n_658;
wire n_616;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_3048;
wire n_2729;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_4060;
wire n_943;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_538;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_1441;
wire n_606;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_3446;
wire n_4158;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_586;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_2347;
wire n_690;
wire n_1886;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_2178;
wire n_701;
wire n_3271;
wire n_950;
wire n_4248;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_1767;
wire n_627;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3253;
wire n_3431;
wire n_3337;
wire n_3209;
wire n_3450;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2750;
wire n_2893;
wire n_2558;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4289;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4288;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1714;
wire n_872;
wire n_1139;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4058;
wire n_4103;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3348;
wire n_3229;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2959;
wire n_2494;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3867;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_745;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_1774;
wire n_2354;
wire n_884;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_474;
wire n_811;
wire n_1207;
wire n_683;
wire n_2442;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2581;
wire n_1363;
wire n_2294;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_4053;
wire n_2748;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3944;
wire n_3909;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2301;
wire n_2209;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3724;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_4056;
wire n_1617;
wire n_3260;
wire n_3816;
wire n_3386;
wire n_3370;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_858;
wire n_4149;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_4355;
wire n_501;
wire n_2276;
wire n_960;
wire n_3234;
wire n_956;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4030;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3276;
wire n_3250;
wire n_1934;
wire n_3194;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_4234;
wire n_4304;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_1037;
wire n_1397;
wire n_621;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_710;
wire n_3730;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_4258;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2760;
wire n_1940;
wire n_1979;
wire n_2560;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3988;
wire n_1974;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4135;
wire n_2871;
wire n_4209;
wire n_4279;
wire n_2688;
wire n_3858;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_2310;
wire n_879;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3562;
wire n_3044;
wire n_3381;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_3305;
wire n_2992;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2923;
wire n_489;
wire n_2885;
wire n_2888;
wire n_2793;
wire n_2715;
wire n_2671;
wire n_1804;
wire n_2761;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_4203;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_2949;
wire n_3726;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2814;
wire n_2528;
wire n_2787;
wire n_2969;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_601;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1785;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1114;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_3473;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_611;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2465;
wire n_1112;
wire n_2275;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_2203;
wire n_1945;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_576;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2615;
wire n_2265;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_2744;
wire n_4309;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_839;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_854;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4105;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1362;
wire n_1156;
wire n_4259;
wire n_3123;
wire n_2600;
wire n_984;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_4104;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4346;
wire n_4351;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2844;
wire n_2490;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_4057;
wire n_679;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_640;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_29),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_224),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_19),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_144),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_309),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_230),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_11),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_253),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_147),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_90),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_251),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_319),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_461),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_328),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_236),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_351),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_232),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_288),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_192),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_9),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_116),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_124),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_394),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_294),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_413),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_125),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_154),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_138),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_284),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_248),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_87),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_298),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_30),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_193),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_169),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_279),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_416),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_276),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_53),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_128),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_348),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_279),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_296),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_95),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_240),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_210),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_251),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_52),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_1),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_414),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_412),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_48),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_400),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_452),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_174),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_350),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_222),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_117),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_259),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_235),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_407),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_150),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_323),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_187),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_143),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_300),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_184),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_32),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_374),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_150),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_148),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_33),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_82),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_55),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_111),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_0),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_437),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_202),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_276),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_128),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_409),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_169),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_355),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_143),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_299),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_411),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_94),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_10),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_226),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_125),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_107),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_230),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_62),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_86),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_403),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_12),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_37),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_327),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_39),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_297),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_71),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_235),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_181),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_391),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_62),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_202),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g577 ( 
.A(n_52),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_448),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_433),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_352),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_90),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_395),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_316),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_361),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_167),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_0),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_297),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_70),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_249),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_21),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_231),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_57),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_267),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_22),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_301),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_4),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_100),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_293),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_267),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_379),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_198),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_201),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_290),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_360),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_300),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_50),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_373),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_122),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_463),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_49),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_141),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_175),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_81),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_320),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_207),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_50),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_94),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_226),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_26),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_86),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_110),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_234),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_385),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_344),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_346),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_426),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_61),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_96),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_111),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_317),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_133),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_449),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_200),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_151),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_244),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_256),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_113),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_378),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_454),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_41),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_248),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_25),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_197),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_243),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_159),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_183),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_464),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_271),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_89),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_380),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_28),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_288),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_357),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_382),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_1),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_183),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_264),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_371),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_367),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_204),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_142),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_188),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_353),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_445),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_349),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_204),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_430),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_363),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_347),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_333),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_425),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_456),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_289),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_105),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_201),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_402),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_162),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_185),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_55),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_404),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_122),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_104),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_289),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_261),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_85),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_272),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_338),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_212),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_428),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_64),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_261),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_167),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_137),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_399),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_71),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_182),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_5),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_165),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_468),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_240),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_193),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_92),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_384),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_59),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_5),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_435),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_188),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_383),
.Y(n_708)
);

BUFx5_ASAP7_75t_L g709 ( 
.A(n_144),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_306),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_141),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_356),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_441),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_368),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_218),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_11),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_174),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_88),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_81),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_178),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_422),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_45),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_120),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_218),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_21),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_158),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_58),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_33),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_106),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_250),
.Y(n_730)
);

BUFx8_ASAP7_75t_SL g731 ( 
.A(n_337),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_341),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_329),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_70),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_78),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_262),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_390),
.Y(n_737)
);

CKINVDCx16_ASAP7_75t_R g738 ( 
.A(n_225),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_189),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_121),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_89),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_99),
.Y(n_742)
);

CKINVDCx16_ASAP7_75t_R g743 ( 
.A(n_69),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_110),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_27),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_292),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_317),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_97),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_278),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_309),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_163),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_377),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_292),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_154),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_53),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_67),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_432),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_197),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_466),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_273),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_7),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_263),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_326),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_275),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_69),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_221),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_315),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_238),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_709),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_709),
.Y(n_770)
);

INVxp33_ASAP7_75t_L g771 ( 
.A(n_678),
.Y(n_771)
);

INVxp33_ASAP7_75t_SL g772 ( 
.A(n_704),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_731),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_482),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_709),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_709),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_709),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_483),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_492),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_709),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_709),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_709),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_709),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_680),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_518),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_494),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_588),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_588),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_510),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_588),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_588),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_588),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_519),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_506),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_607),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_588),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_610),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_518),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_610),
.Y(n_799)
);

INVxp33_ASAP7_75t_SL g800 ( 
.A(n_535),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_610),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_610),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_489),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_610),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_520),
.Y(n_805)
);

CKINVDCx20_ASAP7_75t_R g806 ( 
.A(n_533),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_610),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_722),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_489),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_489),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_539),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_722),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_577),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_489),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_481),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_535),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_722),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_722),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_722),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_712),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_547),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_722),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_736),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_736),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_736),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_736),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_696),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_712),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_736),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_736),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_761),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_761),
.Y(n_832)
);

INVxp33_ASAP7_75t_SL g833 ( 
.A(n_696),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_481),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_553),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_761),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_761),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_556),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_761),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_761),
.Y(n_840)
);

BUFx2_ASAP7_75t_SL g841 ( 
.A(n_624),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_487),
.Y(n_842)
);

CKINVDCx16_ASAP7_75t_R g843 ( 
.A(n_577),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_487),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_487),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_504),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_618),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_501),
.Y(n_848)
);

INVxp33_ASAP7_75t_SL g849 ( 
.A(n_470),
.Y(n_849)
);

INVxp33_ASAP7_75t_SL g850 ( 
.A(n_471),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_501),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_504),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_565),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_501),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_526),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_481),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_618),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_548),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_548),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_548),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_605),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_605),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_605),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_634),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_634),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_634),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_716),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_650),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_650),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_716),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_568),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_716),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_650),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_574),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_735),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_735),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_735),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_748),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_748),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_748),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_766),
.Y(n_881)
);

BUFx2_ASAP7_75t_SL g882 ( 
.A(n_624),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_766),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_766),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_738),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_512),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_512),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_561),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_561),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_578),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_649),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_649),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_698),
.Y(n_893)
);

CKINVDCx14_ASAP7_75t_R g894 ( 
.A(n_575),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_698),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_724),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_724),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_740),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_740),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_504),
.Y(n_900)
);

INVxp33_ASAP7_75t_SL g901 ( 
.A(n_472),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_651),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_651),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_526),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_651),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_675),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_675),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_580),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_732),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_675),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_551),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_728),
.Y(n_912)
);

INVxp67_ASAP7_75t_SL g913 ( 
.A(n_732),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_728),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_728),
.Y(n_915)
);

INVxp67_ASAP7_75t_SL g916 ( 
.A(n_732),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_473),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_738),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_834),
.B(n_522),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_847),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_826),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_855),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_800),
.A2(n_743),
.B1(n_765),
.B2(n_527),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_787),
.Y(n_924)
);

OA21x2_ASAP7_75t_L g925 ( 
.A1(n_911),
.A2(n_579),
.B(n_551),
.Y(n_925)
);

OA22x2_ASAP7_75t_SL g926 ( 
.A1(n_820),
.A2(n_828),
.B1(n_475),
.B2(n_477),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_856),
.B(n_522),
.Y(n_927)
);

AND2x2_ASAP7_75t_SL g928 ( 
.A(n_813),
.B(n_551),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_803),
.B(n_654),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_815),
.Y(n_930)
);

OA21x2_ASAP7_75t_L g931 ( 
.A1(n_911),
.A2(n_668),
.B(n_579),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_868),
.B(n_654),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_787),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_827),
.A2(n_743),
.B1(n_542),
.B2(n_596),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_788),
.A2(n_668),
.B(n_579),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_855),
.Y(n_936)
);

BUFx8_ASAP7_75t_L g937 ( 
.A(n_846),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_855),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_815),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_855),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_855),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_904),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_904),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_841),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_869),
.B(n_584),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_904),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_788),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_826),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_904),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_885),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_836),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_790),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_790),
.Y(n_953)
);

BUFx8_ASAP7_75t_SL g954 ( 
.A(n_773),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_904),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_904),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_791),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_803),
.B(n_668),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_918),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_836),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_840),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_770),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_791),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_840),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_792),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_846),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_770),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_780),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_792),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_809),
.B(n_671),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_780),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_774),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_873),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_809),
.B(n_671),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_810),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_796),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_796),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_797),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_873),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_797),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_849),
.B(n_531),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_799),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_SL g983 ( 
.A(n_813),
.B(n_575),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_909),
.B(n_600),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_852),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_810),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_799),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_900),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_769),
.A2(n_671),
.B(n_757),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_852),
.Y(n_990)
);

OA21x2_ASAP7_75t_L g991 ( 
.A1(n_801),
.A2(n_521),
.B(n_485),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_801),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_900),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_802),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_816),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_769),
.B(n_526),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_775),
.A2(n_757),
.B(n_521),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_802),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_850),
.B(n_667),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_804),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_814),
.B(n_485),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_SL g1002 ( 
.A1(n_833),
.A2(n_589),
.B1(n_636),
.B2(n_619),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_804),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_807),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_807),
.Y(n_1005)
);

AND2x2_ASAP7_75t_SL g1006 ( 
.A(n_843),
.B(n_526),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_775),
.A2(n_777),
.B(n_776),
.Y(n_1007)
);

OA21x2_ASAP7_75t_L g1008 ( 
.A1(n_808),
.A2(n_524),
.B(n_523),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_808),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_901),
.B(n_703),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_776),
.A2(n_524),
.B(n_523),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_779),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_842),
.Y(n_1013)
);

INVxp33_ASAP7_75t_SL g1014 ( 
.A(n_786),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_814),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_812),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_812),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_817),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_857),
.B(n_733),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_817),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_841),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_785),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_818),
.B(n_582),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_818),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_819),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_819),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_822),
.Y(n_1027)
);

OAI22x1_ASAP7_75t_L g1028 ( 
.A1(n_798),
.A2(n_571),
.B1(n_629),
.B2(n_499),
.Y(n_1028)
);

OAI22x1_ASAP7_75t_L g1029 ( 
.A1(n_784),
.A2(n_720),
.B1(n_637),
.B2(n_569),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_772),
.A2(n_744),
.B1(n_717),
.B2(n_474),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_913),
.B(n_473),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_822),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_823),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_823),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_843),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_824),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_771),
.A2(n_480),
.B1(n_484),
.B2(n_478),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_824),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_825),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_825),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_842),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_789),
.Y(n_1042)
);

INVx6_ASAP7_75t_L g1043 ( 
.A(n_916),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_882),
.B(n_609),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_930),
.B(n_902),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_988),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_968),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_968),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_968),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_944),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_921),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_989),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_921),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_989),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_989),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_1035),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1007),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_922),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1007),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_981),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1007),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1002),
.A2(n_794),
.B1(n_795),
.B2(n_778),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_944),
.B(n_919),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_1016),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_966),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_921),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_988),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_988),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_948),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_993),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_993),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1043),
.B(n_793),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_1035),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_993),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_966),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_948),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_985),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_962),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_962),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_922),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_985),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_962),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_948),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_997),
.A2(n_1011),
.B(n_933),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_962),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_990),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_967),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_951),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_951),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_967),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_967),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_967),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_924),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_924),
.Y(n_1094)
);

CKINVDCx6p67_ASAP7_75t_R g1095 ( 
.A(n_1012),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_933),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_922),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_947),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_951),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_947),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_952),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_930),
.B(n_902),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_930),
.B(n_903),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_952),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1043),
.B(n_811),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_953),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_953),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_957),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_1016),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_957),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_960),
.Y(n_1111)
);

OAI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1043),
.A2(n_604),
.B1(n_623),
.B2(n_582),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_963),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_960),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_963),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_965),
.Y(n_1116)
);

NAND2xp33_ASAP7_75t_SL g1117 ( 
.A(n_1022),
.B(n_805),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_922),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1016),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_965),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_960),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_961),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_999),
.B(n_835),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_969),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1043),
.B(n_838),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_969),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_922),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1043),
.B(n_853),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_976),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_939),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_922),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_976),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_977),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_977),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_939),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_978),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_990),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_978),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_961),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_961),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_982),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1010),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_939),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_973),
.B(n_874),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_973),
.B(n_890),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_919),
.B(n_903),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_982),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_964),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_SL g1149 ( 
.A(n_1022),
.B(n_806),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_964),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_987),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_987),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_936),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1006),
.A2(n_928),
.B1(n_821),
.B2(n_871),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_920),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_998),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_973),
.B(n_908),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_998),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_936),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1003),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_972),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_964),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_936),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_950),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_959),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1003),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_979),
.B(n_882),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_971),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_927),
.B(n_905),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1012),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1006),
.B(n_733),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1021),
.B(n_894),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_950),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_927),
.B(n_905),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_936),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_971),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1009),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_979),
.B(n_906),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_971),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1009),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_971),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_L g1182 ( 
.A(n_1044),
.B(n_979),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_997),
.A2(n_781),
.B(n_777),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1020),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1020),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1024),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1024),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1006),
.A2(n_763),
.B1(n_626),
.B2(n_632),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_936),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1038),
.Y(n_1190)
);

OA21x2_ASAP7_75t_L g1191 ( 
.A1(n_997),
.A2(n_1011),
.B(n_1038),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_925),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_925),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_980),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_980),
.Y(n_1195)
);

NAND2x1p5_ASAP7_75t_L g1196 ( 
.A(n_1011),
.B(n_604),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_920),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_945),
.B(n_829),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_980),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_925),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1021),
.B(n_1044),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_992),
.A2(n_782),
.B(n_781),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1023),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_995),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_935),
.A2(n_783),
.B(n_782),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_995),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_925),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_925),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_992),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1031),
.B(n_906),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_992),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_931),
.Y(n_1212)
);

OA21x2_ASAP7_75t_L g1213 ( 
.A1(n_994),
.A2(n_783),
.B(n_829),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1031),
.B(n_907),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_929),
.B(n_907),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_931),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_945),
.B(n_830),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_994),
.A2(n_831),
.B(n_830),
.Y(n_1218)
);

INVx5_ASAP7_75t_L g1219 ( 
.A(n_996),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_931),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_996),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_931),
.Y(n_1222)
);

AND2x2_ASAP7_75t_SL g1223 ( 
.A(n_928),
.B(n_623),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_994),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1012),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_937),
.Y(n_1226)
);

INVxp67_ASAP7_75t_L g1227 ( 
.A(n_983),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_984),
.B(n_831),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_931),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1001),
.Y(n_1230)
);

OA21x2_ASAP7_75t_L g1231 ( 
.A1(n_1000),
.A2(n_837),
.B(n_832),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1001),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1001),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1001),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_984),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_932),
.B(n_832),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_958),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1000),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_958),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_958),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_936),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1000),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_958),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_932),
.B(n_837),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_970),
.Y(n_1245)
);

NAND2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1019),
.B(n_488),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_970),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_940),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_928),
.B(n_910),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_970),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_940),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_983),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_970),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1004),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1004),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_974),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_937),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1037),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_974),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_974),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_974),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1004),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1014),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1029),
.B(n_490),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1023),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1023),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1005),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_940),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1023),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_975),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_929),
.B(n_839),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1050),
.B(n_1037),
.Y(n_1272)
);

AND2x2_ASAP7_75t_SL g1273 ( 
.A(n_1223),
.B(n_526),
.Y(n_1273)
);

NOR3xp33_ASAP7_75t_L g1274 ( 
.A(n_1060),
.B(n_934),
.C(n_1002),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1063),
.B(n_937),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1130),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1203),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1237),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1202),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1218),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1237),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1202),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1063),
.B(n_937),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1142),
.B(n_1042),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1045),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1239),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1201),
.A2(n_1042),
.B1(n_1030),
.B2(n_614),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1164),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1218),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1239),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1202),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1218),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1218),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1045),
.Y(n_1294)
);

AND2x6_ASAP7_75t_L g1295 ( 
.A(n_1192),
.B(n_625),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1240),
.Y(n_1296)
);

AND2x2_ASAP7_75t_SL g1297 ( 
.A(n_1223),
.B(n_526),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1235),
.B(n_929),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1258),
.A2(n_1030),
.B1(n_923),
.B2(n_1042),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1202),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1231),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1240),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1243),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1045),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1243),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1231),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1203),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1198),
.B(n_929),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1217),
.B(n_991),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1245),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1249),
.A2(n_991),
.B1(n_1008),
.B2(n_935),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1228),
.B(n_991),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1231),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1130),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1245),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1188),
.A2(n_923),
.B1(n_934),
.B2(n_672),
.Y(n_1316)
);

BUFx10_ASAP7_75t_L g1317 ( 
.A(n_1172),
.Y(n_1317)
);

NAND2xp33_ASAP7_75t_SL g1318 ( 
.A(n_1171),
.B(n_1029),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1249),
.B(n_708),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1081),
.B(n_1028),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1137),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1247),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1265),
.B(n_708),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1231),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1197),
.B(n_1028),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1067),
.B(n_1068),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1247),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1123),
.B(n_530),
.Y(n_1328)
);

AND2x6_ASAP7_75t_L g1329 ( 
.A(n_1192),
.B(n_625),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1213),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1095),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1086),
.B(n_910),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1213),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1213),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1135),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1067),
.B(n_991),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1213),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1135),
.B(n_672),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1250),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1250),
.Y(n_1340)
);

AND2x6_ASAP7_75t_L g1341 ( 
.A(n_1193),
.B(n_687),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1253),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1253),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1265),
.A2(n_694),
.B1(n_714),
.B2(n_687),
.Y(n_1344)
);

AND3x2_ASAP7_75t_L g1345 ( 
.A(n_1226),
.B(n_612),
.C(n_476),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1143),
.B(n_491),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1068),
.B(n_1008),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1164),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1097),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1070),
.B(n_1008),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1173),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1143),
.B(n_493),
.Y(n_1352)
);

BUFx10_ASAP7_75t_L g1353 ( 
.A(n_1161),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1072),
.B(n_495),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1266),
.B(n_708),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1256),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1256),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1086),
.B(n_912),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1105),
.B(n_1125),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1128),
.B(n_496),
.Y(n_1360)
);

NAND2xp33_ASAP7_75t_L g1361 ( 
.A(n_1057),
.B(n_708),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1266),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1078),
.A2(n_991),
.B1(n_1008),
.B2(n_935),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1065),
.B(n_912),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1259),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1259),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1260),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1269),
.B(n_708),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1146),
.B(n_914),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1260),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1070),
.B(n_1008),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1269),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1261),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1215),
.B(n_694),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1173),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1102),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1146),
.B(n_914),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1261),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_SL g1379 ( 
.A(n_1078),
.B(n_708),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1071),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1079),
.A2(n_935),
.B1(n_996),
.B2(n_721),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1205),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1205),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1227),
.B(n_497),
.Y(n_1384)
);

INVx4_ASAP7_75t_SL g1385 ( 
.A(n_1057),
.Y(n_1385)
);

INVx4_ASAP7_75t_SL g1386 ( 
.A(n_1059),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1071),
.B(n_975),
.Y(n_1387)
);

AND2x6_ASAP7_75t_L g1388 ( 
.A(n_1193),
.B(n_714),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1056),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1074),
.B(n_975),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1252),
.B(n_498),
.Y(n_1391)
);

NOR2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1095),
.B(n_500),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1074),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1052),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1102),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1093),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1046),
.Y(n_1397)
);

AO22x2_ASAP7_75t_L g1398 ( 
.A1(n_1210),
.A2(n_926),
.B1(n_721),
.B2(n_476),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1215),
.B(n_915),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1230),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1210),
.A2(n_639),
.B1(n_647),
.B2(n_638),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1075),
.B(n_915),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1230),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1079),
.A2(n_935),
.B1(n_996),
.B2(n_986),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1102),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1082),
.B(n_975),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1232),
.Y(n_1407)
);

AND2x6_ASAP7_75t_L g1408 ( 
.A(n_1200),
.B(n_475),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1082),
.B(n_975),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1144),
.B(n_502),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1097),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1052),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1232),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1233),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1233),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1161),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1056),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1085),
.B(n_975),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1219),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1234),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1085),
.A2(n_996),
.B1(n_1015),
.B2(n_986),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1154),
.A2(n_658),
.B1(n_659),
.B2(n_653),
.Y(n_1422)
);

AND2x6_ASAP7_75t_L g1423 ( 
.A(n_1200),
.B(n_477),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1093),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1073),
.Y(n_1425)
);

XOR2xp5_ASAP7_75t_L g1426 ( 
.A(n_1062),
.B(n_954),
.Y(n_1426)
);

NOR2x1p5_ASAP7_75t_L g1427 ( 
.A(n_1170),
.B(n_503),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1097),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1087),
.A2(n_996),
.B1(n_1015),
.B2(n_986),
.Y(n_1429)
);

AND3x2_ASAP7_75t_L g1430 ( 
.A(n_1226),
.B(n_486),
.C(n_479),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1097),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1264),
.B(n_1214),
.C(n_1182),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1103),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1145),
.B(n_505),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1087),
.B(n_986),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1103),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1090),
.B(n_986),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1169),
.B(n_1174),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1094),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1234),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1090),
.B(n_986),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1169),
.B(n_575),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1094),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1215),
.B(n_917),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1210),
.A2(n_664),
.B1(n_665),
.B2(n_663),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1091),
.B(n_1092),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1271),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1096),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1174),
.B(n_575),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1206),
.B(n_917),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1091),
.A2(n_1092),
.B1(n_1214),
.B2(n_1055),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1097),
.Y(n_1452)
);

INVx5_ASAP7_75t_L g1453 ( 
.A(n_1118),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1157),
.B(n_507),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1096),
.Y(n_1455)
);

BUFx4f_ASAP7_75t_L g1456 ( 
.A(n_1103),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1178),
.B(n_1015),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1178),
.B(n_844),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1054),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1219),
.B(n_1015),
.Y(n_1460)
);

AND2x6_ASAP7_75t_L g1461 ( 
.A(n_1207),
.B(n_479),
.Y(n_1461)
);

AO22x2_ASAP7_75t_L g1462 ( 
.A1(n_1054),
.A2(n_926),
.B1(n_509),
.B2(n_516),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1098),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1204),
.B(n_511),
.C(n_508),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1098),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1055),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1100),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1100),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1117),
.Y(n_1469)
);

NOR2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1170),
.B(n_1225),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1101),
.A2(n_996),
.B1(n_1015),
.B2(n_1005),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1101),
.Y(n_1472)
);

BUFx10_ASAP7_75t_L g1473 ( 
.A(n_1225),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1178),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1104),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1219),
.B(n_1221),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1077),
.B(n_513),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1104),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1167),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1263),
.B(n_603),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1236),
.B(n_1015),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1219),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1047),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1106),
.A2(n_996),
.B1(n_1005),
.B2(n_1027),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1073),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1106),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1219),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1047),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1107),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1118),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1246),
.B(n_515),
.C(n_514),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1118),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1244),
.B(n_942),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1147),
.B(n_525),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1107),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_SL g1496 ( 
.A(n_1219),
.B(n_669),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1221),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1155),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1108),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1221),
.B(n_670),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1221),
.B(n_676),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1108),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1110),
.A2(n_1032),
.B1(n_1033),
.B2(n_1027),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1221),
.B(n_689),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1110),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1113),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1257),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1113),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1118),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1207),
.B(n_942),
.Y(n_1510)
);

INVx5_ASAP7_75t_L g1511 ( 
.A(n_1118),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1149),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1115),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1115),
.Y(n_1514)
);

AND2x2_ASAP7_75t_SL g1515 ( 
.A(n_1183),
.B(n_509),
.Y(n_1515)
);

NAND2xp33_ASAP7_75t_L g1516 ( 
.A(n_1059),
.B(n_940),
.Y(n_1516)
);

CKINVDCx14_ASAP7_75t_R g1517 ( 
.A(n_1151),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1208),
.B(n_942),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1321),
.B(n_1165),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1348),
.B(n_1152),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1343),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1432),
.A2(n_1158),
.B1(n_1160),
.B2(n_1061),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1456),
.B(n_1061),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1277),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1343),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1359),
.B(n_1116),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1456),
.B(n_1221),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1356),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1356),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1359),
.B(n_1116),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1367),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1367),
.Y(n_1532)
);

NAND2xp33_ASAP7_75t_L g1533 ( 
.A(n_1295),
.B(n_1208),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1479),
.B(n_1294),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1378),
.Y(n_1535)
);

NAND2xp33_ASAP7_75t_L g1536 ( 
.A(n_1295),
.B(n_1212),
.Y(n_1536)
);

NAND2xp33_ASAP7_75t_L g1537 ( 
.A(n_1295),
.B(n_1212),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_SL g1538 ( 
.A(n_1416),
.B(n_733),
.Y(n_1538)
);

AO221x1_ASAP7_75t_L g1539 ( 
.A1(n_1316),
.A2(n_517),
.B1(n_532),
.B2(n_516),
.C(n_486),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1479),
.B(n_1120),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1294),
.B(n_1304),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1304),
.B(n_1120),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1378),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1273),
.A2(n_1126),
.B1(n_1129),
.B2(n_1124),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1351),
.B(n_1124),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1438),
.B(n_603),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1396),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1375),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1456),
.B(n_1216),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1362),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1405),
.B(n_1126),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1362),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1405),
.B(n_1436),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1396),
.Y(n_1554)
);

NAND3xp33_ASAP7_75t_L g1555 ( 
.A(n_1328),
.B(n_1132),
.C(n_1129),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1436),
.B(n_1132),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1474),
.B(n_1133),
.Y(n_1557)
);

AND2x6_ASAP7_75t_L g1558 ( 
.A(n_1330),
.B(n_1216),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1376),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1273),
.B(n_1220),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1474),
.B(n_1447),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1446),
.A2(n_1222),
.B(n_1220),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1297),
.A2(n_1133),
.B1(n_1136),
.B2(n_1134),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1297),
.B(n_1222),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1424),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1277),
.B(n_1362),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1451),
.A2(n_1229),
.B1(n_1196),
.B2(n_1134),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1424),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1417),
.B(n_1136),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1439),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1416),
.B(n_733),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1277),
.B(n_1229),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1277),
.B(n_1196),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1354),
.B(n_1138),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1425),
.B(n_1138),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1376),
.B(n_1141),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1439),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1354),
.B(n_1141),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1360),
.B(n_1156),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_SL g1580 ( 
.A(n_1372),
.B(n_1196),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1360),
.B(n_1448),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1455),
.B(n_1156),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1463),
.B(n_1166),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1443),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1288),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1467),
.B(n_1166),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1443),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1465),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1468),
.B(n_1177),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1485),
.Y(n_1590)
);

INVx8_ASAP7_75t_L g1591 ( 
.A(n_1408),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_L g1592 ( 
.A(n_1295),
.B(n_1177),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1472),
.B(n_1180),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1478),
.B(n_1180),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1465),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1284),
.B(n_1184),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1389),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1475),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1372),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1284),
.B(n_1272),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1285),
.A2(n_1185),
.B1(n_1186),
.B2(n_1184),
.Y(n_1601)
);

BUFx5_ASAP7_75t_L g1602 ( 
.A(n_1515),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1285),
.A2(n_1186),
.B1(n_1187),
.B2(n_1185),
.Y(n_1603)
);

INVx4_ASAP7_75t_L g1604 ( 
.A(n_1349),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_L g1605 ( 
.A(n_1295),
.B(n_1187),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1486),
.B(n_1190),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1489),
.B(n_1190),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1372),
.B(n_1112),
.Y(n_1608)
);

NOR2xp67_ASAP7_75t_SL g1609 ( 
.A(n_1395),
.B(n_1183),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1498),
.Y(n_1610)
);

O2A1O1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1319),
.A2(n_1195),
.B(n_1199),
.C(n_1194),
.Y(n_1611)
);

INVxp33_ASAP7_75t_L g1612 ( 
.A(n_1480),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1395),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1285),
.A2(n_1270),
.B1(n_1176),
.B2(n_1179),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1332),
.B(n_1358),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1485),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1475),
.Y(n_1617)
);

O2A1O1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1319),
.A2(n_1195),
.B(n_1199),
.C(n_1194),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1499),
.B(n_1270),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1502),
.B(n_1048),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1278),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1450),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1281),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1384),
.B(n_528),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1279),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1286),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1505),
.B(n_1048),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1290),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1442),
.B(n_603),
.Y(n_1629)
);

AND2x6_ASAP7_75t_L g1630 ( 
.A(n_1330),
.B(n_1049),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1296),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1495),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1495),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1433),
.A2(n_1183),
.B1(n_1191),
.B2(n_1084),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1384),
.B(n_529),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1506),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1410),
.A2(n_1176),
.B1(n_1179),
.B2(n_1168),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1470),
.B(n_517),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1302),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1276),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1506),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1508),
.B(n_1049),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1433),
.B(n_1127),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1515),
.B(n_1127),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1513),
.B(n_1168),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1303),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1514),
.B(n_1181),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1333),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1305),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1275),
.B(n_532),
.Y(n_1650)
);

NAND2xp33_ASAP7_75t_L g1651 ( 
.A(n_1329),
.B(n_1127),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1310),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1410),
.B(n_1181),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1328),
.A2(n_536),
.B(n_537),
.C(n_534),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1449),
.B(n_603),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1517),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1276),
.Y(n_1657)
);

NAND2xp33_ASAP7_75t_L g1658 ( 
.A(n_1329),
.B(n_1127),
.Y(n_1658)
);

NOR2xp67_ASAP7_75t_L g1659 ( 
.A(n_1464),
.B(n_699),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1391),
.B(n_543),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1391),
.B(n_546),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1274),
.A2(n_1183),
.B1(n_1191),
.B2(n_1084),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1434),
.B(n_1058),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1314),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1315),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1434),
.B(n_1454),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1322),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1298),
.A2(n_536),
.B1(n_537),
.B2(n_534),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1307),
.B(n_1127),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1454),
.B(n_1058),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1346),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1353),
.B(n_655),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1333),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_L g1674 ( 
.A(n_1329),
.B(n_1131),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1318),
.A2(n_1080),
.B1(n_1153),
.B2(n_1058),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1334),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1364),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1308),
.B(n_1080),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1307),
.A2(n_1084),
.B1(n_1191),
.B2(n_1153),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1369),
.B(n_1080),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1334),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1337),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1377),
.B(n_655),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1346),
.B(n_550),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1517),
.A2(n_729),
.B1(n_655),
.B2(n_540),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1307),
.A2(n_1191),
.B1(n_1084),
.B2(n_1189),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1337),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1400),
.B(n_1153),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1403),
.B(n_1189),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1353),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1289),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1352),
.B(n_554),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1327),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1352),
.B(n_555),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1407),
.B(n_1189),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1413),
.B(n_1241),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1289),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1402),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1414),
.B(n_1241),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1419),
.B(n_1131),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1292),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1339),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1415),
.B(n_1420),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1349),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1477),
.B(n_898),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1292),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1419),
.B(n_1131),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1293),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1293),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1440),
.B(n_1458),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1299),
.B(n_559),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1301),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1458),
.B(n_1241),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1318),
.B(n_563),
.C(n_562),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1419),
.B(n_1131),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1458),
.B(n_1340),
.Y(n_1716)
);

O2A1O1Ixp5_ASAP7_75t_L g1717 ( 
.A1(n_1323),
.A2(n_1251),
.B(n_1211),
.C(n_1224),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1342),
.B(n_1251),
.Y(n_1718)
);

INVx8_ASAP7_75t_L g1719 ( 
.A(n_1408),
.Y(n_1719)
);

INVx4_ASAP7_75t_L g1720 ( 
.A(n_1349),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1314),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1457),
.A2(n_1109),
.B(n_1064),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1357),
.B(n_1251),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1482),
.B(n_1131),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1365),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1287),
.B(n_564),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1512),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1482),
.B(n_1159),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1366),
.B(n_1209),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1482),
.B(n_1159),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1487),
.B(n_1497),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1408),
.A2(n_1211),
.B1(n_1224),
.B2(n_1209),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1370),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1301),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1373),
.B(n_1380),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_SL g1736 ( 
.A(n_1353),
.B(n_655),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1313),
.Y(n_1737)
);

NOR3xp33_ASAP7_75t_L g1738 ( 
.A(n_1275),
.B(n_567),
.C(n_566),
.Y(n_1738)
);

INVx4_ASAP7_75t_L g1739 ( 
.A(n_1349),
.Y(n_1739)
);

INVxp33_ASAP7_75t_L g1740 ( 
.A(n_1325),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1393),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1444),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1444),
.B(n_1254),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1487),
.B(n_1159),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1317),
.B(n_570),
.Y(n_1745)
);

NOR2xp67_ASAP7_75t_L g1746 ( 
.A(n_1491),
.B(n_706),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1444),
.B(n_1397),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1487),
.B(n_1159),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1338),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1313),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1399),
.B(n_1494),
.Y(n_1751)
);

NOR2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1507),
.B(n_572),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1408),
.A2(n_1423),
.B1(n_1461),
.B2(n_1374),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1399),
.B(n_1262),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1497),
.B(n_1159),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1399),
.B(n_1267),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1494),
.B(n_1267),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1326),
.Y(n_1758)
);

NAND2xp33_ASAP7_75t_L g1759 ( 
.A(n_1329),
.B(n_1163),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1320),
.B(n_729),
.Y(n_1760)
);

INVxp67_ASAP7_75t_L g1761 ( 
.A(n_1338),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1324),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1497),
.B(n_1279),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1532),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1532),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1666),
.B(n_1335),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1526),
.B(n_1335),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1602),
.B(n_1317),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1530),
.B(n_1338),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1630),
.Y(n_1770)
);

INVx4_ASAP7_75t_L g1771 ( 
.A(n_1704),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1573),
.A2(n_1453),
.B(n_1428),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1535),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1535),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1648),
.Y(n_1775)
);

NOR3xp33_ASAP7_75t_SL g1776 ( 
.A(n_1726),
.B(n_1507),
.C(n_1283),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1548),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1521),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1758),
.B(n_1374),
.Y(n_1779)
);

INVx3_ASAP7_75t_L g1780 ( 
.A(n_1630),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1525),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1528),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1704),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1648),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1690),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1597),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1615),
.B(n_1374),
.Y(n_1787)
);

INVx5_ASAP7_75t_L g1788 ( 
.A(n_1558),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1600),
.B(n_1317),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1656),
.Y(n_1790)
);

O2A1O1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1684),
.A2(n_1283),
.B(n_1344),
.C(n_1422),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1602),
.B(n_1385),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1673),
.Y(n_1793)
);

NAND2x1p5_ASAP7_75t_L g1794 ( 
.A(n_1524),
.B(n_1411),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1616),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1742),
.B(n_1427),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1529),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_SL g1798 ( 
.A(n_1602),
.B(n_1385),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1610),
.Y(n_1799)
);

AOI21x1_ASAP7_75t_L g1800 ( 
.A1(n_1609),
.A2(n_1435),
.B(n_1409),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1612),
.B(n_1473),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1692),
.A2(n_1408),
.B1(n_1461),
.B2(n_1423),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1673),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1531),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1616),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1596),
.B(n_1398),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1585),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1581),
.A2(n_1381),
.B1(n_1412),
.B2(n_1394),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1590),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1519),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1630),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1694),
.A2(n_1635),
.B1(n_1660),
.B2(n_1624),
.Y(n_1812)
);

INVxp67_ASAP7_75t_SL g1813 ( 
.A(n_1704),
.Y(n_1813)
);

NAND2xp33_ASAP7_75t_L g1814 ( 
.A(n_1602),
.B(n_1591),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1543),
.Y(n_1815)
);

INVx5_ASAP7_75t_L g1816 ( 
.A(n_1558),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1622),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1676),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1676),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_SL g1820 ( 
.A(n_1538),
.B(n_1469),
.C(n_1426),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1661),
.A2(n_1423),
.B1(n_1461),
.B2(n_1398),
.Y(n_1821)
);

AND2x6_ASAP7_75t_SL g1822 ( 
.A(n_1711),
.B(n_1638),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1681),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1671),
.B(n_1398),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1640),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1574),
.B(n_1462),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1576),
.B(n_1385),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1630),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1578),
.B(n_1462),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1681),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1547),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1547),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1579),
.B(n_1462),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1630),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1602),
.A2(n_1461),
.B1(n_1423),
.B2(n_1341),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1602),
.A2(n_1461),
.B1(n_1423),
.B2(n_1341),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1751),
.B(n_1279),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1540),
.B(n_1282),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1640),
.Y(n_1839)
);

AND3x2_ASAP7_75t_SL g1840 ( 
.A(n_1539),
.B(n_1469),
.C(n_1361),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1554),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1520),
.Y(n_1842)
);

BUFx3_ASAP7_75t_L g1843 ( 
.A(n_1657),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1683),
.B(n_1282),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1657),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1682),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1561),
.B(n_1621),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1602),
.B(n_1386),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1682),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_R g1850 ( 
.A(n_1672),
.B(n_1331),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1613),
.B(n_1576),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1623),
.B(n_1282),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1576),
.B(n_1386),
.Y(n_1853)
);

OAI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1612),
.A2(n_1445),
.B1(n_1401),
.B2(n_1493),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1626),
.B(n_1291),
.Y(n_1855)
);

INVx4_ASAP7_75t_L g1856 ( 
.A(n_1704),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1554),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1628),
.B(n_1291),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1664),
.Y(n_1859)
);

BUFx4f_ASAP7_75t_L g1860 ( 
.A(n_1613),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1738),
.A2(n_1329),
.B1(n_1388),
.B2(n_1341),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1613),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1613),
.B(n_1386),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1664),
.B(n_1291),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1687),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1546),
.B(n_1300),
.Y(n_1866)
);

OAI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1560),
.A2(n_1347),
.B(n_1336),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1687),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1721),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1677),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1698),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1604),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1710),
.B(n_1300),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1629),
.B(n_1473),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1565),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1631),
.B(n_1300),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1565),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1691),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1727),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1639),
.B(n_1341),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1691),
.Y(n_1881)
);

INVx2_ASAP7_75t_SL g1882 ( 
.A(n_1749),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1697),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1568),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1741),
.Y(n_1885)
);

BUFx2_ASAP7_75t_SL g1886 ( 
.A(n_1524),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1524),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1697),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1568),
.Y(n_1889)
);

NOR3xp33_ASAP7_75t_SL g1890 ( 
.A(n_1714),
.B(n_590),
.C(n_576),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1604),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1716),
.B(n_1411),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1646),
.B(n_1341),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1649),
.B(n_1388),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1570),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1685),
.A2(n_617),
.B1(n_646),
.B2(n_591),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1573),
.A2(n_1453),
.B(n_1428),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1570),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1652),
.B(n_1388),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1757),
.B(n_1411),
.Y(n_1900)
);

O2A1O1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1654),
.A2(n_1361),
.B(n_1355),
.C(n_1323),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1577),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1701),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1577),
.Y(n_1904)
);

AND2x4_ASAP7_75t_L g1905 ( 
.A(n_1761),
.B(n_1392),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1545),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1753),
.B(n_1411),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1655),
.B(n_1324),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1550),
.B(n_1431),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1584),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1584),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1740),
.B(n_1473),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1569),
.B(n_1430),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1701),
.Y(n_1914)
);

XNOR2xp5_ASAP7_75t_L g1915 ( 
.A(n_1752),
.B(n_1345),
.Y(n_1915)
);

BUFx4f_ASAP7_75t_L g1916 ( 
.A(n_1591),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1665),
.B(n_1667),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1740),
.B(n_1331),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1552),
.B(n_1431),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1587),
.B(n_1280),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_1625),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1575),
.B(n_729),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1693),
.B(n_1280),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1650),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1587),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1599),
.B(n_1431),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1588),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1702),
.B(n_1725),
.Y(n_1928)
);

INVx4_ASAP7_75t_L g1929 ( 
.A(n_1604),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1588),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1733),
.B(n_1388),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1595),
.Y(n_1932)
);

INVx4_ASAP7_75t_L g1933 ( 
.A(n_1720),
.Y(n_1933)
);

NAND2x1p5_ASAP7_75t_L g1934 ( 
.A(n_1720),
.B(n_1431),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1534),
.B(n_1388),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1595),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1706),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1598),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1703),
.B(n_1510),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1560),
.A2(n_1412),
.B1(n_1459),
.B2(n_1394),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1745),
.B(n_1518),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1598),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1582),
.B(n_1481),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1638),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1564),
.A2(n_1412),
.B1(n_1459),
.B2(n_1394),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1650),
.B(n_1280),
.Y(n_1946)
);

INVx2_ASAP7_75t_SL g1947 ( 
.A(n_1617),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1650),
.B(n_1306),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1747),
.B(n_1306),
.Y(n_1949)
);

A2O1A1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1654),
.A2(n_1312),
.B(n_1309),
.C(n_1350),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1617),
.B(n_1306),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1632),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1706),
.Y(n_1953)
);

BUFx8_ASAP7_75t_L g1954 ( 
.A(n_1760),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1583),
.B(n_1311),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1632),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1708),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1571),
.B(n_1406),
.Y(n_1958)
);

AOI22xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1559),
.A2(n_595),
.B1(n_597),
.B2(n_594),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1633),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1625),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1633),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1746),
.A2(n_1500),
.B1(n_1501),
.B2(n_1496),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1541),
.B(n_1387),
.Y(n_1964)
);

INVx8_ASAP7_75t_L g1965 ( 
.A(n_1591),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1636),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1638),
.Y(n_1967)
);

OAI31xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1668),
.A2(n_1379),
.A3(n_1368),
.B(n_1355),
.Y(n_1968)
);

OR2x6_ASAP7_75t_L g1969 ( 
.A(n_1591),
.B(n_1719),
.Y(n_1969)
);

NOR2x2_ASAP7_75t_L g1970 ( 
.A(n_1636),
.B(n_1382),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1708),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1659),
.A2(n_1496),
.B1(n_1501),
.B2(n_1500),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1641),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1922),
.B(n_1906),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1812),
.B(n_1736),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1941),
.B(n_1586),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1810),
.B(n_1705),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1842),
.B(n_1789),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1766),
.B(n_1589),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1810),
.B(n_1735),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1767),
.B(n_1769),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1879),
.B(n_1555),
.Y(n_1982)
);

NAND2xp33_ASAP7_75t_SL g1983 ( 
.A(n_1776),
.B(n_1564),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1879),
.B(n_1553),
.Y(n_1984)
);

NAND2xp33_ASAP7_75t_SL g1985 ( 
.A(n_1850),
.B(n_1720),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1786),
.B(n_1593),
.Y(n_1986)
);

NAND2xp33_ASAP7_75t_SL g1987 ( 
.A(n_1850),
.B(n_1739),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1786),
.B(n_1594),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1777),
.B(n_1606),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1874),
.B(n_1607),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1799),
.B(n_1542),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1913),
.B(n_1641),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1870),
.B(n_1551),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1870),
.B(n_1556),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1787),
.B(n_1557),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1871),
.B(n_1653),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1847),
.B(n_1680),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1871),
.B(n_1563),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1779),
.B(n_1544),
.Y(n_1999)
);

NAND2xp33_ASAP7_75t_SL g2000 ( 
.A(n_1785),
.B(n_1739),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1954),
.B(n_1601),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1785),
.B(n_1739),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1959),
.B(n_1743),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1954),
.B(n_1603),
.Y(n_2004)
);

AND2x2_ASAP7_75t_SL g2005 ( 
.A(n_1968),
.B(n_1658),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1827),
.B(n_1713),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1954),
.B(n_1663),
.Y(n_2007)
);

NAND2xp33_ASAP7_75t_SL g2008 ( 
.A(n_1872),
.B(n_1644),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1924),
.B(n_1754),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1958),
.B(n_1670),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1869),
.B(n_1756),
.Y(n_2011)
);

NAND2xp33_ASAP7_75t_SL g2012 ( 
.A(n_1805),
.B(n_1523),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1912),
.B(n_1625),
.Y(n_2013)
);

NAND2xp33_ASAP7_75t_SL g2014 ( 
.A(n_1805),
.B(n_1523),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_SL g2015 ( 
.A(n_1885),
.B(n_1522),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1908),
.B(n_1709),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1885),
.B(n_1549),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1801),
.B(n_1549),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1817),
.B(n_1566),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1795),
.B(n_1807),
.Y(n_2020)
);

NAND2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1890),
.B(n_1644),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1854),
.B(n_1566),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1860),
.B(n_1580),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1860),
.B(n_1580),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1860),
.B(n_1567),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1791),
.B(n_1619),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1859),
.B(n_1678),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1809),
.B(n_1645),
.Y(n_2028)
);

NAND2xp33_ASAP7_75t_SL g2029 ( 
.A(n_1872),
.B(n_1643),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1908),
.B(n_1709),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1825),
.B(n_1647),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1827),
.B(n_1643),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1827),
.B(n_1614),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1825),
.B(n_1729),
.Y(n_2034)
);

NAND2xp33_ASAP7_75t_SL g2035 ( 
.A(n_1872),
.B(n_1527),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1839),
.B(n_1637),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1839),
.B(n_1675),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1843),
.B(n_1734),
.Y(n_2038)
);

NAND2xp33_ASAP7_75t_SL g2039 ( 
.A(n_1872),
.B(n_1527),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1843),
.B(n_1734),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1853),
.B(n_1669),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1845),
.B(n_1737),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1845),
.B(n_1737),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1939),
.B(n_1712),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1864),
.B(n_1750),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1864),
.B(n_1750),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1943),
.B(n_1712),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1844),
.B(n_1917),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1844),
.B(n_1762),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1864),
.B(n_1944),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1928),
.B(n_1762),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1944),
.B(n_1620),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1967),
.B(n_1627),
.Y(n_2053)
);

NAND2xp33_ASAP7_75t_SL g2054 ( 
.A(n_1891),
.B(n_1669),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1967),
.B(n_1642),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1790),
.B(n_1608),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1853),
.B(n_1608),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1866),
.B(n_1558),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1853),
.B(n_1688),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1824),
.B(n_729),
.Y(n_2060)
);

NAND2xp33_ASAP7_75t_SL g2061 ( 
.A(n_1891),
.B(n_1572),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1882),
.B(n_1689),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1882),
.B(n_1695),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1918),
.B(n_1696),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1905),
.B(n_1699),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1905),
.B(n_1718),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1866),
.B(n_1558),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1905),
.B(n_1723),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1796),
.B(n_1452),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_SL g2070 ( 
.A(n_1891),
.B(n_1459),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1796),
.B(n_1452),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1796),
.B(n_1452),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1891),
.B(n_1806),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1862),
.B(n_1452),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1862),
.B(n_1490),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1862),
.B(n_1923),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1862),
.B(n_1490),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1923),
.B(n_1490),
.Y(n_2078)
);

NAND2xp33_ASAP7_75t_SL g2079 ( 
.A(n_1835),
.B(n_1466),
.Y(n_2079)
);

NAND2xp33_ASAP7_75t_SL g2080 ( 
.A(n_1836),
.B(n_1466),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1923),
.B(n_1490),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1788),
.B(n_1492),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1788),
.B(n_1816),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1788),
.B(n_1816),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_SL g2085 ( 
.A(n_1788),
.B(n_1492),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1949),
.B(n_1964),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1788),
.B(n_1492),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1816),
.B(n_1492),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1964),
.B(n_1558),
.Y(n_2089)
);

NAND2xp33_ASAP7_75t_SL g2090 ( 
.A(n_1929),
.B(n_1466),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1816),
.B(n_1509),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1816),
.B(n_1509),
.Y(n_2092)
);

NAND2xp33_ASAP7_75t_L g2093 ( 
.A(n_1965),
.B(n_1719),
.Y(n_2093)
);

NAND2xp33_ASAP7_75t_SL g2094 ( 
.A(n_1929),
.B(n_1933),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1964),
.B(n_1662),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1837),
.B(n_1826),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1946),
.B(n_1509),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_1851),
.B(n_1572),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1948),
.B(n_1509),
.Y(n_2099)
);

NAND2xp33_ASAP7_75t_SL g2100 ( 
.A(n_1929),
.B(n_1763),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1802),
.B(n_1763),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1933),
.B(n_1562),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1933),
.B(n_1732),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1829),
.B(n_1719),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1833),
.B(n_1371),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1935),
.B(n_1719),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1821),
.B(n_1722),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1778),
.B(n_1418),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1781),
.B(n_1437),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1782),
.B(n_1483),
.Y(n_2110)
);

NAND2xp33_ASAP7_75t_SL g2111 ( 
.A(n_1783),
.B(n_1404),
.Y(n_2111)
);

NAND2xp33_ASAP7_75t_SL g2112 ( 
.A(n_1783),
.B(n_1731),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1797),
.B(n_1804),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1815),
.B(n_1483),
.Y(n_2114)
);

NAND2xp33_ASAP7_75t_SL g2115 ( 
.A(n_1783),
.B(n_1731),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1851),
.B(n_1483),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1880),
.B(n_1488),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1915),
.B(n_898),
.Y(n_2118)
);

NAND2xp33_ASAP7_75t_SL g2119 ( 
.A(n_1783),
.B(n_1382),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1893),
.B(n_1488),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1894),
.B(n_1488),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1899),
.B(n_1679),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1931),
.B(n_1686),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1887),
.B(n_1634),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1887),
.B(n_1390),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1861),
.B(n_1700),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1838),
.B(n_1379),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1955),
.B(n_1700),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1972),
.B(n_1963),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1973),
.B(n_886),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1896),
.B(n_1707),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1852),
.B(n_1707),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_SL g2133 ( 
.A(n_1855),
.B(n_1715),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_1858),
.B(n_1715),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1876),
.B(n_1724),
.Y(n_2135)
);

NAND2xp33_ASAP7_75t_SL g2136 ( 
.A(n_1770),
.B(n_1383),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1921),
.B(n_1724),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1921),
.B(n_1728),
.Y(n_2138)
);

NAND2xp33_ASAP7_75t_SL g2139 ( 
.A(n_1770),
.B(n_1383),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1921),
.B(n_1728),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1961),
.B(n_1730),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1961),
.B(n_1730),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1920),
.B(n_1409),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1961),
.B(n_1744),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1771),
.B(n_1744),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1764),
.B(n_886),
.Y(n_2146)
);

NAND2xp33_ASAP7_75t_SL g2147 ( 
.A(n_1770),
.B(n_1748),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1920),
.B(n_1951),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1771),
.B(n_1856),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1771),
.B(n_1748),
.Y(n_2150)
);

NAND2xp33_ASAP7_75t_SL g2151 ( 
.A(n_1780),
.B(n_1755),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1951),
.B(n_1435),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1856),
.B(n_1755),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1831),
.B(n_1832),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1856),
.B(n_1504),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1775),
.B(n_1441),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1904),
.B(n_1504),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1904),
.B(n_713),
.Y(n_2158)
);

NAND2xp33_ASAP7_75t_SL g2159 ( 
.A(n_1780),
.B(n_1811),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_1820),
.B(n_1368),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1911),
.B(n_1947),
.Y(n_2161)
);

NAND2xp33_ASAP7_75t_SL g2162 ( 
.A(n_1780),
.B(n_1651),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1969),
.B(n_1441),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1969),
.B(n_1460),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1911),
.B(n_737),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_SL g2166 ( 
.A(n_1947),
.B(n_752),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1952),
.B(n_759),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_1822),
.B(n_598),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1952),
.B(n_1428),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1960),
.B(n_1428),
.Y(n_2170)
);

NAND2xp33_ASAP7_75t_SL g2171 ( 
.A(n_1811),
.B(n_1828),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1960),
.B(n_1428),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1808),
.B(n_1453),
.Y(n_2173)
);

NAND2xp33_ASAP7_75t_SL g2174 ( 
.A(n_1811),
.B(n_1651),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1765),
.B(n_1453),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1765),
.B(n_1453),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1775),
.B(n_1363),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1773),
.B(n_1511),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1773),
.B(n_1774),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1774),
.B(n_1511),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1828),
.B(n_1511),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1828),
.B(n_1511),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1834),
.B(n_1511),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_1834),
.B(n_1611),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1834),
.B(n_1618),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1841),
.B(n_599),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1784),
.B(n_1533),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_1857),
.B(n_602),
.Y(n_2188)
);

NAND2xp33_ASAP7_75t_SL g2189 ( 
.A(n_1907),
.B(n_1658),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1784),
.B(n_1533),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_SL g2191 ( 
.A(n_1875),
.B(n_613),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1877),
.B(n_616),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1884),
.B(n_620),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1889),
.B(n_1895),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1793),
.B(n_1536),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1793),
.B(n_1536),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_SL g2197 ( 
.A(n_1898),
.B(n_1902),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1910),
.B(n_622),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_SL g2199 ( 
.A(n_1925),
.B(n_628),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_SL g2200 ( 
.A(n_1927),
.B(n_630),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1930),
.B(n_1932),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_1936),
.B(n_635),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_1938),
.B(n_642),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_1942),
.B(n_643),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1803),
.B(n_1537),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1974),
.B(n_1956),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2154),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1981),
.B(n_1962),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_2005),
.B(n_1768),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2179),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_1978),
.B(n_1907),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2016),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_1977),
.B(n_1980),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2030),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2148),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1976),
.B(n_1966),
.Y(n_2216)
);

OAI22xp5_ASAP7_75t_SL g2217 ( 
.A1(n_2168),
.A2(n_645),
.B1(n_648),
.B2(n_644),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1979),
.B(n_1971),
.Y(n_2218)
);

AND2x4_ASAP7_75t_SL g2219 ( 
.A(n_1992),
.B(n_1969),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1997),
.B(n_1971),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_SL g2221 ( 
.A(n_2005),
.B(n_1768),
.Y(n_2221)
);

INVx1_ASAP7_75t_SL g2222 ( 
.A(n_2020),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2156),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2009),
.B(n_1914),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1989),
.B(n_1914),
.Y(n_2225)
);

OAI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2129),
.A2(n_1950),
.B(n_1873),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1975),
.B(n_1937),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2130),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1990),
.B(n_1937),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2146),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2052),
.A2(n_1916),
.B1(n_1969),
.B2(n_1886),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_2118),
.Y(n_2232)
);

A2O1A1Ixp33_ASAP7_75t_L g2233 ( 
.A1(n_2189),
.A2(n_1901),
.B(n_1605),
.C(n_1592),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2060),
.B(n_2048),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2003),
.B(n_1991),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2051),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2032),
.B(n_2086),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2113),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_2000),
.Y(n_2239)
);

INVxp67_ASAP7_75t_L g2240 ( 
.A(n_1984),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2098),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2194),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2032),
.B(n_1803),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2096),
.B(n_1953),
.Y(n_2244)
);

BUFx2_ASAP7_75t_L g2245 ( 
.A(n_2032),
.Y(n_2245)
);

INVxp67_ASAP7_75t_L g2246 ( 
.A(n_1982),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1996),
.B(n_1953),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2098),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2002),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2197),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2011),
.B(n_1813),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1985),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2201),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1993),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2160),
.B(n_1950),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1986),
.B(n_1957),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_2041),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1988),
.B(n_1818),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2010),
.B(n_1957),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2028),
.B(n_1818),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2098),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2187),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_2041),
.B(n_1863),
.Y(n_2263)
);

INVx4_ASAP7_75t_L g2264 ( 
.A(n_2041),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2027),
.B(n_1819),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1983),
.B(n_1892),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1994),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2019),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2190),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_1985),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2195),
.Y(n_2271)
);

HB1xp67_ASAP7_75t_L g2272 ( 
.A(n_2050),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1987),
.Y(n_2273)
);

INVx1_ASAP7_75t_SL g2274 ( 
.A(n_2053),
.Y(n_2274)
);

NOR2xp67_ASAP7_75t_L g2275 ( 
.A(n_2007),
.B(n_1892),
.Y(n_2275)
);

NOR2xp67_ASAP7_75t_L g2276 ( 
.A(n_2055),
.B(n_1819),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2196),
.Y(n_2277)
);

INVx1_ASAP7_75t_SL g2278 ( 
.A(n_1987),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2205),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_1983),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2038),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2056),
.B(n_1823),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_2033),
.B(n_1863),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2006),
.B(n_1823),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2064),
.B(n_1830),
.Y(n_2285)
);

BUFx2_ASAP7_75t_L g2286 ( 
.A(n_2006),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2040),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_SL g2288 ( 
.A1(n_2033),
.A2(n_656),
.B1(n_657),
.B2(n_652),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2021),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_2033),
.B(n_1792),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2177),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_2001),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1995),
.B(n_1888),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2006),
.B(n_1888),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2095),
.B(n_1830),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2049),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2015),
.B(n_1873),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2047),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2042),
.Y(n_2299)
);

AOI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_2004),
.A2(n_1592),
.B1(n_1605),
.B2(n_1674),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2065),
.A2(n_2066),
.B1(n_2068),
.B2(n_2131),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2018),
.B(n_1846),
.Y(n_2302)
);

XNOR2xp5_ASAP7_75t_L g2303 ( 
.A(n_2186),
.B(n_1792),
.Y(n_2303)
);

AND3x1_ASAP7_75t_SL g2304 ( 
.A(n_1998),
.B(n_558),
.C(n_538),
.Y(n_2304)
);

AO22x1_ASAP7_75t_L g2305 ( 
.A1(n_2163),
.A2(n_662),
.B1(n_666),
.B2(n_660),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2044),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2089),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2105),
.B(n_1846),
.Y(n_2308)
);

INVx3_ASAP7_75t_L g2309 ( 
.A(n_2164),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2073),
.B(n_1849),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2069),
.B(n_1849),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2043),
.Y(n_2312)
);

AND3x1_ASAP7_75t_SL g2313 ( 
.A(n_2071),
.B(n_558),
.C(n_538),
.Y(n_2313)
);

AND3x1_ASAP7_75t_SL g2314 ( 
.A(n_2072),
.B(n_573),
.C(n_540),
.Y(n_2314)
);

AOI22xp33_ASAP7_75t_L g2315 ( 
.A1(n_2022),
.A2(n_1999),
.B1(n_2057),
.B2(n_2036),
.Y(n_2315)
);

INVx2_ASAP7_75t_SL g2316 ( 
.A(n_2076),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2161),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2108),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_2164),
.Y(n_2319)
);

INVxp67_ASAP7_75t_L g2320 ( 
.A(n_2188),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2031),
.B(n_1878),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2017),
.B(n_1798),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2109),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2143),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2034),
.B(n_1878),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2152),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2191),
.B(n_1865),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2192),
.B(n_1865),
.Y(n_2328)
);

AND3x1_ASAP7_75t_SL g2329 ( 
.A(n_2193),
.B(n_581),
.C(n_541),
.Y(n_2329)
);

A2O1A1Ixp33_ASAP7_75t_L g2330 ( 
.A1(n_2189),
.A2(n_2025),
.B(n_2026),
.C(n_2008),
.Y(n_2330)
);

O2A1O1Ixp33_ASAP7_75t_L g2331 ( 
.A1(n_2037),
.A2(n_544),
.B(n_545),
.C(n_541),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2062),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2063),
.B(n_2198),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2199),
.B(n_1868),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2200),
.B(n_1903),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2202),
.B(n_1868),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2203),
.B(n_1798),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2204),
.B(n_1903),
.Y(n_2338)
);

AO22x1_ASAP7_75t_L g2339 ( 
.A1(n_2163),
.A2(n_677),
.B1(n_679),
.B2(n_674),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2013),
.B(n_1881),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2045),
.Y(n_2341)
);

NOR2xp67_ASAP7_75t_L g2342 ( 
.A(n_2158),
.B(n_1881),
.Y(n_2342)
);

INVx3_ASAP7_75t_L g2343 ( 
.A(n_2164),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2165),
.B(n_2166),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2167),
.B(n_1883),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2008),
.B(n_1867),
.Y(n_2346)
);

AND2x4_ASAP7_75t_L g2347 ( 
.A(n_2163),
.B(n_1848),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2110),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2046),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2097),
.B(n_1883),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_2094),
.Y(n_2351)
);

AND3x1_ASAP7_75t_SL g2352 ( 
.A(n_2012),
.B(n_583),
.C(n_544),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2059),
.B(n_1900),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2014),
.B(n_1900),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2128),
.B(n_682),
.Y(n_2355)
);

INVx4_ASAP7_75t_L g2356 ( 
.A(n_2094),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2124),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2104),
.B(n_2023),
.Y(n_2358)
);

BUFx3_ASAP7_75t_L g2359 ( 
.A(n_2058),
.Y(n_2359)
);

AND3x1_ASAP7_75t_SL g2360 ( 
.A(n_2024),
.B(n_585),
.C(n_545),
.Y(n_2360)
);

BUFx6f_ASAP7_75t_L g2361 ( 
.A(n_2083),
.Y(n_2361)
);

AND2x2_ASAP7_75t_SL g2362 ( 
.A(n_2093),
.B(n_1814),
.Y(n_2362)
);

CKINVDCx8_ASAP7_75t_R g2363 ( 
.A(n_2029),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2099),
.B(n_683),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2127),
.B(n_684),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2035),
.B(n_1916),
.Y(n_2366)
);

CKINVDCx20_ASAP7_75t_R g2367 ( 
.A(n_2149),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2078),
.B(n_2081),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2137),
.Y(n_2369)
);

AND2x4_ASAP7_75t_L g2370 ( 
.A(n_2084),
.B(n_1848),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2039),
.Y(n_2371)
);

BUFx10_ASAP7_75t_L g2372 ( 
.A(n_2054),
.Y(n_2372)
);

AOI22x1_ASAP7_75t_L g2373 ( 
.A1(n_2147),
.A2(n_1794),
.B1(n_1897),
.B2(n_1772),
.Y(n_2373)
);

BUFx8_ASAP7_75t_SL g2374 ( 
.A(n_2067),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2157),
.B(n_685),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2114),
.B(n_549),
.Y(n_2376)
);

OAI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2103),
.A2(n_1916),
.B1(n_1965),
.B2(n_1794),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2126),
.B(n_2107),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_2159),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2116),
.B(n_1909),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2132),
.B(n_686),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_2061),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2133),
.B(n_688),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2101),
.B(n_1909),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_R g2385 ( 
.A(n_2162),
.B(n_1965),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2138),
.B(n_1919),
.Y(n_2386)
);

AND3x1_ASAP7_75t_SL g2387 ( 
.A(n_2147),
.B(n_586),
.C(n_549),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2140),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_2159),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2134),
.B(n_691),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2112),
.A2(n_2115),
.B1(n_2106),
.B2(n_2162),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2074),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2075),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2077),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2141),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2112),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2135),
.B(n_695),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2142),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2125),
.B(n_700),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_2145),
.B(n_1919),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2144),
.B(n_1926),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2150),
.B(n_1926),
.Y(n_2402)
);

OR2x6_ASAP7_75t_L g2403 ( 
.A(n_2173),
.B(n_1965),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2153),
.Y(n_2404)
);

AOI22xp5_ASAP7_75t_L g2405 ( 
.A1(n_2115),
.A2(n_1674),
.B1(n_1759),
.B2(n_1814),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2174),
.A2(n_1759),
.B1(n_1537),
.B2(n_707),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2175),
.Y(n_2407)
);

INVxp67_ASAP7_75t_L g2408 ( 
.A(n_2176),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2122),
.B(n_1800),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2178),
.Y(n_2410)
);

INVx1_ASAP7_75t_SL g2411 ( 
.A(n_2171),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2180),
.Y(n_2412)
);

INVx1_ASAP7_75t_SL g2413 ( 
.A(n_2171),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2123),
.B(n_1934),
.Y(n_2414)
);

INVx3_ASAP7_75t_L g2415 ( 
.A(n_2174),
.Y(n_2415)
);

OAI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2082),
.A2(n_1934),
.B1(n_1945),
.B2(n_1940),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_2151),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2155),
.B(n_702),
.Y(n_2418)
);

OAI22xp5_ASAP7_75t_L g2419 ( 
.A1(n_2085),
.A2(n_1970),
.B1(n_1840),
.B2(n_718),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2184),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2117),
.B(n_710),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2100),
.B(n_1840),
.Y(n_2422)
);

OAI221xp5_ASAP7_75t_L g2423 ( 
.A1(n_2151),
.A2(n_560),
.B1(n_573),
.B2(n_557),
.C(n_552),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2120),
.B(n_719),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2169),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2100),
.B(n_2090),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2121),
.B(n_725),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2185),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2170),
.B(n_552),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2087),
.B(n_730),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2172),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2088),
.B(n_557),
.Y(n_2432)
);

OAI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2102),
.A2(n_1717),
.B(n_1516),
.Y(n_2433)
);

OAI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2111),
.A2(n_1516),
.B(n_1503),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2181),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2182),
.Y(n_2436)
);

NAND2x1p5_ASAP7_75t_L g2437 ( 
.A(n_2091),
.B(n_1970),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2183),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2092),
.B(n_734),
.Y(n_2439)
);

BUFx4f_ASAP7_75t_L g2440 ( 
.A(n_2070),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2111),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2070),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_SL g2443 ( 
.A(n_2090),
.B(n_887),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2136),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2079),
.B(n_741),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2079),
.B(n_742),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2080),
.B(n_745),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2080),
.B(n_2119),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2136),
.B(n_746),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2139),
.B(n_747),
.Y(n_2450)
);

AO21x1_ASAP7_75t_L g2451 ( 
.A1(n_2119),
.A2(n_581),
.B(n_560),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2139),
.Y(n_2452)
);

BUFx4f_ASAP7_75t_L g2453 ( 
.A(n_2005),
.Y(n_2453)
);

BUFx6f_ASAP7_75t_L g2454 ( 
.A(n_2032),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_1974),
.B(n_583),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2154),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_1976),
.B(n_749),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1976),
.B(n_750),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2154),
.Y(n_2459)
);

OAI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2129),
.A2(n_1429),
.B(n_1421),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2154),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_1974),
.B(n_585),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_1974),
.B(n_586),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2164),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_1992),
.Y(n_2465)
);

OAI22xp5_ASAP7_75t_SL g2466 ( 
.A1(n_2168),
.A2(n_753),
.B1(n_754),
.B2(n_751),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2154),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1976),
.B(n_756),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_1974),
.B(n_587),
.Y(n_2469)
);

CKINVDCx16_ASAP7_75t_R g2470 ( 
.A(n_2118),
.Y(n_2470)
);

AOI22xp5_ASAP7_75t_L g2471 ( 
.A1(n_1975),
.A2(n_767),
.B1(n_768),
.B2(n_762),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2154),
.Y(n_2472)
);

INVx2_ASAP7_75t_SL g2473 ( 
.A(n_2020),
.Y(n_2473)
);

OR2x6_ASAP7_75t_L g2474 ( 
.A(n_2403),
.B(n_1238),
.Y(n_2474)
);

NAND2x1p5_ASAP7_75t_L g2475 ( 
.A(n_2426),
.B(n_1238),
.Y(n_2475)
);

INVx3_ASAP7_75t_L g2476 ( 
.A(n_2347),
.Y(n_2476)
);

AO21x1_ASAP7_75t_L g2477 ( 
.A1(n_2378),
.A2(n_592),
.B(n_587),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2241),
.Y(n_2478)
);

BUFx8_ASAP7_75t_L g2479 ( 
.A(n_2270),
.Y(n_2479)
);

AND2x2_ASAP7_75t_SL g2480 ( 
.A(n_2453),
.B(n_592),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2241),
.Y(n_2481)
);

INVx3_ASAP7_75t_L g2482 ( 
.A(n_2347),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2237),
.B(n_593),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2248),
.Y(n_2484)
);

NAND3xp33_ASAP7_75t_SL g2485 ( 
.A(n_2232),
.B(n_601),
.C(n_593),
.Y(n_2485)
);

OAI21x1_ASAP7_75t_L g2486 ( 
.A1(n_2373),
.A2(n_1254),
.B(n_1242),
.Y(n_2486)
);

INVx8_ASAP7_75t_L g2487 ( 
.A(n_2263),
.Y(n_2487)
);

OAI21xp5_ASAP7_75t_L g2488 ( 
.A1(n_2330),
.A2(n_606),
.B(n_601),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2248),
.Y(n_2489)
);

OAI21x1_ASAP7_75t_L g2490 ( 
.A1(n_2433),
.A2(n_1255),
.B(n_1242),
.Y(n_2490)
);

OAI21x1_ASAP7_75t_L g2491 ( 
.A1(n_2226),
.A2(n_1262),
.B(n_1255),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2234),
.B(n_606),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2261),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2347),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2261),
.Y(n_2495)
);

OAI21xp5_ASAP7_75t_L g2496 ( 
.A1(n_2330),
.A2(n_611),
.B(n_608),
.Y(n_2496)
);

NOR2x1_ASAP7_75t_L g2497 ( 
.A(n_2356),
.B(n_608),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2211),
.B(n_611),
.Y(n_2498)
);

AO21x2_ASAP7_75t_L g2499 ( 
.A1(n_2354),
.A2(n_845),
.B(n_844),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2420),
.Y(n_2500)
);

BUFx2_ASAP7_75t_L g2501 ( 
.A(n_2309),
.Y(n_2501)
);

AO21x1_ASAP7_75t_SL g2502 ( 
.A1(n_2405),
.A2(n_621),
.B(n_615),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2232),
.Y(n_2503)
);

BUFx3_ASAP7_75t_L g2504 ( 
.A(n_2465),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_2465),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2470),
.Y(n_2506)
);

HB1xp67_ASAP7_75t_L g2507 ( 
.A(n_2207),
.Y(n_2507)
);

AO21x2_ASAP7_75t_L g2508 ( 
.A1(n_2354),
.A2(n_2346),
.B(n_2255),
.Y(n_2508)
);

OAI21x1_ASAP7_75t_L g2509 ( 
.A1(n_2426),
.A2(n_2415),
.B(n_2441),
.Y(n_2509)
);

INVx2_ASAP7_75t_SL g2510 ( 
.A(n_2207),
.Y(n_2510)
);

OAI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2457),
.A2(n_621),
.B(n_615),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2307),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2420),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_2309),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2274),
.B(n_627),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2309),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2428),
.Y(n_2517)
);

INVx5_ASAP7_75t_L g2518 ( 
.A(n_2356),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2428),
.Y(n_2519)
);

INVx3_ASAP7_75t_L g2520 ( 
.A(n_2319),
.Y(n_2520)
);

AO21x2_ASAP7_75t_L g2521 ( 
.A1(n_2346),
.A2(n_848),
.B(n_845),
.Y(n_2521)
);

BUFx12f_ASAP7_75t_L g2522 ( 
.A(n_2289),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2357),
.Y(n_2523)
);

OAI21x1_ASAP7_75t_L g2524 ( 
.A1(n_2415),
.A2(n_1460),
.B(n_1053),
.Y(n_2524)
);

BUFx12f_ASAP7_75t_L g2525 ( 
.A(n_2289),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2319),
.Y(n_2526)
);

OAI21x1_ASAP7_75t_L g2527 ( 
.A1(n_2415),
.A2(n_1053),
.B(n_1051),
.Y(n_2527)
);

OAI21x1_ASAP7_75t_L g2528 ( 
.A1(n_2441),
.A2(n_1066),
.B(n_1051),
.Y(n_2528)
);

AO21x2_ASAP7_75t_L g2529 ( 
.A1(n_2255),
.A2(n_851),
.B(n_848),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2319),
.B(n_318),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2307),
.Y(n_2531)
);

BUFx10_ASAP7_75t_L g2532 ( 
.A(n_2337),
.Y(n_2532)
);

OAI21x1_ASAP7_75t_SL g2533 ( 
.A1(n_2451),
.A2(n_2358),
.B(n_2315),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2343),
.Y(n_2534)
);

NAND2x1p5_ASAP7_75t_L g2535 ( 
.A(n_2362),
.B(n_1064),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2237),
.B(n_627),
.Y(n_2536)
);

INVx4_ASAP7_75t_L g2537 ( 
.A(n_2440),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_L g2538 ( 
.A(n_2362),
.B(n_1064),
.Y(n_2538)
);

BUFx3_ASAP7_75t_L g2539 ( 
.A(n_2206),
.Y(n_2539)
);

CKINVDCx14_ASAP7_75t_R g2540 ( 
.A(n_2455),
.Y(n_2540)
);

AO21x2_ASAP7_75t_L g2541 ( 
.A1(n_2422),
.A2(n_2448),
.B(n_2297),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2343),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2343),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2453),
.B(n_2295),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2464),
.Y(n_2545)
);

BUFx2_ASAP7_75t_L g2546 ( 
.A(n_2464),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2464),
.Y(n_2547)
);

INVx4_ASAP7_75t_L g2548 ( 
.A(n_2440),
.Y(n_2548)
);

AO21x1_ASAP7_75t_L g2549 ( 
.A1(n_2378),
.A2(n_633),
.B(n_631),
.Y(n_2549)
);

OAI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2458),
.A2(n_633),
.B(n_631),
.Y(n_2550)
);

OAI21x1_ASAP7_75t_L g2551 ( 
.A1(n_2379),
.A2(n_1069),
.B(n_1066),
.Y(n_2551)
);

AND2x4_ASAP7_75t_L g2552 ( 
.A(n_2290),
.B(n_321),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_2379),
.Y(n_2553)
);

AO21x2_ASAP7_75t_L g2554 ( 
.A1(n_2422),
.A2(n_854),
.B(n_851),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2459),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2459),
.Y(n_2556)
);

INVx2_ASAP7_75t_SL g2557 ( 
.A(n_2472),
.Y(n_2557)
);

OA21x2_ASAP7_75t_L g2558 ( 
.A1(n_2448),
.A2(n_858),
.B(n_854),
.Y(n_2558)
);

OAI21x1_ASAP7_75t_L g2559 ( 
.A1(n_2379),
.A2(n_1076),
.B(n_1069),
.Y(n_2559)
);

OAI21x1_ASAP7_75t_L g2560 ( 
.A1(n_2266),
.A2(n_1083),
.B(n_1076),
.Y(n_2560)
);

BUFx8_ASAP7_75t_L g2561 ( 
.A(n_2462),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2357),
.Y(n_2562)
);

BUFx3_ASAP7_75t_L g2563 ( 
.A(n_2472),
.Y(n_2563)
);

OAI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_2468),
.A2(n_641),
.B(n_640),
.Y(n_2564)
);

HB1xp67_ASAP7_75t_L g2565 ( 
.A(n_2456),
.Y(n_2565)
);

AOI22xp33_ASAP7_75t_L g2566 ( 
.A1(n_2453),
.A2(n_641),
.B1(n_661),
.B2(n_640),
.Y(n_2566)
);

OAI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2365),
.A2(n_673),
.B(n_661),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2409),
.Y(n_2568)
);

BUFx2_ASAP7_75t_L g2569 ( 
.A(n_2359),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2409),
.Y(n_2570)
);

AO21x2_ASAP7_75t_L g2571 ( 
.A1(n_2297),
.A2(n_859),
.B(n_858),
.Y(n_2571)
);

OAI21x1_ASAP7_75t_SL g2572 ( 
.A1(n_2301),
.A2(n_870),
.B(n_861),
.Y(n_2572)
);

BUFx3_ASAP7_75t_L g2573 ( 
.A(n_2374),
.Y(n_2573)
);

BUFx4_ASAP7_75t_SL g2574 ( 
.A(n_2292),
.Y(n_2574)
);

INVxp67_ASAP7_75t_SL g2575 ( 
.A(n_2298),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2395),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2369),
.Y(n_2577)
);

INVx2_ASAP7_75t_SL g2578 ( 
.A(n_2257),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2369),
.Y(n_2579)
);

INVx2_ASAP7_75t_SL g2580 ( 
.A(n_2257),
.Y(n_2580)
);

OAI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2445),
.A2(n_681),
.B(n_673),
.Y(n_2581)
);

BUFx2_ASAP7_75t_L g2582 ( 
.A(n_2359),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2295),
.B(n_681),
.Y(n_2583)
);

HB1xp67_ASAP7_75t_L g2584 ( 
.A(n_2461),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2257),
.Y(n_2585)
);

CKINVDCx11_ASAP7_75t_R g2586 ( 
.A(n_2222),
.Y(n_2586)
);

OAI21x1_ASAP7_75t_L g2587 ( 
.A1(n_2266),
.A2(n_1088),
.B(n_1083),
.Y(n_2587)
);

AO21x2_ASAP7_75t_L g2588 ( 
.A1(n_2233),
.A2(n_860),
.B(n_859),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2388),
.Y(n_2589)
);

HB1xp67_ASAP7_75t_L g2590 ( 
.A(n_2467),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2290),
.Y(n_2591)
);

AND2x4_ASAP7_75t_L g2592 ( 
.A(n_2290),
.B(n_322),
.Y(n_2592)
);

AO21x2_ASAP7_75t_L g2593 ( 
.A1(n_2233),
.A2(n_862),
.B(n_860),
.Y(n_2593)
);

AO21x2_ASAP7_75t_L g2594 ( 
.A1(n_2209),
.A2(n_863),
.B(n_862),
.Y(n_2594)
);

BUFx3_ASAP7_75t_L g2595 ( 
.A(n_2374),
.Y(n_2595)
);

OR2x6_ASAP7_75t_L g2596 ( 
.A(n_2403),
.B(n_861),
.Y(n_2596)
);

AO21x2_ASAP7_75t_L g2597 ( 
.A1(n_2209),
.A2(n_2221),
.B(n_2391),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2417),
.Y(n_2598)
);

NOR2x1_ASAP7_75t_L g2599 ( 
.A(n_2356),
.B(n_690),
.Y(n_2599)
);

INVx2_ASAP7_75t_SL g2600 ( 
.A(n_2257),
.Y(n_2600)
);

INVx4_ASAP7_75t_L g2601 ( 
.A(n_2440),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2454),
.Y(n_2602)
);

CKINVDCx20_ASAP7_75t_R g2603 ( 
.A(n_2367),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2243),
.B(n_690),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2388),
.Y(n_2605)
);

INVx3_ASAP7_75t_SL g2606 ( 
.A(n_2239),
.Y(n_2606)
);

AOI22x1_ASAP7_75t_L g2607 ( 
.A1(n_2280),
.A2(n_693),
.B1(n_697),
.B2(n_692),
.Y(n_2607)
);

INVx1_ASAP7_75t_SL g2608 ( 
.A(n_2213),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2211),
.B(n_692),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2398),
.Y(n_2610)
);

OAI21x1_ASAP7_75t_L g2611 ( 
.A1(n_2444),
.A2(n_1089),
.B(n_1088),
.Y(n_2611)
);

OAI21xp5_ASAP7_75t_L g2612 ( 
.A1(n_2446),
.A2(n_697),
.B(n_693),
.Y(n_2612)
);

OAI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2447),
.A2(n_705),
.B(n_701),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2243),
.B(n_701),
.Y(n_2614)
);

BUFx4f_ASAP7_75t_L g2615 ( 
.A(n_2437),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2398),
.Y(n_2616)
);

OAI21x1_ASAP7_75t_L g2617 ( 
.A1(n_2452),
.A2(n_1099),
.B(n_1089),
.Y(n_2617)
);

BUFx2_ASAP7_75t_L g2618 ( 
.A(n_2389),
.Y(n_2618)
);

OAI21x1_ASAP7_75t_L g2619 ( 
.A1(n_2416),
.A2(n_1111),
.B(n_1099),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2262),
.Y(n_2620)
);

BUFx12f_ASAP7_75t_L g2621 ( 
.A(n_2463),
.Y(n_2621)
);

BUFx3_ASAP7_75t_L g2622 ( 
.A(n_2251),
.Y(n_2622)
);

BUFx3_ASAP7_75t_L g2623 ( 
.A(n_2473),
.Y(n_2623)
);

AOI21x1_ASAP7_75t_L g2624 ( 
.A1(n_2443),
.A2(n_864),
.B(n_863),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2293),
.Y(n_2625)
);

NAND2x1p5_ASAP7_75t_L g2626 ( 
.A(n_2366),
.B(n_1109),
.Y(n_2626)
);

OAI21x1_ASAP7_75t_L g2627 ( 
.A1(n_2434),
.A2(n_1114),
.B(n_1111),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2298),
.Y(n_2628)
);

AO21x2_ASAP7_75t_L g2629 ( 
.A1(n_2221),
.A2(n_865),
.B(n_864),
.Y(n_2629)
);

OAI21x1_ASAP7_75t_L g2630 ( 
.A1(n_2442),
.A2(n_1121),
.B(n_1114),
.Y(n_2630)
);

OAI21x1_ASAP7_75t_L g2631 ( 
.A1(n_2366),
.A2(n_1122),
.B(n_1121),
.Y(n_2631)
);

AO21x2_ASAP7_75t_L g2632 ( 
.A1(n_2443),
.A2(n_866),
.B(n_865),
.Y(n_2632)
);

OAI21x1_ASAP7_75t_L g2633 ( 
.A1(n_2353),
.A2(n_2377),
.B(n_2269),
.Y(n_2633)
);

BUFx2_ASAP7_75t_R g2634 ( 
.A(n_2292),
.Y(n_2634)
);

AND2x4_ASAP7_75t_L g2635 ( 
.A(n_2264),
.B(n_324),
.Y(n_2635)
);

OAI21x1_ASAP7_75t_L g2636 ( 
.A1(n_2262),
.A2(n_2269),
.B(n_2310),
.Y(n_2636)
);

BUFx2_ASAP7_75t_R g2637 ( 
.A(n_2252),
.Y(n_2637)
);

OA21x2_ASAP7_75t_L g2638 ( 
.A1(n_2384),
.A2(n_867),
.B(n_866),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2306),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2306),
.Y(n_2640)
);

INVx4_ASAP7_75t_L g2641 ( 
.A(n_2351),
.Y(n_2641)
);

OR2x6_ASAP7_75t_SL g2642 ( 
.A(n_2396),
.B(n_705),
.Y(n_2642)
);

AO21x2_ASAP7_75t_L g2643 ( 
.A1(n_2384),
.A2(n_872),
.B(n_867),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2215),
.B(n_711),
.Y(n_2644)
);

INVx4_ASAP7_75t_L g2645 ( 
.A(n_2351),
.Y(n_2645)
);

INVxp67_ASAP7_75t_SL g2646 ( 
.A(n_2296),
.Y(n_2646)
);

INVx3_ASAP7_75t_L g2647 ( 
.A(n_2264),
.Y(n_2647)
);

AOI22x1_ASAP7_75t_L g2648 ( 
.A1(n_2280),
.A2(n_715),
.B1(n_723),
.B2(n_711),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2246),
.B(n_715),
.Y(n_2649)
);

INVx8_ASAP7_75t_L g2650 ( 
.A(n_2263),
.Y(n_2650)
);

INVx4_ASAP7_75t_L g2651 ( 
.A(n_2372),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2245),
.B(n_723),
.Y(n_2652)
);

OAI21x1_ASAP7_75t_SL g2653 ( 
.A1(n_2227),
.A2(n_875),
.B(n_870),
.Y(n_2653)
);

CKINVDCx11_ASAP7_75t_R g2654 ( 
.A(n_2363),
.Y(n_2654)
);

AOI22x1_ASAP7_75t_L g2655 ( 
.A1(n_2303),
.A2(n_727),
.B1(n_739),
.B2(n_726),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2404),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2323),
.Y(n_2657)
);

NAND2x1p5_ASAP7_75t_L g2658 ( 
.A(n_2278),
.B(n_1109),
.Y(n_2658)
);

BUFx2_ASAP7_75t_L g2659 ( 
.A(n_2400),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2323),
.Y(n_2660)
);

BUFx2_ASAP7_75t_R g2661 ( 
.A(n_2252),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2324),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2215),
.B(n_726),
.Y(n_2663)
);

INVx8_ASAP7_75t_L g2664 ( 
.A(n_2263),
.Y(n_2664)
);

OAI21x1_ASAP7_75t_L g2665 ( 
.A1(n_2436),
.A2(n_1139),
.B(n_1122),
.Y(n_2665)
);

OAI21x1_ASAP7_75t_L g2666 ( 
.A1(n_2436),
.A2(n_2438),
.B(n_2340),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2473),
.Y(n_2667)
);

OAI21x1_ASAP7_75t_SL g2668 ( 
.A1(n_2282),
.A2(n_881),
.B(n_875),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2236),
.Y(n_2669)
);

BUFx3_ASAP7_75t_L g2670 ( 
.A(n_2454),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2236),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2291),
.B(n_727),
.Y(n_2672)
);

AND2x4_ASAP7_75t_L g2673 ( 
.A(n_2264),
.B(n_325),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2259),
.Y(n_2674)
);

BUFx2_ASAP7_75t_SL g2675 ( 
.A(n_2363),
.Y(n_2675)
);

BUFx6f_ASAP7_75t_L g2676 ( 
.A(n_2454),
.Y(n_2676)
);

INVx4_ASAP7_75t_L g2677 ( 
.A(n_2372),
.Y(n_2677)
);

OA21x2_ASAP7_75t_L g2678 ( 
.A1(n_2386),
.A2(n_876),
.B(n_872),
.Y(n_2678)
);

OAI21xp5_ASAP7_75t_L g2679 ( 
.A1(n_2355),
.A2(n_755),
.B(n_739),
.Y(n_2679)
);

NAND2x1p5_ASAP7_75t_L g2680 ( 
.A(n_2400),
.B(n_1119),
.Y(n_2680)
);

AO21x2_ASAP7_75t_L g2681 ( 
.A1(n_2275),
.A2(n_877),
.B(n_876),
.Y(n_2681)
);

HB1xp67_ASAP7_75t_L g2682 ( 
.A(n_2272),
.Y(n_2682)
);

AO21x2_ASAP7_75t_L g2683 ( 
.A1(n_2385),
.A2(n_878),
.B(n_877),
.Y(n_2683)
);

INVx3_ASAP7_75t_SL g2684 ( 
.A(n_2239),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2216),
.A2(n_1476),
.B(n_1471),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2302),
.Y(n_2686)
);

INVx4_ASAP7_75t_L g2687 ( 
.A(n_2372),
.Y(n_2687)
);

HB1xp67_ASAP7_75t_L g2688 ( 
.A(n_2258),
.Y(n_2688)
);

OAI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2320),
.A2(n_758),
.B(n_755),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2210),
.Y(n_2690)
);

BUFx12f_ASAP7_75t_L g2691 ( 
.A(n_2469),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2454),
.Y(n_2692)
);

OAI21x1_ASAP7_75t_L g2693 ( 
.A1(n_2438),
.A2(n_1140),
.B(n_1139),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2324),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2291),
.B(n_758),
.Y(n_2695)
);

BUFx2_ASAP7_75t_R g2696 ( 
.A(n_2273),
.Y(n_2696)
);

INVx5_ASAP7_75t_L g2697 ( 
.A(n_2403),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2210),
.Y(n_2698)
);

OAI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2381),
.A2(n_764),
.B(n_760),
.Y(n_2699)
);

OAI21x1_ASAP7_75t_L g2700 ( 
.A1(n_2414),
.A2(n_1148),
.B(n_1140),
.Y(n_2700)
);

BUFx8_ASAP7_75t_L g2701 ( 
.A(n_2344),
.Y(n_2701)
);

AOI22x1_ASAP7_75t_L g2702 ( 
.A1(n_2396),
.A2(n_764),
.B1(n_760),
.B2(n_887),
.Y(n_2702)
);

HB1xp67_ASAP7_75t_L g2703 ( 
.A(n_2254),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2224),
.B(n_881),
.Y(n_2704)
);

AOI22xp33_ASAP7_75t_L g2705 ( 
.A1(n_2288),
.A2(n_889),
.B1(n_891),
.B2(n_888),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2229),
.Y(n_2706)
);

OAI21x1_ASAP7_75t_L g2707 ( 
.A1(n_2414),
.A2(n_1150),
.B(n_1148),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2326),
.Y(n_2708)
);

AO21x2_ASAP7_75t_L g2709 ( 
.A1(n_2385),
.A2(n_879),
.B(n_878),
.Y(n_2709)
);

AO21x2_ASAP7_75t_L g2710 ( 
.A1(n_2300),
.A2(n_880),
.B(n_879),
.Y(n_2710)
);

BUFx3_ASAP7_75t_L g2711 ( 
.A(n_2361),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_2235),
.B(n_888),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2361),
.Y(n_2713)
);

AO21x2_ASAP7_75t_L g2714 ( 
.A1(n_2449),
.A2(n_883),
.B(n_880),
.Y(n_2714)
);

BUFx4f_ASAP7_75t_SL g2715 ( 
.A(n_2367),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2326),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_L g2717 ( 
.A(n_2240),
.B(n_330),
.Y(n_2717)
);

CKINVDCx20_ASAP7_75t_R g2718 ( 
.A(n_2286),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2247),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2223),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_L g2721 ( 
.A1(n_2283),
.A2(n_891),
.B1(n_892),
.B2(n_889),
.Y(n_2721)
);

AO21x2_ASAP7_75t_L g2722 ( 
.A1(n_2450),
.A2(n_884),
.B(n_883),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2223),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2283),
.B(n_331),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_2249),
.Y(n_2725)
);

INVx4_ASAP7_75t_L g2726 ( 
.A(n_2273),
.Y(n_2726)
);

BUFx3_ASAP7_75t_L g2727 ( 
.A(n_2361),
.Y(n_2727)
);

OA21x2_ASAP7_75t_L g2728 ( 
.A1(n_2386),
.A2(n_884),
.B(n_892),
.Y(n_2728)
);

OAI21x1_ASAP7_75t_L g2729 ( 
.A1(n_2231),
.A2(n_1162),
.B(n_1150),
.Y(n_2729)
);

NAND2x1p5_ASAP7_75t_L g2730 ( 
.A(n_2400),
.B(n_2411),
.Y(n_2730)
);

OAI21x1_ASAP7_75t_L g2731 ( 
.A1(n_2401),
.A2(n_1162),
.B(n_1484),
.Y(n_2731)
);

BUFx12f_ASAP7_75t_L g2732 ( 
.A(n_2249),
.Y(n_2732)
);

OR2x6_ASAP7_75t_L g2733 ( 
.A(n_2403),
.B(n_893),
.Y(n_2733)
);

BUFx3_ASAP7_75t_L g2734 ( 
.A(n_2361),
.Y(n_2734)
);

BUFx8_ASAP7_75t_L g2735 ( 
.A(n_2522),
.Y(n_2735)
);

INVx3_ASAP7_75t_SL g2736 ( 
.A(n_2503),
.Y(n_2736)
);

AOI22xp33_ASAP7_75t_L g2737 ( 
.A1(n_2480),
.A2(n_2283),
.B1(n_2337),
.B2(n_2423),
.Y(n_2737)
);

AOI22xp33_ASAP7_75t_L g2738 ( 
.A1(n_2480),
.A2(n_2430),
.B1(n_2268),
.B2(n_2217),
.Y(n_2738)
);

CKINVDCx20_ASAP7_75t_R g2739 ( 
.A(n_2654),
.Y(n_2739)
);

BUFx3_ASAP7_75t_L g2740 ( 
.A(n_2573),
.Y(n_2740)
);

INVx4_ASAP7_75t_L g2741 ( 
.A(n_2651),
.Y(n_2741)
);

AOI22xp33_ASAP7_75t_SL g2742 ( 
.A1(n_2480),
.A2(n_2655),
.B1(n_2715),
.B2(n_2689),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2656),
.Y(n_2743)
);

OAI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2642),
.A2(n_2382),
.B1(n_2371),
.B2(n_2230),
.Y(n_2744)
);

INVx4_ASAP7_75t_L g2745 ( 
.A(n_2651),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2544),
.B(n_2267),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2656),
.Y(n_2747)
);

AOI22xp33_ASAP7_75t_L g2748 ( 
.A1(n_2655),
.A2(n_2430),
.B1(n_2466),
.B2(n_2322),
.Y(n_2748)
);

AOI22xp33_ASAP7_75t_L g2749 ( 
.A1(n_2621),
.A2(n_2322),
.B1(n_2419),
.B2(n_2318),
.Y(n_2749)
);

BUFx2_ASAP7_75t_R g2750 ( 
.A(n_2675),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2576),
.Y(n_2751)
);

AOI22xp33_ASAP7_75t_L g2752 ( 
.A1(n_2621),
.A2(n_2418),
.B1(n_2228),
.B2(n_2390),
.Y(n_2752)
);

AOI22xp33_ASAP7_75t_L g2753 ( 
.A1(n_2691),
.A2(n_2383),
.B1(n_2397),
.B2(n_2332),
.Y(n_2753)
);

HB1xp67_ASAP7_75t_L g2754 ( 
.A(n_2508),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2556),
.Y(n_2755)
);

AOI22xp33_ASAP7_75t_L g2756 ( 
.A1(n_2691),
.A2(n_2376),
.B1(n_2333),
.B2(n_2345),
.Y(n_2756)
);

AOI22xp5_ASAP7_75t_L g2757 ( 
.A1(n_2581),
.A2(n_2613),
.B1(n_2612),
.B2(n_2550),
.Y(n_2757)
);

INVx1_ASAP7_75t_SL g2758 ( 
.A(n_2586),
.Y(n_2758)
);

INVx6_ASAP7_75t_L g2759 ( 
.A(n_2561),
.Y(n_2759)
);

INVx4_ASAP7_75t_L g2760 ( 
.A(n_2651),
.Y(n_2760)
);

AOI22xp33_ASAP7_75t_L g2761 ( 
.A1(n_2511),
.A2(n_2370),
.B1(n_2375),
.B2(n_2429),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2576),
.Y(n_2762)
);

INVx3_ASAP7_75t_L g2763 ( 
.A(n_2556),
.Y(n_2763)
);

CKINVDCx16_ASAP7_75t_R g2764 ( 
.A(n_2603),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2563),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2657),
.Y(n_2766)
);

AOI22xp33_ASAP7_75t_L g2767 ( 
.A1(n_2564),
.A2(n_2699),
.B1(n_2679),
.B2(n_2567),
.Y(n_2767)
);

AOI22xp33_ASAP7_75t_L g2768 ( 
.A1(n_2724),
.A2(n_2370),
.B1(n_2316),
.B2(n_2328),
.Y(n_2768)
);

OAI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2642),
.A2(n_2382),
.B1(n_2371),
.B2(n_2406),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2724),
.A2(n_2370),
.B1(n_2316),
.B2(n_2334),
.Y(n_2770)
);

AOI22xp33_ASAP7_75t_SL g2771 ( 
.A1(n_2561),
.A2(n_2413),
.B1(n_2304),
.B2(n_2238),
.Y(n_2771)
);

INVx6_ASAP7_75t_L g2772 ( 
.A(n_2561),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2657),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2701),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2660),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2574),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2660),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2575),
.B(n_2271),
.Y(n_2778)
);

CKINVDCx5p33_ASAP7_75t_R g2779 ( 
.A(n_2503),
.Y(n_2779)
);

CKINVDCx20_ASAP7_75t_R g2780 ( 
.A(n_2718),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2540),
.A2(n_2329),
.B1(n_2360),
.B2(n_2352),
.Y(n_2781)
);

OAI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2566),
.A2(n_2437),
.B1(n_2471),
.B2(n_2250),
.Y(n_2782)
);

INVx2_ASAP7_75t_SL g2783 ( 
.A(n_2539),
.Y(n_2783)
);

HB1xp67_ASAP7_75t_L g2784 ( 
.A(n_2508),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2634),
.A2(n_2253),
.B1(n_2242),
.B2(n_2277),
.Y(n_2785)
);

BUFx10_ASAP7_75t_L g2786 ( 
.A(n_2515),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2577),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_SL g2788 ( 
.A1(n_2561),
.A2(n_2219),
.B1(n_2317),
.B2(n_2432),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2577),
.Y(n_2789)
);

OAI22xp33_ASAP7_75t_L g2790 ( 
.A1(n_2498),
.A2(n_2399),
.B1(n_2364),
.B2(n_2276),
.Y(n_2790)
);

CKINVDCx5p33_ASAP7_75t_R g2791 ( 
.A(n_2522),
.Y(n_2791)
);

CKINVDCx11_ASAP7_75t_R g2792 ( 
.A(n_2525),
.Y(n_2792)
);

AOI22xp5_ASAP7_75t_L g2793 ( 
.A1(n_2485),
.A2(n_2339),
.B1(n_2305),
.B2(n_2387),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2563),
.Y(n_2794)
);

OAI22xp33_ASAP7_75t_L g2795 ( 
.A1(n_2609),
.A2(n_2279),
.B1(n_2349),
.B2(n_2341),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2579),
.Y(n_2796)
);

BUFx3_ASAP7_75t_L g2797 ( 
.A(n_2573),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2579),
.Y(n_2798)
);

CKINVDCx20_ASAP7_75t_R g2799 ( 
.A(n_2701),
.Y(n_2799)
);

AOI22xp33_ASAP7_75t_L g2800 ( 
.A1(n_2724),
.A2(n_2336),
.B1(n_2327),
.B2(n_2219),
.Y(n_2800)
);

BUFx8_ASAP7_75t_L g2801 ( 
.A(n_2525),
.Y(n_2801)
);

BUFx3_ASAP7_75t_L g2802 ( 
.A(n_2595),
.Y(n_2802)
);

BUFx6f_ASAP7_75t_L g2803 ( 
.A(n_2713),
.Y(n_2803)
);

INVx3_ASAP7_75t_L g2804 ( 
.A(n_2713),
.Y(n_2804)
);

OAI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2539),
.A2(n_2608),
.B1(n_2496),
.B2(n_2488),
.Y(n_2805)
);

AOI22xp33_ASAP7_75t_SL g2806 ( 
.A1(n_2607),
.A2(n_2402),
.B1(n_2401),
.B2(n_2208),
.Y(n_2806)
);

OAI22xp33_ASAP7_75t_L g2807 ( 
.A1(n_2506),
.A2(n_2439),
.B1(n_2424),
.B2(n_2427),
.Y(n_2807)
);

OAI22x1_ASAP7_75t_SL g2808 ( 
.A1(n_2506),
.A2(n_895),
.B1(n_896),
.B2(n_893),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_SL g2809 ( 
.A1(n_2607),
.A2(n_2402),
.B1(n_2208),
.B2(n_2296),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2615),
.A2(n_2408),
.B1(n_2214),
.B2(n_2212),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2713),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2610),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2713),
.Y(n_2813)
);

INVx1_ASAP7_75t_SL g2814 ( 
.A(n_2606),
.Y(n_2814)
);

BUFx12f_ASAP7_75t_L g2815 ( 
.A(n_2732),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2610),
.Y(n_2816)
);

INVx2_ASAP7_75t_R g2817 ( 
.A(n_2518),
.Y(n_2817)
);

CKINVDCx20_ASAP7_75t_R g2818 ( 
.A(n_2701),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2555),
.Y(n_2819)
);

INVx4_ASAP7_75t_L g2820 ( 
.A(n_2677),
.Y(n_2820)
);

CKINVDCx11_ASAP7_75t_R g2821 ( 
.A(n_2606),
.Y(n_2821)
);

INVx6_ASAP7_75t_L g2822 ( 
.A(n_2479),
.Y(n_2822)
);

AOI22xp5_ASAP7_75t_L g2823 ( 
.A1(n_2675),
.A2(n_2314),
.B1(n_2313),
.B2(n_2342),
.Y(n_2823)
);

OAI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2615),
.A2(n_2214),
.B1(n_2212),
.B2(n_2225),
.Y(n_2824)
);

BUFx3_ASAP7_75t_L g2825 ( 
.A(n_2595),
.Y(n_2825)
);

BUFx4f_ASAP7_75t_L g2826 ( 
.A(n_2732),
.Y(n_2826)
);

AOI22xp33_ASAP7_75t_L g2827 ( 
.A1(n_2724),
.A2(n_2349),
.B1(n_2341),
.B2(n_2348),
.Y(n_2827)
);

INVx1_ASAP7_75t_SL g2828 ( 
.A(n_2606),
.Y(n_2828)
);

CKINVDCx11_ASAP7_75t_R g2829 ( 
.A(n_2684),
.Y(n_2829)
);

INVx3_ASAP7_75t_L g2830 ( 
.A(n_2713),
.Y(n_2830)
);

AND2x4_ASAP7_75t_SL g2831 ( 
.A(n_2537),
.B(n_2284),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_SL g2832 ( 
.A1(n_2648),
.A2(n_2380),
.B1(n_2460),
.B2(n_2287),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2616),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2616),
.Y(n_2834)
);

AOI22xp33_ASAP7_75t_SL g2835 ( 
.A1(n_2648),
.A2(n_2380),
.B1(n_2299),
.B2(n_2312),
.Y(n_2835)
);

AOI22xp33_ASAP7_75t_SL g2836 ( 
.A1(n_2541),
.A2(n_2281),
.B1(n_2368),
.B2(n_2425),
.Y(n_2836)
);

BUFx6f_ASAP7_75t_L g2837 ( 
.A(n_2734),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2555),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2646),
.B(n_2244),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2544),
.B(n_2622),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2568),
.B(n_2285),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_SL g2842 ( 
.A1(n_2541),
.A2(n_2431),
.B1(n_2407),
.B2(n_2412),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2507),
.Y(n_2843)
);

NAND2x1p5_ASAP7_75t_L g2844 ( 
.A(n_2518),
.B(n_2697),
.Y(n_2844)
);

INVx2_ASAP7_75t_SL g2845 ( 
.A(n_2725),
.Y(n_2845)
);

AOI22xp33_ASAP7_75t_SL g2846 ( 
.A1(n_2541),
.A2(n_2701),
.B1(n_2702),
.B2(n_2597),
.Y(n_2846)
);

CKINVDCx6p67_ASAP7_75t_R g2847 ( 
.A(n_2684),
.Y(n_2847)
);

CKINVDCx5p33_ASAP7_75t_R g2848 ( 
.A(n_2725),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2565),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_SL g2850 ( 
.A1(n_2702),
.A2(n_2410),
.B1(n_2435),
.B2(n_2350),
.Y(n_2850)
);

INVx4_ASAP7_75t_L g2851 ( 
.A(n_2677),
.Y(n_2851)
);

CKINVDCx11_ASAP7_75t_R g2852 ( 
.A(n_2684),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2584),
.Y(n_2853)
);

CKINVDCx6p67_ASAP7_75t_R g2854 ( 
.A(n_2483),
.Y(n_2854)
);

AOI22xp33_ASAP7_75t_L g2855 ( 
.A1(n_2552),
.A2(n_2421),
.B1(n_2335),
.B2(n_2338),
.Y(n_2855)
);

BUFx8_ASAP7_75t_SL g2856 ( 
.A(n_2598),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2510),
.Y(n_2857)
);

BUFx2_ASAP7_75t_L g2858 ( 
.A(n_2479),
.Y(n_2858)
);

INVx6_ASAP7_75t_L g2859 ( 
.A(n_2479),
.Y(n_2859)
);

INVx6_ASAP7_75t_L g2860 ( 
.A(n_2479),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2510),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2590),
.Y(n_2862)
);

CKINVDCx6p67_ASAP7_75t_R g2863 ( 
.A(n_2483),
.Y(n_2863)
);

AOI22xp33_ASAP7_75t_L g2864 ( 
.A1(n_2552),
.A2(n_2294),
.B1(n_895),
.B2(n_897),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2552),
.A2(n_896),
.B1(n_899),
.B2(n_897),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_2637),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2690),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2690),
.Y(n_2868)
);

BUFx2_ASAP7_75t_SL g2869 ( 
.A(n_2623),
.Y(n_2869)
);

INVx4_ASAP7_75t_L g2870 ( 
.A(n_2677),
.Y(n_2870)
);

BUFx3_ASAP7_75t_L g2871 ( 
.A(n_2504),
.Y(n_2871)
);

INVx6_ASAP7_75t_L g2872 ( 
.A(n_2687),
.Y(n_2872)
);

INVx4_ASAP7_75t_L g2873 ( 
.A(n_2687),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2622),
.B(n_2311),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2698),
.Y(n_2875)
);

INVx4_ASAP7_75t_L g2876 ( 
.A(n_2687),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2698),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2537),
.A2(n_2260),
.B1(n_2265),
.B2(n_2256),
.Y(n_2878)
);

AOI22xp33_ASAP7_75t_SL g2879 ( 
.A1(n_2597),
.A2(n_2393),
.B1(n_2394),
.B2(n_2392),
.Y(n_2879)
);

AOI22xp33_ASAP7_75t_L g2880 ( 
.A1(n_2552),
.A2(n_899),
.B1(n_2218),
.B2(n_2321),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2592),
.A2(n_2325),
.B1(n_2220),
.B2(n_2308),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_L g2882 ( 
.A1(n_2592),
.A2(n_839),
.B1(n_1041),
.B2(n_1013),
.Y(n_2882)
);

BUFx4f_ASAP7_75t_SL g2883 ( 
.A(n_2504),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2661),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2703),
.Y(n_2885)
);

CKINVDCx11_ASAP7_75t_R g2886 ( 
.A(n_2532),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_L g2887 ( 
.A1(n_2592),
.A2(n_1041),
.B1(n_1013),
.B2(n_1032),
.Y(n_2887)
);

AOI22xp33_ASAP7_75t_SL g2888 ( 
.A1(n_2597),
.A2(n_2331),
.B1(n_4),
.B2(n_2),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2592),
.A2(n_1041),
.B1(n_1013),
.B2(n_1032),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2568),
.B(n_2),
.Y(n_2890)
);

INVx6_ASAP7_75t_L g2891 ( 
.A(n_2537),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2688),
.B(n_3),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2570),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2532),
.A2(n_1041),
.B1(n_1013),
.B2(n_1033),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2734),
.Y(n_2895)
);

AOI22xp33_ASAP7_75t_L g2896 ( 
.A1(n_2532),
.A2(n_1033),
.B1(n_1039),
.B2(n_1027),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2570),
.Y(n_2897)
);

OAI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2615),
.A2(n_2696),
.B1(n_2618),
.B2(n_2705),
.Y(n_2898)
);

INVx2_ASAP7_75t_SL g2899 ( 
.A(n_2623),
.Y(n_2899)
);

AOI22xp33_ASAP7_75t_L g2900 ( 
.A1(n_2532),
.A2(n_1039),
.B1(n_1017),
.B2(n_1018),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2569),
.B(n_3),
.Y(n_2901)
);

AOI22xp33_ASAP7_75t_SL g2902 ( 
.A1(n_2508),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_2667),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2536),
.A2(n_1039),
.B1(n_1017),
.B2(n_1018),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2557),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2548),
.A2(n_1017),
.B1(n_1018),
.B2(n_1016),
.Y(n_2906)
);

AOI22xp33_ASAP7_75t_L g2907 ( 
.A1(n_2536),
.A2(n_1017),
.B1(n_1018),
.B2(n_1016),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2500),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2500),
.Y(n_2909)
);

BUFx12f_ASAP7_75t_L g2910 ( 
.A(n_2604),
.Y(n_2910)
);

AOI22xp33_ASAP7_75t_L g2911 ( 
.A1(n_2502),
.A2(n_1017),
.B1(n_1018),
.B2(n_1016),
.Y(n_2911)
);

OAI22xp33_ASAP7_75t_L g2912 ( 
.A1(n_2601),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_2912)
);

AOI22xp33_ASAP7_75t_L g2913 ( 
.A1(n_2502),
.A2(n_1018),
.B1(n_1025),
.B2(n_1017),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2513),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2513),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2557),
.Y(n_2916)
);

OAI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2618),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2517),
.Y(n_2918)
);

BUFx12f_ASAP7_75t_L g2919 ( 
.A(n_2604),
.Y(n_2919)
);

INVx6_ASAP7_75t_L g2920 ( 
.A(n_2548),
.Y(n_2920)
);

INVx2_ASAP7_75t_SL g2921 ( 
.A(n_2667),
.Y(n_2921)
);

BUFx3_ASAP7_75t_L g2922 ( 
.A(n_2505),
.Y(n_2922)
);

BUFx2_ASAP7_75t_L g2923 ( 
.A(n_2505),
.Y(n_2923)
);

AOI22xp5_ASAP7_75t_SL g2924 ( 
.A1(n_2641),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2517),
.Y(n_2925)
);

CKINVDCx11_ASAP7_75t_R g2926 ( 
.A(n_2676),
.Y(n_2926)
);

INVx2_ASAP7_75t_SL g2927 ( 
.A(n_2711),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2674),
.B(n_14),
.Y(n_2928)
);

CKINVDCx11_ASAP7_75t_R g2929 ( 
.A(n_2676),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2519),
.Y(n_2930)
);

AOI22xp33_ASAP7_75t_L g2931 ( 
.A1(n_2533),
.A2(n_1026),
.B1(n_1034),
.B2(n_1025),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2589),
.Y(n_2932)
);

INVx6_ASAP7_75t_L g2933 ( 
.A(n_2548),
.Y(n_2933)
);

INVx1_ASAP7_75t_SL g2934 ( 
.A(n_2569),
.Y(n_2934)
);

BUFx3_ASAP7_75t_L g2935 ( 
.A(n_2711),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2582),
.B(n_15),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2533),
.A2(n_1026),
.B1(n_1034),
.B2(n_1025),
.Y(n_2937)
);

AOI22xp33_ASAP7_75t_SL g2938 ( 
.A1(n_2601),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_2938)
);

OAI21xp5_ASAP7_75t_SL g2939 ( 
.A1(n_2649),
.A2(n_16),
.B(n_17),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2730),
.A2(n_2598),
.B1(n_2492),
.B2(n_2641),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2519),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2589),
.Y(n_2942)
);

INVx1_ASAP7_75t_SL g2943 ( 
.A(n_2582),
.Y(n_2943)
);

INVx8_ASAP7_75t_L g2944 ( 
.A(n_2635),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2523),
.Y(n_2945)
);

AOI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2601),
.A2(n_1026),
.B1(n_1034),
.B2(n_1025),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2523),
.Y(n_2947)
);

INVx2_ASAP7_75t_SL g2948 ( 
.A(n_2727),
.Y(n_2948)
);

BUFx6f_ASAP7_75t_L g2949 ( 
.A(n_2727),
.Y(n_2949)
);

CKINVDCx20_ASAP7_75t_R g2950 ( 
.A(n_2670),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2605),
.Y(n_2951)
);

CKINVDCx6p67_ASAP7_75t_R g2952 ( 
.A(n_2670),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2562),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2562),
.Y(n_2954)
);

BUFx6f_ASAP7_75t_L g2955 ( 
.A(n_2676),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2605),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2720),
.Y(n_2957)
);

BUFx4_ASAP7_75t_SL g2958 ( 
.A(n_2733),
.Y(n_2958)
);

INVx5_ASAP7_75t_L g2959 ( 
.A(n_2733),
.Y(n_2959)
);

A2O1A1Ixp33_ASAP7_75t_L g2960 ( 
.A1(n_2757),
.A2(n_2717),
.B(n_2599),
.C(n_2497),
.Y(n_2960)
);

HB1xp67_ASAP7_75t_L g2961 ( 
.A(n_2934),
.Y(n_2961)
);

AO21x2_ASAP7_75t_L g2962 ( 
.A1(n_2754),
.A2(n_2549),
.B(n_2477),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2767),
.A2(n_2518),
.B(n_2658),
.Y(n_2963)
);

OAI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2902),
.A2(n_2730),
.B1(n_2497),
.B2(n_2599),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2885),
.B(n_2849),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2853),
.B(n_2674),
.Y(n_2966)
);

AOI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2742),
.A2(n_2805),
.B1(n_2748),
.B2(n_2790),
.Y(n_2967)
);

AOI21x1_ASAP7_75t_L g2968 ( 
.A1(n_2785),
.A2(n_2549),
.B(n_2477),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2743),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2862),
.B(n_2720),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_L g2971 ( 
.A(n_2814),
.B(n_2682),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2755),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2747),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_SL g2974 ( 
.A(n_2750),
.B(n_2601),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2751),
.Y(n_2975)
);

BUFx10_ASAP7_75t_L g2976 ( 
.A(n_2776),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2795),
.B(n_2641),
.Y(n_2977)
);

AOI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2805),
.A2(n_2518),
.B(n_2658),
.Y(n_2978)
);

A2O1A1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_2742),
.A2(n_2697),
.B(n_2635),
.C(n_2673),
.Y(n_2979)
);

OAI22x1_ASAP7_75t_L g2980 ( 
.A1(n_2903),
.A2(n_2736),
.B1(n_2828),
.B2(n_2783),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2762),
.B(n_2723),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2843),
.B(n_2723),
.Y(n_2982)
);

AOI21xp5_ASAP7_75t_L g2983 ( 
.A1(n_2795),
.A2(n_2518),
.B(n_2658),
.Y(n_2983)
);

OA21x2_ASAP7_75t_L g2984 ( 
.A1(n_2754),
.A2(n_2633),
.B(n_2509),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2765),
.Y(n_2985)
);

OAI21x1_ASAP7_75t_L g2986 ( 
.A1(n_2844),
.A2(n_2617),
.B(n_2611),
.Y(n_2986)
);

BUFx2_ASAP7_75t_L g2987 ( 
.A(n_2923),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2893),
.Y(n_2988)
);

AOI222xp33_ASAP7_75t_L g2989 ( 
.A1(n_2939),
.A2(n_2583),
.B1(n_2652),
.B2(n_2614),
.C1(n_2644),
.C2(n_2663),
.Y(n_2989)
);

OA21x2_ASAP7_75t_L g2990 ( 
.A1(n_2784),
.A2(n_2633),
.B(n_2509),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2824),
.A2(n_2518),
.B(n_2697),
.Y(n_2991)
);

OAI21x1_ASAP7_75t_L g2992 ( 
.A1(n_2844),
.A2(n_2617),
.B(n_2611),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2897),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2943),
.B(n_2628),
.Y(n_2994)
);

AOI22xp33_ASAP7_75t_L g2995 ( 
.A1(n_2938),
.A2(n_2650),
.B1(n_2664),
.B2(n_2487),
.Y(n_2995)
);

OAI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2832),
.A2(n_2888),
.B(n_2793),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2902),
.A2(n_2730),
.B1(n_2645),
.B2(n_2726),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2841),
.B(n_2628),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2938),
.A2(n_2650),
.B1(n_2664),
.B2(n_2487),
.Y(n_2999)
);

AOI222xp33_ASAP7_75t_L g3000 ( 
.A1(n_2808),
.A2(n_2583),
.B1(n_2652),
.B2(n_2614),
.C1(n_2663),
.C2(n_2672),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2766),
.Y(n_3001)
);

AO31x2_ASAP7_75t_L g3002 ( 
.A1(n_2940),
.A2(n_2824),
.A3(n_2810),
.B(n_2745),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2840),
.B(n_2659),
.Y(n_3003)
);

AO31x2_ASAP7_75t_L g3004 ( 
.A1(n_2940),
.A2(n_2526),
.A3(n_2546),
.B(n_2501),
.Y(n_3004)
);

AO21x2_ASAP7_75t_L g3005 ( 
.A1(n_2784),
.A2(n_2643),
.B(n_2653),
.Y(n_3005)
);

AO21x2_ASAP7_75t_L g3006 ( 
.A1(n_2890),
.A2(n_2643),
.B(n_2653),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2794),
.Y(n_3007)
);

HB1xp67_ASAP7_75t_L g3008 ( 
.A(n_2763),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2874),
.B(n_2476),
.Y(n_3009)
);

A2O1A1Ixp33_ASAP7_75t_L g3010 ( 
.A1(n_2924),
.A2(n_2738),
.B(n_2888),
.C(n_2832),
.Y(n_3010)
);

OAI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2810),
.A2(n_2630),
.B(n_2668),
.Y(n_3011)
);

AO31x2_ASAP7_75t_L g3012 ( 
.A1(n_2741),
.A2(n_2526),
.A3(n_2546),
.B(n_2501),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2737),
.A2(n_2645),
.B1(n_2726),
.B2(n_2733),
.Y(n_3013)
);

CKINVDCx11_ASAP7_75t_R g3014 ( 
.A(n_2739),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2807),
.A2(n_2697),
.B(n_2710),
.Y(n_3015)
);

AND2x4_ASAP7_75t_L g3016 ( 
.A(n_2763),
.B(n_2697),
.Y(n_3016)
);

AO31x2_ASAP7_75t_L g3017 ( 
.A1(n_2741),
.A2(n_2542),
.A3(n_2543),
.B(n_2534),
.Y(n_3017)
);

OA21x2_ASAP7_75t_L g3018 ( 
.A1(n_2890),
.A2(n_2666),
.B(n_2636),
.Y(n_3018)
);

OA21x2_ASAP7_75t_L g3019 ( 
.A1(n_2928),
.A2(n_2666),
.B(n_2636),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2932),
.Y(n_3020)
);

AOI222xp33_ASAP7_75t_L g3021 ( 
.A1(n_2912),
.A2(n_2672),
.B1(n_2695),
.B2(n_2712),
.C1(n_2706),
.C2(n_2686),
.Y(n_3021)
);

OAI21x1_ASAP7_75t_L g3022 ( 
.A1(n_2931),
.A2(n_2630),
.B(n_2668),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2841),
.B(n_2639),
.Y(n_3023)
);

AO21x2_ASAP7_75t_L g3024 ( 
.A1(n_2912),
.A2(n_2643),
.B(n_2572),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2942),
.Y(n_3025)
);

AOI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2778),
.A2(n_2697),
.B(n_2710),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2773),
.Y(n_3027)
);

HB1xp67_ASAP7_75t_L g3028 ( 
.A(n_2857),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2951),
.Y(n_3029)
);

HB1xp67_ASAP7_75t_L g3030 ( 
.A(n_2861),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2746),
.B(n_2476),
.Y(n_3031)
);

OR2x2_ASAP7_75t_L g3032 ( 
.A(n_2775),
.B(n_2659),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2777),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2871),
.B(n_2476),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2787),
.Y(n_3035)
);

CKINVDCx5p33_ASAP7_75t_R g3036 ( 
.A(n_2764),
.Y(n_3036)
);

A2O1A1Ixp33_ASAP7_75t_L g3037 ( 
.A1(n_2846),
.A2(n_2635),
.B(n_2673),
.C(n_2530),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2956),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2789),
.B(n_2639),
.Y(n_3039)
);

AOI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2778),
.A2(n_2710),
.B(n_2714),
.Y(n_3040)
);

AOI21x1_ASAP7_75t_L g3041 ( 
.A1(n_2785),
.A2(n_2695),
.B(n_2704),
.Y(n_3041)
);

AOI21xp5_ASAP7_75t_L g3042 ( 
.A1(n_2839),
.A2(n_2722),
.B(n_2714),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2819),
.Y(n_3043)
);

HB1xp67_ASAP7_75t_L g3044 ( 
.A(n_2905),
.Y(n_3044)
);

AOI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2839),
.A2(n_2846),
.B(n_2865),
.Y(n_3045)
);

OAI21x1_ASAP7_75t_L g3046 ( 
.A1(n_2937),
.A2(n_2707),
.B(n_2700),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2796),
.Y(n_3047)
);

AOI221xp5_ASAP7_75t_L g3048 ( 
.A1(n_2917),
.A2(n_2706),
.B1(n_2719),
.B2(n_2686),
.C(n_2625),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2798),
.B(n_2640),
.Y(n_3049)
);

OR2x2_ASAP7_75t_L g3050 ( 
.A(n_2812),
.B(n_2482),
.Y(n_3050)
);

OAI21x1_ASAP7_75t_SL g3051 ( 
.A1(n_2928),
.A2(n_2760),
.B(n_2745),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2816),
.Y(n_3052)
);

AO21x2_ASAP7_75t_L g3053 ( 
.A1(n_2833),
.A2(n_2572),
.B(n_2588),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2959),
.A2(n_2782),
.B(n_2864),
.Y(n_3054)
);

OAI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2854),
.A2(n_2733),
.B1(n_2596),
.B2(n_2645),
.Y(n_3055)
);

INVx4_ASAP7_75t_L g3056 ( 
.A(n_2847),
.Y(n_3056)
);

AOI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_2910),
.A2(n_2650),
.B1(n_2664),
.B2(n_2487),
.Y(n_3057)
);

HB1xp67_ASAP7_75t_L g3058 ( 
.A(n_2916),
.Y(n_3058)
);

AO21x2_ASAP7_75t_L g3059 ( 
.A1(n_2834),
.A2(n_2593),
.B(n_2588),
.Y(n_3059)
);

OAI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2835),
.A2(n_2721),
.B(n_2475),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2867),
.B(n_2640),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2838),
.Y(n_3062)
);

BUFx6f_ASAP7_75t_L g3063 ( 
.A(n_2821),
.Y(n_3063)
);

AOI21x1_ASAP7_75t_L g3064 ( 
.A1(n_2744),
.A2(n_2728),
.B(n_2638),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2868),
.B(n_2669),
.Y(n_3065)
);

OAI221xp5_ASAP7_75t_L g3066 ( 
.A1(n_2753),
.A2(n_2733),
.B1(n_2726),
.B2(n_2719),
.C(n_2625),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2875),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2877),
.Y(n_3068)
);

BUFx3_ASAP7_75t_L g3069 ( 
.A(n_2780),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2957),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2908),
.B(n_2669),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2909),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_SL g3073 ( 
.A(n_2786),
.B(n_2676),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2922),
.B(n_2482),
.Y(n_3074)
);

INVx3_ASAP7_75t_L g3075 ( 
.A(n_2935),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2914),
.Y(n_3076)
);

OAI22x1_ASAP7_75t_L g3077 ( 
.A1(n_2736),
.A2(n_2482),
.B1(n_2494),
.B2(n_2591),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2915),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2959),
.A2(n_2722),
.B(n_2714),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2918),
.B(n_2671),
.Y(n_3080)
);

A2O1A1Ixp33_ASAP7_75t_L g3081 ( 
.A1(n_2781),
.A2(n_2898),
.B(n_2761),
.C(n_2771),
.Y(n_3081)
);

OAI21x1_ASAP7_75t_L g3082 ( 
.A1(n_2804),
.A2(n_2707),
.B(n_2700),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2925),
.B(n_2671),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2930),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2959),
.A2(n_2722),
.B(n_2593),
.Y(n_3085)
);

A2O1A1Ixp33_ASAP7_75t_L g3086 ( 
.A1(n_2898),
.A2(n_2673),
.B(n_2635),
.C(n_2530),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_2863),
.B(n_2494),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2941),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2945),
.B(n_2716),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2947),
.B(n_2716),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2953),
.B(n_2662),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2954),
.B(n_2662),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2869),
.Y(n_3093)
);

OA21x2_ASAP7_75t_L g3094 ( 
.A1(n_2756),
.A2(n_2559),
.B(n_2551),
.Y(n_3094)
);

OAI21xp33_ASAP7_75t_L g3095 ( 
.A1(n_2836),
.A2(n_2495),
.B(n_2478),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2899),
.Y(n_3096)
);

OAI21x1_ASAP7_75t_L g3097 ( 
.A1(n_2804),
.A2(n_2559),
.B(n_2551),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2921),
.B(n_2494),
.Y(n_3098)
);

AO21x2_ASAP7_75t_L g3099 ( 
.A1(n_2769),
.A2(n_2593),
.B(n_2588),
.Y(n_3099)
);

OAI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_2917),
.A2(n_2596),
.B1(n_2474),
.B2(n_2558),
.Y(n_3100)
);

OA21x2_ASAP7_75t_L g3101 ( 
.A1(n_2749),
.A2(n_2527),
.B(n_2528),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2836),
.B(n_2694),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2959),
.A2(n_2709),
.B(n_2683),
.Y(n_3103)
);

BUFx2_ASAP7_75t_L g3104 ( 
.A(n_2856),
.Y(n_3104)
);

BUFx2_ASAP7_75t_L g3105 ( 
.A(n_2774),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2830),
.B(n_2591),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2842),
.B(n_2694),
.Y(n_3107)
);

OA21x2_ASAP7_75t_L g3108 ( 
.A1(n_2827),
.A2(n_2527),
.B(n_2528),
.Y(n_3108)
);

AOI221xp5_ASAP7_75t_L g3109 ( 
.A1(n_2744),
.A2(n_2495),
.B1(n_2478),
.B2(n_2708),
.C(n_2542),
.Y(n_3109)
);

NAND2x1p5_ASAP7_75t_L g3110 ( 
.A(n_2760),
.B(n_2553),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2858),
.B(n_2591),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2782),
.A2(n_2709),
.B(n_2683),
.Y(n_3112)
);

OAI211xp5_ASAP7_75t_L g3113 ( 
.A1(n_2835),
.A2(n_2708),
.B(n_2512),
.C(n_2531),
.Y(n_3113)
);

OAI21x1_ASAP7_75t_SL g3114 ( 
.A1(n_2820),
.A2(n_2531),
.B(n_2512),
.Y(n_3114)
);

AND2x4_ASAP7_75t_L g3115 ( 
.A(n_2830),
.B(n_2534),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_L g3116 ( 
.A1(n_2919),
.A2(n_2487),
.B1(n_2664),
.B2(n_2650),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2803),
.Y(n_3117)
);

OAI22xp33_ASAP7_75t_SL g3118 ( 
.A1(n_2759),
.A2(n_2596),
.B1(n_2474),
.B2(n_2538),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2842),
.B(n_2620),
.Y(n_3119)
);

AOI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_2944),
.A2(n_2709),
.B(n_2683),
.Y(n_3120)
);

OR2x2_ASAP7_75t_L g3121 ( 
.A(n_2927),
.B(n_2481),
.Y(n_3121)
);

OAI21x1_ASAP7_75t_L g3122 ( 
.A1(n_2855),
.A2(n_2619),
.B(n_2486),
.Y(n_3122)
);

OAI22xp5_ASAP7_75t_SL g3123 ( 
.A1(n_2799),
.A2(n_2596),
.B1(n_2474),
.B2(n_2673),
.Y(n_3123)
);

OAI21x1_ASAP7_75t_L g3124 ( 
.A1(n_2881),
.A2(n_2619),
.B(n_2486),
.Y(n_3124)
);

OAI21x1_ASAP7_75t_L g3125 ( 
.A1(n_2906),
.A2(n_2490),
.B(n_2560),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2879),
.B(n_2620),
.Y(n_3126)
);

OA21x2_ASAP7_75t_L g3127 ( 
.A1(n_2768),
.A2(n_2770),
.B(n_2800),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2879),
.B(n_2481),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2948),
.Y(n_3129)
);

A2O1A1Ixp33_ASAP7_75t_L g3130 ( 
.A1(n_2771),
.A2(n_2530),
.B(n_2650),
.C(n_2487),
.Y(n_3130)
);

INVx5_ASAP7_75t_L g3131 ( 
.A(n_2759),
.Y(n_3131)
);

NAND3xp33_ASAP7_75t_L g3132 ( 
.A(n_2850),
.B(n_2545),
.C(n_2543),
.Y(n_3132)
);

OAI21x1_ASAP7_75t_L g3133 ( 
.A1(n_2878),
.A2(n_2490),
.B(n_2560),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2803),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_SL g3135 ( 
.A1(n_2786),
.A2(n_2759),
.B1(n_2772),
.B2(n_2818),
.Y(n_3135)
);

AO31x2_ASAP7_75t_L g3136 ( 
.A1(n_2820),
.A2(n_2547),
.A3(n_2545),
.B(n_2484),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2803),
.Y(n_3137)
);

OAI22xp33_ASAP7_75t_L g3138 ( 
.A1(n_2823),
.A2(n_2596),
.B1(n_2474),
.B2(n_2664),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2811),
.Y(n_3139)
);

OAI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_2850),
.A2(n_2475),
.B(n_2530),
.Y(n_3140)
);

AND2x6_ASAP7_75t_SL g3141 ( 
.A(n_2792),
.B(n_2474),
.Y(n_3141)
);

AOI22xp33_ASAP7_75t_L g3142 ( 
.A1(n_2886),
.A2(n_2676),
.B1(n_2692),
.B2(n_2554),
.Y(n_3142)
);

INVx2_ASAP7_75t_SL g3143 ( 
.A(n_2740),
.Y(n_3143)
);

OAI221xp5_ASAP7_75t_SL g3144 ( 
.A1(n_2752),
.A2(n_2547),
.B1(n_2493),
.B2(n_2489),
.C(n_2484),
.Y(n_3144)
);

A2O1A1Ixp33_ASAP7_75t_L g3145 ( 
.A1(n_2826),
.A2(n_2553),
.B(n_2647),
.C(n_2516),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2809),
.B(n_2489),
.Y(n_3146)
);

OA21x2_ASAP7_75t_L g3147 ( 
.A1(n_2901),
.A2(n_2693),
.B(n_2665),
.Y(n_3147)
);

AOI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2944),
.A2(n_2558),
.B(n_2638),
.Y(n_3148)
);

OAI221xp5_ASAP7_75t_L g3149 ( 
.A1(n_2788),
.A2(n_2578),
.B1(n_2600),
.B2(n_2585),
.C(n_2580),
.Y(n_3149)
);

INVx3_ASAP7_75t_L g3150 ( 
.A(n_2872),
.Y(n_3150)
);

OAI21xp33_ASAP7_75t_L g3151 ( 
.A1(n_3010),
.A2(n_2806),
.B(n_2809),
.Y(n_3151)
);

INVx8_ASAP7_75t_L g3152 ( 
.A(n_3063),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_3063),
.B(n_2883),
.Y(n_3153)
);

AOI21xp33_ASAP7_75t_L g3154 ( 
.A1(n_2996),
.A2(n_2936),
.B(n_2892),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_2996),
.A2(n_2788),
.B1(n_2806),
.B2(n_2772),
.Y(n_3155)
);

AOI22xp33_ASAP7_75t_L g3156 ( 
.A1(n_2967),
.A2(n_2772),
.B1(n_2859),
.B2(n_2822),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_3013),
.A2(n_2822),
.B1(n_2860),
.B2(n_2859),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2969),
.Y(n_3158)
);

AOI21x1_ASAP7_75t_L g3159 ( 
.A1(n_3041),
.A2(n_2728),
.B(n_2638),
.Y(n_3159)
);

AOI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_3013),
.A2(n_2822),
.B1(n_2860),
.B2(n_2859),
.Y(n_3160)
);

INVx4_ASAP7_75t_L g3161 ( 
.A(n_3063),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2973),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2987),
.B(n_2797),
.Y(n_3163)
);

AOI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_2963),
.A2(n_2826),
.B(n_2944),
.Y(n_3164)
);

OR2x6_ASAP7_75t_L g3165 ( 
.A(n_2983),
.B(n_2860),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2975),
.Y(n_3166)
);

AO31x2_ASAP7_75t_L g3167 ( 
.A1(n_3079),
.A2(n_2870),
.A3(n_2873),
.B(n_2851),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_3001),
.Y(n_3168)
);

AOI221xp5_ASAP7_75t_L g3169 ( 
.A1(n_3081),
.A2(n_2758),
.B1(n_2880),
.B2(n_2845),
.C(n_2802),
.Y(n_3169)
);

BUFx3_ASAP7_75t_L g3170 ( 
.A(n_3014),
.Y(n_3170)
);

OAI22xp5_ASAP7_75t_L g3171 ( 
.A1(n_2960),
.A2(n_2750),
.B1(n_2950),
.B2(n_2884),
.Y(n_3171)
);

AO221x1_ASAP7_75t_L g3172 ( 
.A1(n_3077),
.A2(n_2813),
.B1(n_2811),
.B2(n_2955),
.C(n_2895),
.Y(n_3172)
);

HB1xp67_ASAP7_75t_L g3173 ( 
.A(n_2961),
.Y(n_3173)
);

INVx3_ASAP7_75t_L g3174 ( 
.A(n_3150),
.Y(n_3174)
);

AOI22xp33_ASAP7_75t_L g3175 ( 
.A1(n_3127),
.A2(n_2891),
.B1(n_2933),
.B2(n_2920),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_3150),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_SL g3177 ( 
.A1(n_2997),
.A2(n_2891),
.B1(n_2933),
.B2(n_2920),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_3056),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3027),
.Y(n_3179)
);

INVx2_ASAP7_75t_L g3180 ( 
.A(n_2972),
.Y(n_3180)
);

AOI22xp33_ASAP7_75t_L g3181 ( 
.A1(n_3127),
.A2(n_2891),
.B1(n_2933),
.B2(n_2920),
.Y(n_3181)
);

NAND2xp33_ASAP7_75t_SL g3182 ( 
.A(n_2980),
.B(n_2866),
.Y(n_3182)
);

OAI21x1_ASAP7_75t_L g3183 ( 
.A1(n_2991),
.A2(n_2638),
.B(n_2728),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_SL g3184 ( 
.A1(n_2997),
.A2(n_2831),
.B1(n_2735),
.B2(n_2801),
.Y(n_3184)
);

AOI22xp33_ASAP7_75t_L g3185 ( 
.A1(n_3054),
.A2(n_2815),
.B1(n_2852),
.B2(n_2829),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3033),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_2964),
.A2(n_2825),
.B1(n_2889),
.B2(n_2887),
.Y(n_3187)
);

INVx6_ASAP7_75t_L g3188 ( 
.A(n_2976),
.Y(n_3188)
);

AOI22xp33_ASAP7_75t_SL g3189 ( 
.A1(n_2964),
.A2(n_3066),
.B1(n_2974),
.B2(n_2978),
.Y(n_3189)
);

BUFx6f_ASAP7_75t_L g3190 ( 
.A(n_2976),
.Y(n_3190)
);

AOI22xp5_ASAP7_75t_L g3191 ( 
.A1(n_3123),
.A2(n_2872),
.B1(n_2952),
.B2(n_2791),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3035),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3047),
.Y(n_3193)
);

OAI22xp5_ASAP7_75t_L g3194 ( 
.A1(n_2995),
.A2(n_2553),
.B1(n_2779),
.B2(n_2848),
.Y(n_3194)
);

AOI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_3138),
.A2(n_2882),
.B1(n_2735),
.B2(n_2801),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2965),
.B(n_2966),
.Y(n_3196)
);

OR2x2_ASAP7_75t_L g3197 ( 
.A(n_3003),
.B(n_2493),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3052),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3067),
.Y(n_3199)
);

INVx6_ASAP7_75t_L g3200 ( 
.A(n_3056),
.Y(n_3200)
);

OAI221xp5_ASAP7_75t_L g3201 ( 
.A1(n_2979),
.A2(n_2872),
.B1(n_2873),
.B2(n_2870),
.C(n_2851),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_2977),
.A2(n_2692),
.B1(n_2647),
.B2(n_2554),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_2985),
.Y(n_3203)
);

AOI22xp33_ASAP7_75t_L g3204 ( 
.A1(n_2999),
.A2(n_2692),
.B1(n_2647),
.B2(n_2554),
.Y(n_3204)
);

AOI22xp33_ASAP7_75t_L g3205 ( 
.A1(n_2989),
.A2(n_2692),
.B1(n_2895),
.B2(n_2837),
.Y(n_3205)
);

OAI33xp33_ASAP7_75t_L g3206 ( 
.A1(n_2965),
.A2(n_20),
.A3(n_23),
.B1(n_18),
.B2(n_19),
.B3(n_22),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_3009),
.B(n_2817),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_3031),
.B(n_2817),
.Y(n_3208)
);

OAI211xp5_ASAP7_75t_L g3209 ( 
.A1(n_2989),
.A2(n_2929),
.B(n_2926),
.C(n_2907),
.Y(n_3209)
);

AOI22xp33_ASAP7_75t_L g3210 ( 
.A1(n_3045),
.A2(n_2692),
.B1(n_2895),
.B2(n_2837),
.Y(n_3210)
);

AOI22xp33_ASAP7_75t_L g3211 ( 
.A1(n_3000),
.A2(n_2949),
.B1(n_2837),
.B2(n_2876),
.Y(n_3211)
);

AOI221xp5_ASAP7_75t_L g3212 ( 
.A1(n_3095),
.A2(n_2949),
.B1(n_2904),
.B2(n_2520),
.C(n_2516),
.Y(n_3212)
);

AOI22xp33_ASAP7_75t_L g3213 ( 
.A1(n_3000),
.A2(n_2949),
.B1(n_2876),
.B2(n_2580),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2966),
.B(n_2728),
.Y(n_3214)
);

AOI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_3105),
.A2(n_2585),
.B1(n_2600),
.B2(n_2578),
.Y(n_3215)
);

AND2x6_ASAP7_75t_L g3216 ( 
.A(n_3087),
.B(n_2958),
.Y(n_3216)
);

AND2x2_ASAP7_75t_L g3217 ( 
.A(n_3008),
.B(n_2811),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_3111),
.B(n_2813),
.Y(n_3218)
);

AND2x2_ASAP7_75t_L g3219 ( 
.A(n_3098),
.B(n_2813),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3007),
.Y(n_3220)
);

AOI222xp33_ASAP7_75t_SL g3221 ( 
.A1(n_3100),
.A2(n_24),
.B1(n_26),
.B2(n_20),
.C1(n_23),
.C2(n_25),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3068),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3076),
.Y(n_3223)
);

AOI22xp33_ASAP7_75t_L g3224 ( 
.A1(n_3021),
.A2(n_2602),
.B1(n_2681),
.B2(n_2516),
.Y(n_3224)
);

AND2x2_ASAP7_75t_L g3225 ( 
.A(n_3034),
.B(n_2955),
.Y(n_3225)
);

OAI21x1_ASAP7_75t_L g3226 ( 
.A1(n_3015),
.A2(n_2678),
.B(n_2520),
.Y(n_3226)
);

OAI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_3086),
.A2(n_2475),
.B1(n_2558),
.B2(n_2538),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3021),
.A2(n_2602),
.B1(n_2681),
.B2(n_2520),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_3051),
.A2(n_2681),
.B1(n_2514),
.B2(n_2538),
.Y(n_3229)
);

INVx2_ASAP7_75t_SL g3230 ( 
.A(n_3143),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_3078),
.Y(n_3231)
);

OAI21xp33_ASAP7_75t_SL g3232 ( 
.A1(n_3073),
.A2(n_2958),
.B(n_2514),
.Y(n_3232)
);

AOI22xp33_ASAP7_75t_L g3233 ( 
.A1(n_3055),
.A2(n_2514),
.B1(n_2535),
.B2(n_2499),
.Y(n_3233)
);

O2A1O1Ixp33_ASAP7_75t_L g3234 ( 
.A1(n_3112),
.A2(n_2680),
.B(n_2535),
.C(n_2626),
.Y(n_3234)
);

OAI22xp5_ASAP7_75t_L g3235 ( 
.A1(n_3037),
.A2(n_2558),
.B1(n_2535),
.B2(n_2900),
.Y(n_3235)
);

OAI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_2974),
.A2(n_2680),
.B1(n_2626),
.B2(n_2955),
.Y(n_3236)
);

AOI22xp33_ASAP7_75t_L g3237 ( 
.A1(n_3099),
.A2(n_2499),
.B1(n_2629),
.B2(n_2594),
.Y(n_3237)
);

INVx2_ASAP7_75t_SL g3238 ( 
.A(n_3075),
.Y(n_3238)
);

OAI222xp33_ASAP7_75t_L g3239 ( 
.A1(n_3135),
.A2(n_2680),
.B1(n_2626),
.B2(n_2946),
.C1(n_2913),
.C2(n_2911),
.Y(n_3239)
);

OAI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_3132),
.A2(n_2678),
.B1(n_2896),
.B2(n_2894),
.Y(n_3240)
);

OAI221xp5_ASAP7_75t_L g3241 ( 
.A1(n_3140),
.A2(n_2678),
.B1(n_2685),
.B2(n_28),
.C(n_24),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3074),
.B(n_2678),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_3099),
.A2(n_2499),
.B1(n_2629),
.B2(n_2594),
.Y(n_3243)
);

OAI221xp5_ASAP7_75t_L g3244 ( 
.A1(n_3130),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.C(n_31),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2971),
.A2(n_2629),
.B1(n_2594),
.B2(n_2571),
.Y(n_3245)
);

HB1xp67_ASAP7_75t_L g3246 ( 
.A(n_3028),
.Y(n_3246)
);

OAI221xp5_ASAP7_75t_L g3247 ( 
.A1(n_3140),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.C(n_35),
.Y(n_3247)
);

CKINVDCx5p33_ASAP7_75t_R g3248 ( 
.A(n_3036),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3020),
.B(n_2529),
.Y(n_3249)
);

AOI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_3042),
.A2(n_2571),
.B(n_2529),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3025),
.B(n_2529),
.Y(n_3251)
);

AOI22xp33_ASAP7_75t_SL g3252 ( 
.A1(n_3100),
.A2(n_2571),
.B1(n_2521),
.B2(n_2632),
.Y(n_3252)
);

OAI33xp33_ASAP7_75t_L g3253 ( 
.A1(n_2970),
.A2(n_36),
.A3(n_38),
.B1(n_34),
.B2(n_35),
.B3(n_37),
.Y(n_3253)
);

OAI221xp5_ASAP7_75t_L g3254 ( 
.A1(n_3060),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.C(n_40),
.Y(n_3254)
);

OA21x2_ASAP7_75t_L g3255 ( 
.A1(n_3107),
.A2(n_2693),
.B(n_2665),
.Y(n_3255)
);

AND2x4_ASAP7_75t_L g3256 ( 
.A(n_3106),
.B(n_2521),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_3137),
.Y(n_3257)
);

AOI21xp33_ASAP7_75t_L g3258 ( 
.A1(n_3048),
.A2(n_40),
.B(n_41),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_SL g3259 ( 
.A1(n_3118),
.A2(n_2521),
.B1(n_2632),
.B2(n_2731),
.Y(n_3259)
);

AOI221xp5_ASAP7_75t_L g3260 ( 
.A1(n_3144),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.C(n_45),
.Y(n_3260)
);

AOI22xp33_ASAP7_75t_L g3261 ( 
.A1(n_3060),
.A2(n_2632),
.B1(n_2627),
.B2(n_2729),
.Y(n_3261)
);

AOI22xp33_ASAP7_75t_L g3262 ( 
.A1(n_3149),
.A2(n_2627),
.B1(n_2729),
.B2(n_2491),
.Y(n_3262)
);

BUFx6f_ASAP7_75t_L g3263 ( 
.A(n_3104),
.Y(n_3263)
);

INVx2_ASAP7_75t_SL g3264 ( 
.A(n_3075),
.Y(n_3264)
);

INVx5_ASAP7_75t_SL g3265 ( 
.A(n_3006),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3139),
.Y(n_3266)
);

BUFx2_ASAP7_75t_L g3267 ( 
.A(n_3106),
.Y(n_3267)
);

AOI21xp33_ASAP7_75t_L g3268 ( 
.A1(n_2962),
.A2(n_42),
.B(n_43),
.Y(n_3268)
);

AOI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_3093),
.A2(n_3024),
.B1(n_3109),
.B2(n_3057),
.Y(n_3269)
);

OAI21x1_ASAP7_75t_L g3270 ( 
.A1(n_3026),
.A2(n_2587),
.B(n_2524),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_3024),
.A2(n_2491),
.B1(n_2731),
.B2(n_2631),
.Y(n_3271)
);

OR2x2_ASAP7_75t_L g3272 ( 
.A(n_3032),
.B(n_2587),
.Y(n_3272)
);

AOI22xp33_ASAP7_75t_L g3273 ( 
.A1(n_3116),
.A2(n_2631),
.B1(n_2524),
.B2(n_1026),
.Y(n_3273)
);

INVx2_ASAP7_75t_SL g3274 ( 
.A(n_3117),
.Y(n_3274)
);

INVx6_ASAP7_75t_L g3275 ( 
.A(n_3069),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_2968),
.A2(n_2624),
.B1(n_47),
.B2(n_44),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2988),
.Y(n_3277)
);

OAI221xp5_ASAP7_75t_L g3278 ( 
.A1(n_3145),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.C(n_49),
.Y(n_3278)
);

OAI221xp5_ASAP7_75t_SL g3279 ( 
.A1(n_3113),
.A2(n_54),
.B1(n_46),
.B2(n_51),
.C(n_56),
.Y(n_3279)
);

AOI221xp5_ASAP7_75t_L g3280 ( 
.A1(n_3102),
.A2(n_56),
.B1(n_51),
.B2(n_54),
.C(n_57),
.Y(n_3280)
);

OAI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_3131),
.A2(n_2624),
.B1(n_60),
.B2(n_58),
.Y(n_3281)
);

AOI22xp33_ASAP7_75t_L g3282 ( 
.A1(n_3006),
.A2(n_1026),
.B1(n_1034),
.B2(n_1025),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3084),
.Y(n_3283)
);

AOI22xp33_ASAP7_75t_L g3284 ( 
.A1(n_3146),
.A2(n_1026),
.B1(n_1034),
.B2(n_1025),
.Y(n_3284)
);

INVx2_ASAP7_75t_L g3285 ( 
.A(n_2993),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_3146),
.A2(n_1036),
.B1(n_1040),
.B2(n_1034),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3088),
.Y(n_3287)
);

OAI221xp5_ASAP7_75t_L g3288 ( 
.A1(n_3102),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.C(n_63),
.Y(n_3288)
);

OAI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_3040),
.A2(n_63),
.B(n_64),
.Y(n_3289)
);

OAI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_3142),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_3290)
);

OAI211xp5_ASAP7_75t_L g3291 ( 
.A1(n_3128),
.A2(n_68),
.B(n_65),
.C(n_66),
.Y(n_3291)
);

AOI221xp5_ASAP7_75t_L g3292 ( 
.A1(n_3128),
.A2(n_73),
.B1(n_68),
.B2(n_72),
.C(n_74),
.Y(n_3292)
);

AOI211xp5_ASAP7_75t_L g3293 ( 
.A1(n_3096),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3120),
.A2(n_1040),
.B1(n_1036),
.B2(n_1119),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3070),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_3085),
.A2(n_1040),
.B(n_1036),
.Y(n_3296)
);

OAI21x1_ASAP7_75t_L g3297 ( 
.A1(n_3148),
.A2(n_941),
.B(n_938),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3016),
.A2(n_3129),
.B1(n_3131),
.B2(n_3126),
.Y(n_3298)
);

OAI22xp33_ASAP7_75t_L g3299 ( 
.A1(n_3131),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3299)
);

OR2x6_ASAP7_75t_L g3300 ( 
.A(n_3103),
.B(n_1036),
.Y(n_3300)
);

INVx3_ASAP7_75t_L g3301 ( 
.A(n_3016),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_3131),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_3302)
);

AND2x4_ASAP7_75t_L g3303 ( 
.A(n_3134),
.B(n_78),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3072),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2970),
.Y(n_3305)
);

INVx2_ASAP7_75t_SL g3306 ( 
.A(n_3121),
.Y(n_3306)
);

OAI22xp5_ASAP7_75t_L g3307 ( 
.A1(n_3126),
.A2(n_82),
.B1(n_79),
.B2(n_80),
.Y(n_3307)
);

AND2x4_ASAP7_75t_L g3308 ( 
.A(n_3115),
.B(n_3012),
.Y(n_3308)
);

AOI22xp33_ASAP7_75t_L g3309 ( 
.A1(n_2962),
.A2(n_1040),
.B1(n_1036),
.B2(n_1119),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3158),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3162),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3301),
.B(n_3002),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_3308),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_3166),
.Y(n_3314)
);

HB1xp67_ASAP7_75t_L g3315 ( 
.A(n_3246),
.Y(n_3315)
);

HB1xp67_ASAP7_75t_L g3316 ( 
.A(n_3173),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3168),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3308),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3301),
.B(n_3002),
.Y(n_3319)
);

AND2x2_ASAP7_75t_L g3320 ( 
.A(n_3267),
.B(n_3002),
.Y(n_3320)
);

AND2x4_ASAP7_75t_SL g3321 ( 
.A(n_3190),
.B(n_3030),
.Y(n_3321)
);

AO21x2_ASAP7_75t_L g3322 ( 
.A1(n_3289),
.A2(n_3268),
.B(n_3296),
.Y(n_3322)
);

INVxp67_ASAP7_75t_SL g3323 ( 
.A(n_3196),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3207),
.B(n_3004),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3179),
.Y(n_3325)
);

AOI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_3221),
.A2(n_3107),
.B1(n_3119),
.B2(n_3053),
.Y(n_3326)
);

INVx3_ASAP7_75t_SL g3327 ( 
.A(n_3152),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3186),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3277),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3208),
.B(n_3004),
.Y(n_3330)
);

OR2x2_ASAP7_75t_L g3331 ( 
.A(n_3196),
.B(n_3004),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3305),
.B(n_3044),
.Y(n_3332)
);

BUFx2_ASAP7_75t_L g3333 ( 
.A(n_3165),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3192),
.Y(n_3334)
);

OR2x2_ASAP7_75t_L g3335 ( 
.A(n_3306),
.B(n_3119),
.Y(n_3335)
);

AND2x4_ASAP7_75t_SL g3336 ( 
.A(n_3190),
.B(n_3058),
.Y(n_3336)
);

OR2x2_ASAP7_75t_L g3337 ( 
.A(n_3197),
.B(n_2994),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_3214),
.B(n_2994),
.Y(n_3338)
);

AND2x4_ASAP7_75t_SL g3339 ( 
.A(n_3190),
.B(n_3115),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3193),
.Y(n_3340)
);

BUFx3_ASAP7_75t_L g3341 ( 
.A(n_3152),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3285),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3269),
.B(n_2998),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3198),
.Y(n_3344)
);

INVxp67_ASAP7_75t_L g3345 ( 
.A(n_3199),
.Y(n_3345)
);

AND2x4_ASAP7_75t_L g3346 ( 
.A(n_3165),
.B(n_3012),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_3174),
.B(n_3019),
.Y(n_3347)
);

BUFx2_ASAP7_75t_L g3348 ( 
.A(n_3165),
.Y(n_3348)
);

AND2x4_ASAP7_75t_L g3349 ( 
.A(n_3167),
.B(n_3012),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3174),
.B(n_3019),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3222),
.Y(n_3351)
);

OAI211xp5_ASAP7_75t_L g3352 ( 
.A1(n_3151),
.A2(n_2982),
.B(n_3023),
.C(n_2998),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3223),
.Y(n_3353)
);

HB1xp67_ASAP7_75t_L g3354 ( 
.A(n_3295),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_L g3355 ( 
.A(n_3188),
.B(n_3141),
.Y(n_3355)
);

AND2x4_ASAP7_75t_L g3356 ( 
.A(n_3167),
.B(n_3017),
.Y(n_3356)
);

AND2x2_ASAP7_75t_L g3357 ( 
.A(n_3176),
.B(n_3018),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3231),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_3176),
.B(n_3018),
.Y(n_3359)
);

AND2x4_ASAP7_75t_L g3360 ( 
.A(n_3167),
.B(n_3017),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3283),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3287),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3304),
.Y(n_3363)
);

AND2x2_ASAP7_75t_L g3364 ( 
.A(n_3217),
.B(n_3029),
.Y(n_3364)
);

AOI21xp33_ASAP7_75t_L g3365 ( 
.A1(n_3289),
.A2(n_3114),
.B(n_2982),
.Y(n_3365)
);

BUFx2_ASAP7_75t_L g3366 ( 
.A(n_3232),
.Y(n_3366)
);

HB1xp67_ASAP7_75t_L g3367 ( 
.A(n_3180),
.Y(n_3367)
);

OR2x2_ASAP7_75t_L g3368 ( 
.A(n_3214),
.B(n_3050),
.Y(n_3368)
);

NAND2x1_ASAP7_75t_L g3369 ( 
.A(n_3172),
.B(n_2984),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3203),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3220),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3257),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3218),
.B(n_3038),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3266),
.Y(n_3374)
);

INVx3_ASAP7_75t_L g3375 ( 
.A(n_3200),
.Y(n_3375)
);

BUFx2_ASAP7_75t_L g3376 ( 
.A(n_3216),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3242),
.B(n_3023),
.Y(n_3377)
);

INVxp67_ASAP7_75t_L g3378 ( 
.A(n_3182),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3272),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3249),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3225),
.B(n_3043),
.Y(n_3381)
);

BUFx2_ASAP7_75t_L g3382 ( 
.A(n_3216),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_3219),
.B(n_3238),
.Y(n_3383)
);

OR2x2_ASAP7_75t_L g3384 ( 
.A(n_3265),
.B(n_3062),
.Y(n_3384)
);

NOR4xp25_ASAP7_75t_SL g3385 ( 
.A(n_3201),
.B(n_3064),
.C(n_3110),
.D(n_2984),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3264),
.B(n_2990),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3175),
.B(n_2981),
.Y(n_3387)
);

INVx2_ASAP7_75t_L g3388 ( 
.A(n_3265),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3265),
.Y(n_3389)
);

HB1xp67_ASAP7_75t_L g3390 ( 
.A(n_3249),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3251),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_3256),
.Y(n_3392)
);

INVx3_ASAP7_75t_L g3393 ( 
.A(n_3200),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3251),
.Y(n_3394)
);

BUFx2_ASAP7_75t_L g3395 ( 
.A(n_3216),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_SL g3396 ( 
.A1(n_3247),
.A2(n_3110),
.B1(n_2990),
.B2(n_3053),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3163),
.B(n_3017),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3181),
.B(n_3210),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3274),
.Y(n_3399)
);

BUFx2_ASAP7_75t_L g3400 ( 
.A(n_3216),
.Y(n_3400)
);

AND2x4_ASAP7_75t_SL g3401 ( 
.A(n_3178),
.B(n_3161),
.Y(n_3401)
);

INVx1_ASAP7_75t_SL g3402 ( 
.A(n_3170),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3256),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3303),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3303),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3298),
.B(n_3136),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3230),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3226),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3177),
.B(n_3136),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3178),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3245),
.Y(n_3411)
);

OAI211xp5_ASAP7_75t_L g3412 ( 
.A1(n_3293),
.A2(n_3039),
.B(n_3061),
.C(n_3049),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3164),
.B(n_3136),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3159),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3300),
.Y(n_3415)
);

OAI21xp33_ASAP7_75t_L g3416 ( 
.A1(n_3254),
.A2(n_2981),
.B(n_3039),
.Y(n_3416)
);

HB1xp67_ASAP7_75t_L g3417 ( 
.A(n_3300),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3300),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3255),
.Y(n_3419)
);

INVx3_ASAP7_75t_L g3420 ( 
.A(n_3188),
.Y(n_3420)
);

OR2x2_ASAP7_75t_L g3421 ( 
.A(n_3227),
.B(n_3091),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3255),
.Y(n_3422)
);

AO21x2_ASAP7_75t_L g3423 ( 
.A1(n_3268),
.A2(n_3005),
.B(n_3049),
.Y(n_3423)
);

AOI222xp33_ASAP7_75t_L g3424 ( 
.A1(n_3254),
.A2(n_3083),
.B1(n_3065),
.B2(n_3090),
.C1(n_3089),
.C2(n_3061),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3157),
.B(n_3005),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_3189),
.A2(n_3101),
.B1(n_3094),
.B2(n_3059),
.Y(n_3426)
);

BUFx2_ASAP7_75t_L g3427 ( 
.A(n_3161),
.Y(n_3427)
);

AOI221xp5_ASAP7_75t_L g3428 ( 
.A1(n_3288),
.A2(n_3071),
.B1(n_3083),
.B2(n_3080),
.C(n_3065),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3183),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3160),
.B(n_3059),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3270),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3234),
.Y(n_3432)
);

AND2x2_ASAP7_75t_L g3433 ( 
.A(n_3184),
.B(n_3147),
.Y(n_3433)
);

BUFx3_ASAP7_75t_L g3434 ( 
.A(n_3152),
.Y(n_3434)
);

BUFx2_ASAP7_75t_L g3435 ( 
.A(n_3263),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3191),
.B(n_3147),
.Y(n_3436)
);

HB1xp67_ASAP7_75t_L g3437 ( 
.A(n_3227),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3276),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3263),
.Y(n_3439)
);

AND2x4_ASAP7_75t_L g3440 ( 
.A(n_3215),
.B(n_3091),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3263),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3276),
.Y(n_3442)
);

INVx3_ASAP7_75t_L g3443 ( 
.A(n_3356),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3411),
.B(n_3154),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_R g3445 ( 
.A(n_3327),
.B(n_3248),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3311),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3311),
.Y(n_3447)
);

OA21x2_ASAP7_75t_L g3448 ( 
.A1(n_3419),
.A2(n_3258),
.B(n_3297),
.Y(n_3448)
);

INVx2_ASAP7_75t_SL g3449 ( 
.A(n_3401),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3356),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3333),
.B(n_3211),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3322),
.A2(n_3247),
.B1(n_3171),
.B2(n_3241),
.Y(n_3452)
);

INVx4_ASAP7_75t_L g3453 ( 
.A(n_3327),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3314),
.Y(n_3454)
);

AO31x2_ASAP7_75t_L g3455 ( 
.A1(n_3366),
.A2(n_3307),
.A3(n_3171),
.B(n_3302),
.Y(n_3455)
);

BUFx2_ASAP7_75t_L g3456 ( 
.A(n_3427),
.Y(n_3456)
);

AOI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_3424),
.A2(n_3307),
.B(n_3244),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3356),
.Y(n_3458)
);

OA21x2_ASAP7_75t_L g3459 ( 
.A1(n_3419),
.A2(n_3258),
.B(n_3154),
.Y(n_3459)
);

BUFx3_ASAP7_75t_L g3460 ( 
.A(n_3427),
.Y(n_3460)
);

NAND2x1_ASAP7_75t_L g3461 ( 
.A(n_3333),
.B(n_3275),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3432),
.B(n_3213),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3432),
.B(n_3205),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3314),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_3326),
.A2(n_3155),
.B1(n_3185),
.B2(n_3241),
.Y(n_3465)
);

INVx2_ASAP7_75t_SL g3466 ( 
.A(n_3401),
.Y(n_3466)
);

INVx2_ASAP7_75t_SL g3467 ( 
.A(n_3321),
.Y(n_3467)
);

OA21x2_ASAP7_75t_L g3468 ( 
.A1(n_3422),
.A2(n_3250),
.B(n_3169),
.Y(n_3468)
);

OR2x2_ASAP7_75t_L g3469 ( 
.A(n_3335),
.B(n_3092),
.Y(n_3469)
);

HB1xp67_ASAP7_75t_L g3470 ( 
.A(n_3316),
.Y(n_3470)
);

AOI21xp33_ASAP7_75t_L g3471 ( 
.A1(n_3396),
.A2(n_3278),
.B(n_3291),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_3341),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3352),
.B(n_3202),
.Y(n_3473)
);

OAI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3343),
.A2(n_3292),
.B(n_3280),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3360),
.Y(n_3475)
);

AO31x2_ASAP7_75t_L g3476 ( 
.A1(n_3366),
.A2(n_3302),
.A3(n_3290),
.B(n_3235),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3360),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3317),
.Y(n_3478)
);

AND2x6_ASAP7_75t_L g3479 ( 
.A(n_3375),
.B(n_3221),
.Y(n_3479)
);

INVx5_ASAP7_75t_L g3480 ( 
.A(n_3376),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3360),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3317),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3361),
.Y(n_3483)
);

BUFx3_ASAP7_75t_L g3484 ( 
.A(n_3341),
.Y(n_3484)
);

INVxp67_ASAP7_75t_SL g3485 ( 
.A(n_3315),
.Y(n_3485)
);

OR2x6_ASAP7_75t_L g3486 ( 
.A(n_3376),
.B(n_3153),
.Y(n_3486)
);

OAI21xp33_ASAP7_75t_L g3487 ( 
.A1(n_3426),
.A2(n_3279),
.B(n_3260),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3361),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3329),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3348),
.B(n_3156),
.Y(n_3490)
);

INVxp67_ASAP7_75t_L g3491 ( 
.A(n_3435),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3329),
.Y(n_3492)
);

OA21x2_ASAP7_75t_L g3493 ( 
.A1(n_3422),
.A2(n_3229),
.B(n_3237),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_L g3494 ( 
.A(n_3420),
.B(n_3275),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3328),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3440),
.B(n_3224),
.Y(n_3496)
);

AO21x2_ASAP7_75t_L g3497 ( 
.A1(n_3414),
.A2(n_3299),
.B(n_3281),
.Y(n_3497)
);

NOR2xp33_ASAP7_75t_L g3498 ( 
.A(n_3420),
.B(n_3402),
.Y(n_3498)
);

AOI22xp33_ASAP7_75t_L g3499 ( 
.A1(n_3322),
.A2(n_3235),
.B1(n_3206),
.B2(n_3253),
.Y(n_3499)
);

OAI221xp5_ASAP7_75t_SL g3500 ( 
.A1(n_3412),
.A2(n_3209),
.B1(n_3228),
.B2(n_3187),
.C(n_3212),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3328),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3344),
.Y(n_3502)
);

AOI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3442),
.A2(n_3290),
.B1(n_3194),
.B2(n_3236),
.Y(n_3503)
);

NOR2x1_ASAP7_75t_L g3504 ( 
.A(n_3420),
.B(n_3194),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3440),
.B(n_3204),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3344),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3348),
.B(n_3259),
.Y(n_3507)
);

BUFx2_ASAP7_75t_L g3508 ( 
.A(n_3435),
.Y(n_3508)
);

OA21x2_ASAP7_75t_L g3509 ( 
.A1(n_3408),
.A2(n_3243),
.B(n_3282),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3351),
.Y(n_3510)
);

NAND2xp33_ASAP7_75t_L g3511 ( 
.A(n_3416),
.B(n_3195),
.Y(n_3511)
);

HB1xp67_ASAP7_75t_L g3512 ( 
.A(n_3354),
.Y(n_3512)
);

INVxp67_ASAP7_75t_L g3513 ( 
.A(n_3398),
.Y(n_3513)
);

AOI22xp5_ASAP7_75t_L g3514 ( 
.A1(n_3438),
.A2(n_3233),
.B1(n_3252),
.B2(n_3240),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3342),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_3342),
.Y(n_3516)
);

AOI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3322),
.A2(n_3294),
.B1(n_3240),
.B2(n_3261),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3363),
.Y(n_3518)
);

INVx3_ASAP7_75t_L g3519 ( 
.A(n_3349),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3363),
.Y(n_3520)
);

A2O1A1Ixp33_ASAP7_75t_L g3521 ( 
.A1(n_3438),
.A2(n_3239),
.B(n_3309),
.C(n_3286),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3351),
.Y(n_3522)
);

BUFx3_ASAP7_75t_L g3523 ( 
.A(n_3434),
.Y(n_3523)
);

OAI21x1_ASAP7_75t_L g3524 ( 
.A1(n_3369),
.A2(n_2992),
.B(n_2986),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3353),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3353),
.Y(n_3526)
);

INVx3_ASAP7_75t_L g3527 ( 
.A(n_3349),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3358),
.Y(n_3528)
);

A2O1A1Ixp33_ASAP7_75t_L g3529 ( 
.A1(n_3378),
.A2(n_3284),
.B(n_3262),
.C(n_3271),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3358),
.Y(n_3530)
);

INVx1_ASAP7_75t_SL g3531 ( 
.A(n_3321),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3434),
.Y(n_3532)
);

O2A1O1Ixp33_ASAP7_75t_L g3533 ( 
.A1(n_3437),
.A2(n_3092),
.B(n_3080),
.C(n_3089),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3384),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3384),
.Y(n_3535)
);

BUFx2_ASAP7_75t_L g3536 ( 
.A(n_3382),
.Y(n_3536)
);

OA21x2_ASAP7_75t_L g3537 ( 
.A1(n_3408),
.A2(n_3082),
.B(n_3122),
.Y(n_3537)
);

AND2x2_ASAP7_75t_L g3538 ( 
.A(n_3382),
.B(n_3395),
.Y(n_3538)
);

AO21x2_ASAP7_75t_L g3539 ( 
.A1(n_3414),
.A2(n_3090),
.B(n_3071),
.Y(n_3539)
);

INVx3_ASAP7_75t_L g3540 ( 
.A(n_3349),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3440),
.B(n_3101),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3347),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3395),
.B(n_3133),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3347),
.Y(n_3544)
);

INVxp67_ASAP7_75t_SL g3545 ( 
.A(n_3439),
.Y(n_3545)
);

AO21x2_ASAP7_75t_L g3546 ( 
.A1(n_3388),
.A2(n_3011),
.B(n_3124),
.Y(n_3546)
);

A2O1A1Ixp33_ASAP7_75t_L g3547 ( 
.A1(n_3365),
.A2(n_3022),
.B(n_3273),
.C(n_3046),
.Y(n_3547)
);

OAI21x1_ASAP7_75t_L g3548 ( 
.A1(n_3369),
.A2(n_3097),
.B(n_3125),
.Y(n_3548)
);

OAI31xp33_ASAP7_75t_L g3549 ( 
.A1(n_3400),
.A2(n_83),
.A3(n_79),
.B(n_80),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3400),
.B(n_3094),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3350),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3362),
.Y(n_3552)
);

OAI21x1_ASAP7_75t_L g3553 ( 
.A1(n_3388),
.A2(n_3108),
.B(n_83),
.Y(n_3553)
);

OR2x2_ASAP7_75t_L g3554 ( 
.A(n_3421),
.B(n_3108),
.Y(n_3554)
);

BUFx3_ASAP7_75t_L g3555 ( 
.A(n_3375),
.Y(n_3555)
);

OAI21x1_ASAP7_75t_L g3556 ( 
.A1(n_3389),
.A2(n_84),
.B(n_85),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3362),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3310),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_L g3559 ( 
.A1(n_3433),
.A2(n_1040),
.B1(n_1036),
.B2(n_88),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_3387),
.B(n_3428),
.Y(n_3560)
);

AO21x2_ASAP7_75t_L g3561 ( 
.A1(n_3389),
.A2(n_3431),
.B(n_3429),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3323),
.B(n_84),
.Y(n_3562)
);

BUFx6f_ASAP7_75t_L g3563 ( 
.A(n_3439),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3325),
.Y(n_3564)
);

A2O1A1Ixp33_ASAP7_75t_L g3565 ( 
.A1(n_3355),
.A2(n_92),
.B(n_87),
.C(n_91),
.Y(n_3565)
);

BUFx2_ASAP7_75t_L g3566 ( 
.A(n_3375),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3334),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_3350),
.Y(n_3568)
);

AOI22xp33_ASAP7_75t_L g3569 ( 
.A1(n_3433),
.A2(n_1040),
.B1(n_95),
.B2(n_91),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3446),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3460),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3460),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3447),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3454),
.Y(n_3574)
);

BUFx2_ASAP7_75t_L g3575 ( 
.A(n_3445),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3464),
.Y(n_3576)
);

AND2x2_ASAP7_75t_L g3577 ( 
.A(n_3538),
.B(n_3393),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_3470),
.Y(n_3578)
);

OR2x2_ASAP7_75t_L g3579 ( 
.A(n_3485),
.B(n_3476),
.Y(n_3579)
);

OR2x2_ASAP7_75t_L g3580 ( 
.A(n_3476),
.B(n_3444),
.Y(n_3580)
);

OR2x2_ASAP7_75t_L g3581 ( 
.A(n_3476),
.B(n_3421),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3538),
.B(n_3393),
.Y(n_3582)
);

OR2x2_ASAP7_75t_L g3583 ( 
.A(n_3476),
.B(n_3463),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3512),
.Y(n_3584)
);

NOR2x1p5_ASAP7_75t_L g3585 ( 
.A(n_3453),
.B(n_3393),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3479),
.B(n_3513),
.Y(n_3586)
);

INVx2_ASAP7_75t_L g3587 ( 
.A(n_3456),
.Y(n_3587)
);

INVx1_ASAP7_75t_SL g3588 ( 
.A(n_3445),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3508),
.Y(n_3589)
);

OAI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3452),
.A2(n_3441),
.B1(n_3336),
.B2(n_3385),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3536),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3478),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3482),
.Y(n_3593)
);

NAND3xp33_ASAP7_75t_L g3594 ( 
.A(n_3471),
.B(n_3418),
.C(n_3415),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3480),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3486),
.B(n_3320),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3486),
.B(n_3441),
.Y(n_3597)
);

INVx4_ASAP7_75t_L g3598 ( 
.A(n_3453),
.Y(n_3598)
);

AND2x2_ASAP7_75t_L g3599 ( 
.A(n_3486),
.B(n_3339),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3480),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3495),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3501),
.Y(n_3602)
);

OR2x2_ASAP7_75t_L g3603 ( 
.A(n_3496),
.B(n_3335),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3480),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3502),
.Y(n_3605)
);

BUFx2_ASAP7_75t_L g3606 ( 
.A(n_3486),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3479),
.B(n_3404),
.Y(n_3607)
);

INVxp33_ASAP7_75t_SL g3608 ( 
.A(n_3498),
.Y(n_3608)
);

OR2x2_ASAP7_75t_L g3609 ( 
.A(n_3462),
.B(n_3368),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3506),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3449),
.B(n_3320),
.Y(n_3611)
);

INVx4_ASAP7_75t_L g3612 ( 
.A(n_3453),
.Y(n_3612)
);

BUFx3_ASAP7_75t_L g3613 ( 
.A(n_3472),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3510),
.Y(n_3614)
);

AND2x4_ASAP7_75t_L g3615 ( 
.A(n_3480),
.B(n_3346),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_3449),
.B(n_3409),
.Y(n_3616)
);

NAND3xp33_ASAP7_75t_L g3617 ( 
.A(n_3499),
.B(n_3418),
.C(n_3415),
.Y(n_3617)
);

AO21x2_ASAP7_75t_L g3618 ( 
.A1(n_3562),
.A2(n_3319),
.B(n_3312),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3522),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_3531),
.B(n_3490),
.Y(n_3620)
);

AND2x2_ASAP7_75t_L g3621 ( 
.A(n_3490),
.B(n_3339),
.Y(n_3621)
);

INVxp67_ASAP7_75t_L g3622 ( 
.A(n_3479),
.Y(n_3622)
);

AOI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_3511),
.A2(n_3425),
.B1(n_3430),
.B2(n_3423),
.Y(n_3623)
);

AO31x2_ASAP7_75t_L g3624 ( 
.A1(n_3566),
.A2(n_3431),
.A3(n_3313),
.B(n_3318),
.Y(n_3624)
);

AOI22xp5_ASAP7_75t_L g3625 ( 
.A1(n_3487),
.A2(n_3436),
.B1(n_3425),
.B2(n_3409),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3525),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3479),
.B(n_3404),
.Y(n_3627)
);

BUFx2_ASAP7_75t_L g3628 ( 
.A(n_3555),
.Y(n_3628)
);

AND2x2_ASAP7_75t_L g3629 ( 
.A(n_3466),
.B(n_3336),
.Y(n_3629)
);

HB1xp67_ASAP7_75t_L g3630 ( 
.A(n_3483),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3466),
.B(n_3397),
.Y(n_3631)
);

BUFx2_ASAP7_75t_L g3632 ( 
.A(n_3555),
.Y(n_3632)
);

INVxp67_ASAP7_75t_SL g3633 ( 
.A(n_3468),
.Y(n_3633)
);

NOR2xp33_ASAP7_75t_L g3634 ( 
.A(n_3498),
.B(n_3405),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3526),
.Y(n_3635)
);

AOI22xp33_ASAP7_75t_L g3636 ( 
.A1(n_3511),
.A2(n_3430),
.B1(n_3423),
.B2(n_3436),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3467),
.B(n_3484),
.Y(n_3637)
);

AND2x4_ASAP7_75t_SL g3638 ( 
.A(n_3472),
.B(n_3405),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3480),
.B(n_3313),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_L g3640 ( 
.A(n_3560),
.B(n_3345),
.Y(n_3640)
);

OAI33xp33_ASAP7_75t_L g3641 ( 
.A1(n_3465),
.A2(n_3391),
.A3(n_3394),
.B1(n_3380),
.B2(n_3331),
.B3(n_3338),
.Y(n_3641)
);

OR2x2_ASAP7_75t_L g3642 ( 
.A(n_3469),
.B(n_3368),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3528),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3479),
.B(n_3457),
.Y(n_3644)
);

BUFx3_ASAP7_75t_L g3645 ( 
.A(n_3472),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3467),
.B(n_3318),
.Y(n_3646)
);

NAND2x1_ASAP7_75t_SL g3647 ( 
.A(n_3504),
.B(n_3346),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3451),
.B(n_3392),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3484),
.B(n_3397),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3530),
.Y(n_3650)
);

OR2x2_ASAP7_75t_L g3651 ( 
.A(n_3505),
.B(n_3338),
.Y(n_3651)
);

NAND3xp33_ASAP7_75t_L g3652 ( 
.A(n_3474),
.B(n_3417),
.C(n_3429),
.Y(n_3652)
);

HB1xp67_ASAP7_75t_L g3653 ( 
.A(n_3483),
.Y(n_3653)
);

INVxp67_ASAP7_75t_L g3654 ( 
.A(n_3479),
.Y(n_3654)
);

AOI33xp33_ASAP7_75t_L g3655 ( 
.A1(n_3517),
.A2(n_3406),
.A3(n_3413),
.B1(n_3379),
.B2(n_3312),
.B3(n_3319),
.Y(n_3655)
);

AOI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_3497),
.A2(n_3423),
.B1(n_3406),
.B2(n_3407),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3451),
.B(n_3392),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3552),
.Y(n_3658)
);

OR2x2_ASAP7_75t_L g3659 ( 
.A(n_3473),
.B(n_3379),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3563),
.Y(n_3660)
);

INVxp67_ASAP7_75t_SL g3661 ( 
.A(n_3468),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3557),
.Y(n_3662)
);

BUFx2_ASAP7_75t_L g3663 ( 
.A(n_3523),
.Y(n_3663)
);

OAI211xp5_ASAP7_75t_L g3664 ( 
.A1(n_3549),
.A2(n_3413),
.B(n_3331),
.C(n_3390),
.Y(n_3664)
);

AND2x4_ASAP7_75t_L g3665 ( 
.A(n_3491),
.B(n_3346),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3563),
.Y(n_3666)
);

AOI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3521),
.A2(n_3332),
.B(n_3403),
.Y(n_3667)
);

AOI22xp33_ASAP7_75t_L g3668 ( 
.A1(n_3497),
.A2(n_3330),
.B1(n_3324),
.B2(n_3410),
.Y(n_3668)
);

AND2x2_ASAP7_75t_L g3669 ( 
.A(n_3523),
.B(n_3383),
.Y(n_3669)
);

OR2x2_ASAP7_75t_L g3670 ( 
.A(n_3534),
.B(n_3377),
.Y(n_3670)
);

INVx1_ASAP7_75t_SL g3671 ( 
.A(n_3532),
.Y(n_3671)
);

INVx4_ASAP7_75t_L g3672 ( 
.A(n_3472),
.Y(n_3672)
);

OAI321xp33_ASAP7_75t_L g3673 ( 
.A1(n_3500),
.A2(n_3324),
.A3(n_3330),
.B1(n_3399),
.B2(n_3340),
.C(n_3357),
.Y(n_3673)
);

OR2x2_ASAP7_75t_L g3674 ( 
.A(n_3534),
.B(n_3337),
.Y(n_3674)
);

OR2x2_ASAP7_75t_L g3675 ( 
.A(n_3535),
.B(n_3337),
.Y(n_3675)
);

BUFx2_ASAP7_75t_L g3676 ( 
.A(n_3532),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3563),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3558),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3543),
.B(n_3383),
.Y(n_3679)
);

OR2x2_ASAP7_75t_L g3680 ( 
.A(n_3535),
.B(n_3367),
.Y(n_3680)
);

NAND4xp25_ASAP7_75t_L g3681 ( 
.A(n_3521),
.B(n_3359),
.C(n_3357),
.D(n_3386),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3494),
.B(n_3364),
.Y(n_3682)
);

INVx2_ASAP7_75t_SL g3683 ( 
.A(n_3563),
.Y(n_3683)
);

AND2x4_ASAP7_75t_SL g3684 ( 
.A(n_3494),
.B(n_3364),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3584),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3584),
.Y(n_3686)
);

OR2x2_ASAP7_75t_L g3687 ( 
.A(n_3603),
.B(n_3455),
.Y(n_3687)
);

OR2x2_ASAP7_75t_L g3688 ( 
.A(n_3609),
.B(n_3455),
.Y(n_3688)
);

AND2x2_ASAP7_75t_L g3689 ( 
.A(n_3620),
.B(n_3461),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_SL g3690 ( 
.A1(n_3644),
.A2(n_3565),
.B(n_3459),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3578),
.Y(n_3691)
);

AND2x2_ASAP7_75t_L g3692 ( 
.A(n_3577),
.B(n_3545),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3613),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3582),
.B(n_3507),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3578),
.Y(n_3695)
);

OR2x2_ASAP7_75t_L g3696 ( 
.A(n_3617),
.B(n_3455),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3630),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3630),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_SL g3699 ( 
.A(n_3673),
.B(n_3503),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3671),
.B(n_3455),
.Y(n_3700)
);

INVxp67_ASAP7_75t_SL g3701 ( 
.A(n_3647),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3587),
.B(n_3497),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3587),
.B(n_3514),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3653),
.Y(n_3704)
);

INVx5_ASAP7_75t_L g3705 ( 
.A(n_3598),
.Y(n_3705)
);

AND2x2_ASAP7_75t_L g3706 ( 
.A(n_3637),
.B(n_3507),
.Y(n_3706)
);

BUFx2_ASAP7_75t_SL g3707 ( 
.A(n_3613),
.Y(n_3707)
);

BUFx3_ASAP7_75t_L g3708 ( 
.A(n_3575),
.Y(n_3708)
);

OR2x2_ASAP7_75t_L g3709 ( 
.A(n_3659),
.B(n_3651),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3645),
.Y(n_3710)
);

INVx4_ASAP7_75t_L g3711 ( 
.A(n_3598),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3621),
.B(n_3543),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3645),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3663),
.Y(n_3714)
);

OR2x2_ASAP7_75t_L g3715 ( 
.A(n_3680),
.B(n_3459),
.Y(n_3715)
);

OAI22xp5_ASAP7_75t_L g3716 ( 
.A1(n_3668),
.A2(n_3529),
.B1(n_3569),
.B2(n_3559),
.Y(n_3716)
);

AND2x2_ASAP7_75t_L g3717 ( 
.A(n_3676),
.B(n_3629),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3588),
.B(n_3459),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3638),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3591),
.B(n_3468),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3638),
.B(n_3550),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3599),
.B(n_3550),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3591),
.B(n_3564),
.Y(n_3723)
);

OR2x2_ASAP7_75t_L g3724 ( 
.A(n_3607),
.B(n_3567),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3571),
.B(n_3533),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3669),
.B(n_3381),
.Y(n_3726)
);

AND2x4_ASAP7_75t_L g3727 ( 
.A(n_3585),
.B(n_3519),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3653),
.Y(n_3728)
);

HB1xp67_ASAP7_75t_L g3729 ( 
.A(n_3589),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3672),
.Y(n_3730)
);

OAI22xp5_ASAP7_75t_L g3731 ( 
.A1(n_3668),
.A2(n_3529),
.B1(n_3547),
.B2(n_3565),
.Y(n_3731)
);

OR2x2_ASAP7_75t_L g3732 ( 
.A(n_3627),
.B(n_3493),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3606),
.B(n_3450),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3608),
.B(n_3541),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3628),
.B(n_3450),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3632),
.B(n_3458),
.Y(n_3736)
);

NOR2xp33_ASAP7_75t_L g3737 ( 
.A(n_3608),
.B(n_3489),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3571),
.B(n_3493),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3570),
.Y(n_3739)
);

AND2x2_ASAP7_75t_L g3740 ( 
.A(n_3596),
.B(n_3458),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3573),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3596),
.B(n_3475),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3580),
.B(n_3493),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3597),
.B(n_3475),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3574),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3572),
.B(n_3556),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3572),
.B(n_3556),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3611),
.B(n_3477),
.Y(n_3748)
);

AND2x2_ASAP7_75t_L g3749 ( 
.A(n_3611),
.B(n_3477),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3576),
.Y(n_3750)
);

HB1xp67_ASAP7_75t_L g3751 ( 
.A(n_3589),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_SL g3752 ( 
.A(n_3656),
.B(n_3633),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3684),
.B(n_3481),
.Y(n_3753)
);

INVxp67_ASAP7_75t_SL g3754 ( 
.A(n_3633),
.Y(n_3754)
);

OR2x2_ASAP7_75t_L g3755 ( 
.A(n_3583),
.B(n_3489),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3672),
.Y(n_3756)
);

OR2x2_ASAP7_75t_L g3757 ( 
.A(n_3674),
.B(n_3492),
.Y(n_3757)
);

HB1xp67_ASAP7_75t_L g3758 ( 
.A(n_3595),
.Y(n_3758)
);

OR2x2_ASAP7_75t_L g3759 ( 
.A(n_3675),
.B(n_3492),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3672),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3592),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3593),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_3594),
.B(n_3579),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3634),
.B(n_3515),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_SL g3765 ( 
.A(n_3656),
.B(n_3661),
.Y(n_3765)
);

NAND2xp5_ASAP7_75t_L g3766 ( 
.A(n_3634),
.B(n_3515),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3601),
.Y(n_3767)
);

INVx4_ASAP7_75t_L g3768 ( 
.A(n_3598),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3612),
.B(n_3516),
.Y(n_3769)
);

INVx1_ASAP7_75t_SL g3770 ( 
.A(n_3684),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3648),
.B(n_3481),
.Y(n_3771)
);

AND3x2_ASAP7_75t_L g3772 ( 
.A(n_3661),
.B(n_3516),
.C(n_3488),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3602),
.Y(n_3773)
);

INVx2_ASAP7_75t_SL g3774 ( 
.A(n_3615),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3648),
.B(n_3519),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3657),
.B(n_3519),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3754),
.Y(n_3777)
);

NAND4xp75_ASAP7_75t_SL g3778 ( 
.A(n_3734),
.B(n_3616),
.C(n_3640),
.D(n_3639),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3729),
.Y(n_3779)
);

XOR2x2_ASAP7_75t_L g3780 ( 
.A(n_3699),
.B(n_3586),
.Y(n_3780)
);

NAND4xp75_ASAP7_75t_SL g3781 ( 
.A(n_3734),
.B(n_3616),
.C(n_3640),
.D(n_3639),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3717),
.B(n_3682),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3751),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3772),
.Y(n_3784)
);

NAND4xp75_ASAP7_75t_L g3785 ( 
.A(n_3752),
.B(n_3625),
.C(n_3600),
.D(n_3604),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3708),
.Y(n_3786)
);

INVx4_ASAP7_75t_L g3787 ( 
.A(n_3705),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3708),
.Y(n_3788)
);

BUFx2_ASAP7_75t_L g3789 ( 
.A(n_3774),
.Y(n_3789)
);

INVx1_ASAP7_75t_SL g3790 ( 
.A(n_3707),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3705),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3758),
.Y(n_3792)
);

BUFx2_ASAP7_75t_L g3793 ( 
.A(n_3774),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3685),
.Y(n_3794)
);

INVx2_ASAP7_75t_SL g3795 ( 
.A(n_3705),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3705),
.Y(n_3796)
);

BUFx2_ASAP7_75t_L g3797 ( 
.A(n_3714),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3705),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3717),
.B(n_3689),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3706),
.B(n_3657),
.Y(n_3800)
);

INVxp67_ASAP7_75t_L g3801 ( 
.A(n_3718),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3686),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3706),
.B(n_3649),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3691),
.Y(n_3804)
);

INVx2_ASAP7_75t_SL g3805 ( 
.A(n_3775),
.Y(n_3805)
);

BUFx3_ASAP7_75t_L g3806 ( 
.A(n_3714),
.Y(n_3806)
);

OR2x2_ASAP7_75t_L g3807 ( 
.A(n_3709),
.B(n_3622),
.Y(n_3807)
);

XNOR2xp5_ASAP7_75t_L g3808 ( 
.A(n_3699),
.B(n_3681),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3693),
.B(n_3654),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3693),
.B(n_3612),
.Y(n_3810)
);

AND2x4_ASAP7_75t_L g3811 ( 
.A(n_3719),
.B(n_3711),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3721),
.Y(n_3812)
);

XOR2x2_ASAP7_75t_L g3813 ( 
.A(n_3731),
.B(n_3590),
.Y(n_3813)
);

XNOR2xp5_ASAP7_75t_L g3814 ( 
.A(n_3716),
.B(n_3664),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3721),
.B(n_3646),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3695),
.Y(n_3816)
);

NAND4xp75_ASAP7_75t_L g3817 ( 
.A(n_3752),
.B(n_3595),
.C(n_3604),
.D(n_3600),
.Y(n_3817)
);

NAND4xp75_ASAP7_75t_L g3818 ( 
.A(n_3765),
.B(n_3683),
.C(n_3667),
.D(n_3666),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3710),
.B(n_3612),
.Y(n_3819)
);

XOR2x2_ASAP7_75t_L g3820 ( 
.A(n_3765),
.B(n_3652),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3697),
.Y(n_3821)
);

HB1xp67_ASAP7_75t_L g3822 ( 
.A(n_3698),
.Y(n_3822)
);

NAND4xp75_ASAP7_75t_SL g3823 ( 
.A(n_3718),
.B(n_3646),
.C(n_3631),
.D(n_3679),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_3704),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3728),
.Y(n_3825)
);

INVx4_ASAP7_75t_L g3826 ( 
.A(n_3711),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3755),
.Y(n_3827)
);

XOR2x2_ASAP7_75t_L g3828 ( 
.A(n_3696),
.B(n_3623),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3710),
.B(n_3713),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3775),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3739),
.Y(n_3831)
);

NAND4xp75_ASAP7_75t_L g3832 ( 
.A(n_3702),
.B(n_3683),
.C(n_3660),
.D(n_3677),
.Y(n_3832)
);

INVx1_ASAP7_75t_SL g3833 ( 
.A(n_3692),
.Y(n_3833)
);

INVx2_ASAP7_75t_SL g3834 ( 
.A(n_3776),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_3694),
.B(n_3665),
.Y(n_3835)
);

OAI21xp33_ASAP7_75t_L g3836 ( 
.A1(n_3690),
.A2(n_3655),
.B(n_3636),
.Y(n_3836)
);

XNOR2xp5_ASAP7_75t_L g3837 ( 
.A(n_3770),
.B(n_3636),
.Y(n_3837)
);

NAND4xp75_ASAP7_75t_L g3838 ( 
.A(n_3720),
.B(n_3666),
.C(n_3677),
.D(n_3660),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3741),
.Y(n_3839)
);

NOR2x1_ASAP7_75t_L g3840 ( 
.A(n_3711),
.B(n_3581),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3694),
.B(n_3665),
.Y(n_3841)
);

NAND4xp75_ASAP7_75t_L g3842 ( 
.A(n_3700),
.B(n_3641),
.C(n_3623),
.D(n_3678),
.Y(n_3842)
);

NOR4xp25_ASAP7_75t_L g3843 ( 
.A(n_3763),
.B(n_3655),
.C(n_3547),
.D(n_3610),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3776),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3768),
.Y(n_3845)
);

AND2x4_ASAP7_75t_L g3846 ( 
.A(n_3719),
.B(n_3615),
.Y(n_3846)
);

AND2x4_ASAP7_75t_L g3847 ( 
.A(n_3768),
.B(n_3615),
.Y(n_3847)
);

AOI22xp5_ASAP7_75t_L g3848 ( 
.A1(n_3701),
.A2(n_3665),
.B1(n_3618),
.B2(n_3679),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3745),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3692),
.B(n_3712),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3750),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3712),
.B(n_3618),
.Y(n_3852)
);

AOI22xp33_ASAP7_75t_L g3853 ( 
.A1(n_3703),
.A2(n_3448),
.B1(n_3509),
.B2(n_3605),
.Y(n_3853)
);

NOR4xp25_ASAP7_75t_L g3854 ( 
.A(n_3713),
.B(n_3614),
.C(n_3626),
.D(n_3619),
.Y(n_3854)
);

XOR2xp5_ASAP7_75t_L g3855 ( 
.A(n_3688),
.B(n_3670),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3768),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3722),
.B(n_3735),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3730),
.Y(n_3858)
);

XNOR2xp5_ASAP7_75t_L g3859 ( 
.A(n_3722),
.B(n_3635),
.Y(n_3859)
);

INVx2_ASAP7_75t_SL g3860 ( 
.A(n_3727),
.Y(n_3860)
);

INVx1_ASAP7_75t_SL g3861 ( 
.A(n_3735),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3761),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3737),
.B(n_3643),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3762),
.Y(n_3864)
);

AND2x2_ASAP7_75t_L g3865 ( 
.A(n_3736),
.B(n_3527),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3730),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3756),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3767),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3822),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3861),
.B(n_3737),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_3833),
.B(n_3756),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_3799),
.B(n_3753),
.Y(n_3872)
);

OAI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3818),
.A2(n_3743),
.B(n_3725),
.Y(n_3873)
);

OR2x2_ASAP7_75t_L g3874 ( 
.A(n_3786),
.B(n_3687),
.Y(n_3874)
);

NOR2xp67_ASAP7_75t_L g3875 ( 
.A(n_3787),
.B(n_3727),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3806),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3828),
.B(n_3760),
.Y(n_3877)
);

AOI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_3836),
.A2(n_3738),
.B1(n_3732),
.B2(n_3746),
.Y(n_3878)
);

AND2x4_ASAP7_75t_L g3879 ( 
.A(n_3806),
.B(n_3760),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3828),
.B(n_3773),
.Y(n_3880)
);

NAND2x1p5_ASAP7_75t_L g3881 ( 
.A(n_3790),
.B(n_3727),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3820),
.B(n_3723),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3820),
.B(n_3843),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3822),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3799),
.B(n_3753),
.Y(n_3885)
);

AOI22xp33_ASAP7_75t_SL g3886 ( 
.A1(n_3784),
.A2(n_3715),
.B1(n_3736),
.B2(n_3771),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3797),
.Y(n_3887)
);

NAND3xp33_ASAP7_75t_L g3888 ( 
.A(n_3801),
.B(n_3769),
.C(n_3747),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3789),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3857),
.B(n_3726),
.Y(n_3890)
);

OAI22xp33_ASAP7_75t_L g3891 ( 
.A1(n_3784),
.A2(n_3766),
.B1(n_3764),
.B2(n_3724),
.Y(n_3891)
);

NAND2x1p5_ASAP7_75t_L g3892 ( 
.A(n_3787),
.B(n_3733),
.Y(n_3892)
);

OR2x2_ASAP7_75t_L g3893 ( 
.A(n_3786),
.B(n_3757),
.Y(n_3893)
);

INVx1_ASAP7_75t_SL g3894 ( 
.A(n_3793),
.Y(n_3894)
);

INVx1_ASAP7_75t_SL g3895 ( 
.A(n_3817),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3792),
.Y(n_3896)
);

AND2x2_ASAP7_75t_L g3897 ( 
.A(n_3857),
.B(n_3744),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3860),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3850),
.B(n_3800),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3830),
.Y(n_3900)
);

OR2x2_ASAP7_75t_L g3901 ( 
.A(n_3788),
.B(n_3759),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3850),
.B(n_3744),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3830),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3844),
.Y(n_3904)
);

OR2x2_ASAP7_75t_L g3905 ( 
.A(n_3788),
.B(n_3829),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3844),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3860),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3800),
.B(n_3771),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3782),
.B(n_3733),
.Y(n_3909)
);

OR2x2_ASAP7_75t_L g3910 ( 
.A(n_3807),
.B(n_3809),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3858),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3812),
.B(n_3769),
.Y(n_3912)
);

INVxp67_ASAP7_75t_SL g3913 ( 
.A(n_3840),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3858),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3842),
.B(n_3650),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3808),
.B(n_3658),
.Y(n_3916)
);

INVxp67_ASAP7_75t_L g3917 ( 
.A(n_3815),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3866),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3812),
.B(n_3740),
.Y(n_3919)
);

INVxp67_ASAP7_75t_SL g3920 ( 
.A(n_3815),
.Y(n_3920)
);

NAND2x1p5_ASAP7_75t_L g3921 ( 
.A(n_3787),
.B(n_3740),
.Y(n_3921)
);

INVxp67_ASAP7_75t_L g3922 ( 
.A(n_3835),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_L g3923 ( 
.A(n_3810),
.B(n_3742),
.Y(n_3923)
);

OR2x2_ASAP7_75t_L g3924 ( 
.A(n_3805),
.B(n_3642),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3866),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3867),
.Y(n_3926)
);

NAND2x2_ASAP7_75t_L g3927 ( 
.A(n_3805),
.B(n_3554),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3835),
.B(n_3742),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3867),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3779),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3841),
.B(n_3748),
.Y(n_3931)
);

AOI32xp33_ASAP7_75t_L g3932 ( 
.A1(n_3841),
.A2(n_3749),
.A3(n_3748),
.B1(n_3662),
.B2(n_3540),
.Y(n_3932)
);

AND2x2_ASAP7_75t_L g3933 ( 
.A(n_3803),
.B(n_3749),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3846),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3783),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3777),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3834),
.Y(n_3937)
);

NAND3xp33_ASAP7_75t_L g3938 ( 
.A(n_3814),
.B(n_3448),
.C(n_3554),
.Y(n_3938)
);

OR2x2_ASAP7_75t_L g3939 ( 
.A(n_3834),
.B(n_3542),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3803),
.B(n_3488),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3854),
.B(n_3518),
.Y(n_3941)
);

OR2x2_ASAP7_75t_L g3942 ( 
.A(n_3863),
.B(n_3542),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3846),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3846),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3865),
.B(n_3518),
.Y(n_3945)
);

OR2x2_ASAP7_75t_L g3946 ( 
.A(n_3827),
.B(n_3544),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3865),
.B(n_3520),
.Y(n_3947)
);

INVx2_ASAP7_75t_SL g3948 ( 
.A(n_3847),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3794),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3811),
.B(n_3520),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3811),
.B(n_3837),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3802),
.Y(n_3952)
);

OR2x6_ASAP7_75t_L g3953 ( 
.A(n_3826),
.B(n_3553),
.Y(n_3953)
);

INVxp67_ASAP7_75t_L g3954 ( 
.A(n_3838),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3804),
.Y(n_3955)
);

NAND2x1p5_ASAP7_75t_L g3956 ( 
.A(n_3847),
.B(n_3553),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3816),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3821),
.Y(n_3958)
);

OAI22xp5_ASAP7_75t_L g3959 ( 
.A1(n_3883),
.A2(n_3785),
.B1(n_3853),
.B2(n_3855),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3894),
.B(n_3811),
.Y(n_3960)
);

OAI21xp33_ASAP7_75t_L g3961 ( 
.A1(n_3883),
.A2(n_3813),
.B(n_3780),
.Y(n_3961)
);

AOI22xp5_ASAP7_75t_L g3962 ( 
.A1(n_3895),
.A2(n_3813),
.B1(n_3780),
.B2(n_3832),
.Y(n_3962)
);

NAND3xp33_ASAP7_75t_L g3963 ( 
.A(n_3873),
.B(n_3853),
.C(n_3848),
.Y(n_3963)
);

INVx2_ASAP7_75t_SL g3964 ( 
.A(n_3879),
.Y(n_3964)
);

AOI221xp5_ASAP7_75t_L g3965 ( 
.A1(n_3895),
.A2(n_3824),
.B1(n_3825),
.B2(n_3859),
.C(n_3819),
.Y(n_3965)
);

OAI31xp33_ASAP7_75t_L g3966 ( 
.A1(n_3938),
.A2(n_3852),
.A3(n_3781),
.B(n_3778),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3920),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3869),
.Y(n_3968)
);

AOI211x1_ASAP7_75t_L g3969 ( 
.A1(n_3873),
.A2(n_3852),
.B(n_3831),
.C(n_3849),
.Y(n_3969)
);

NOR2xp33_ASAP7_75t_L g3970 ( 
.A(n_3881),
.B(n_3826),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3884),
.Y(n_3971)
);

OAI22xp5_ASAP7_75t_L g3972 ( 
.A1(n_3882),
.A2(n_3795),
.B1(n_3847),
.B2(n_3845),
.Y(n_3972)
);

AOI22xp5_ASAP7_75t_L g3973 ( 
.A1(n_3954),
.A2(n_3795),
.B1(n_3851),
.B2(n_3839),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3899),
.Y(n_3974)
);

AOI22xp5_ASAP7_75t_L g3975 ( 
.A1(n_3882),
.A2(n_3856),
.B1(n_3845),
.B2(n_3796),
.Y(n_3975)
);

AOI22xp5_ASAP7_75t_L g3976 ( 
.A1(n_3880),
.A2(n_3862),
.B1(n_3868),
.B2(n_3864),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3934),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3892),
.Y(n_3978)
);

OAI211xp5_ASAP7_75t_L g3979 ( 
.A1(n_3878),
.A2(n_3826),
.B(n_3856),
.C(n_3796),
.Y(n_3979)
);

AO21x1_ASAP7_75t_L g3980 ( 
.A1(n_3913),
.A2(n_3798),
.B(n_3791),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3943),
.Y(n_3981)
);

OR2x2_ASAP7_75t_L g3982 ( 
.A(n_3894),
.B(n_3877),
.Y(n_3982)
);

OAI22xp33_ASAP7_75t_SL g3983 ( 
.A1(n_3927),
.A2(n_3798),
.B1(n_3791),
.B2(n_3823),
.Y(n_3983)
);

NOR2xp33_ASAP7_75t_SL g3984 ( 
.A(n_3872),
.B(n_3544),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3944),
.Y(n_3985)
);

A2O1A1Ixp33_ASAP7_75t_L g3986 ( 
.A1(n_3938),
.A2(n_3548),
.B(n_3524),
.C(n_3540),
.Y(n_3986)
);

AOI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3880),
.A2(n_3448),
.B1(n_3509),
.B2(n_3561),
.Y(n_3987)
);

AOI32xp33_ASAP7_75t_L g3988 ( 
.A1(n_3915),
.A2(n_3540),
.A3(n_3527),
.B1(n_3443),
.B2(n_3551),
.Y(n_3988)
);

NOR2xp33_ASAP7_75t_L g3989 ( 
.A(n_3951),
.B(n_3910),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3937),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_3879),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3921),
.Y(n_3992)
);

OAI221xp5_ASAP7_75t_L g3993 ( 
.A1(n_3878),
.A2(n_3527),
.B1(n_3568),
.B2(n_3551),
.C(n_3443),
.Y(n_3993)
);

AOI211xp5_ASAP7_75t_L g3994 ( 
.A1(n_3915),
.A2(n_3548),
.B(n_3568),
.C(n_3524),
.Y(n_3994)
);

OAI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3888),
.A2(n_3509),
.B(n_3443),
.Y(n_3995)
);

OR2x2_ASAP7_75t_L g3996 ( 
.A(n_3877),
.B(n_3624),
.Y(n_3996)
);

OAI22xp33_ASAP7_75t_SL g3997 ( 
.A1(n_3941),
.A2(n_3624),
.B1(n_3374),
.B2(n_3372),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3908),
.Y(n_3998)
);

AND2x4_ASAP7_75t_L g3999 ( 
.A(n_3875),
.B(n_3624),
.Y(n_3999)
);

AOI211xp5_ASAP7_75t_SL g4000 ( 
.A1(n_3891),
.A2(n_3359),
.B(n_3386),
.C(n_3624),
.Y(n_4000)
);

AOI21xp33_ASAP7_75t_SL g4001 ( 
.A1(n_3870),
.A2(n_3561),
.B(n_93),
.Y(n_4001)
);

NAND3xp33_ASAP7_75t_L g4002 ( 
.A(n_3886),
.B(n_3537),
.C(n_3371),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3887),
.Y(n_4003)
);

XNOR2xp5_ASAP7_75t_L g4004 ( 
.A(n_3928),
.B(n_93),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3948),
.Y(n_4005)
);

OAI21xp5_ASAP7_75t_SL g4006 ( 
.A1(n_3922),
.A2(n_3370),
.B(n_3381),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3900),
.Y(n_4007)
);

OAI31xp33_ASAP7_75t_L g4008 ( 
.A1(n_3941),
.A2(n_3539),
.A3(n_3373),
.B(n_3561),
.Y(n_4008)
);

NAND4xp75_ASAP7_75t_L g4009 ( 
.A(n_3875),
.B(n_3537),
.C(n_3373),
.D(n_98),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3916),
.A2(n_3537),
.B1(n_3539),
.B2(n_3546),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3885),
.B(n_3902),
.Y(n_4011)
);

XNOR2xp5_ASAP7_75t_L g4012 ( 
.A(n_3931),
.B(n_96),
.Y(n_4012)
);

OAI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_3888),
.A2(n_3539),
.B(n_3546),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3903),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_L g4015 ( 
.A(n_3923),
.B(n_3909),
.Y(n_4015)
);

OAI31xp33_ASAP7_75t_L g4016 ( 
.A1(n_3956),
.A2(n_3546),
.A3(n_99),
.B(n_97),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3904),
.Y(n_4017)
);

OAI21xp5_ASAP7_75t_L g4018 ( 
.A1(n_3917),
.A2(n_98),
.B(n_100),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3897),
.B(n_101),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3906),
.Y(n_4020)
);

OAI21xp33_ASAP7_75t_L g4021 ( 
.A1(n_3933),
.A2(n_101),
.B(n_102),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3898),
.Y(n_4022)
);

AOI21xp33_ASAP7_75t_L g4023 ( 
.A1(n_3893),
.A2(n_102),
.B(n_103),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3907),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3911),
.Y(n_4025)
);

BUFx2_ASAP7_75t_SL g4026 ( 
.A(n_3876),
.Y(n_4026)
);

OAI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3953),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3890),
.B(n_106),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3889),
.Y(n_4029)
);

INVxp67_ASAP7_75t_L g4030 ( 
.A(n_3924),
.Y(n_4030)
);

OAI21xp33_ASAP7_75t_L g4031 ( 
.A1(n_3916),
.A2(n_107),
.B(n_108),
.Y(n_4031)
);

INVxp67_ASAP7_75t_L g4032 ( 
.A(n_3919),
.Y(n_4032)
);

AOI22xp33_ASAP7_75t_L g4033 ( 
.A1(n_3936),
.A2(n_112),
.B1(n_108),
.B2(n_109),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3950),
.B(n_109),
.Y(n_4034)
);

CKINVDCx14_ASAP7_75t_R g4035 ( 
.A(n_3905),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3914),
.Y(n_4036)
);

INVx1_ASAP7_75t_SL g4037 ( 
.A(n_3901),
.Y(n_4037)
);

AOI21xp33_ASAP7_75t_L g4038 ( 
.A1(n_3871),
.A2(n_112),
.B(n_113),
.Y(n_4038)
);

OAI22xp33_ASAP7_75t_SL g4039 ( 
.A1(n_3874),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_4039)
);

INVx1_ASAP7_75t_SL g4040 ( 
.A(n_3939),
.Y(n_4040)
);

OAI22xp5_ASAP7_75t_L g4041 ( 
.A1(n_3912),
.A2(n_117),
.B1(n_114),
.B2(n_115),
.Y(n_4041)
);

OAI22xp33_ASAP7_75t_L g4042 ( 
.A1(n_3953),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3960),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_4011),
.B(n_3896),
.Y(n_4044)
);

OAI21xp33_ASAP7_75t_L g4045 ( 
.A1(n_3961),
.A2(n_3932),
.B(n_3930),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_4005),
.B(n_3935),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3964),
.B(n_3918),
.Y(n_4047)
);

AOI22xp5_ASAP7_75t_L g4048 ( 
.A1(n_3959),
.A2(n_3940),
.B1(n_3947),
.B2(n_3945),
.Y(n_4048)
);

OR2x2_ASAP7_75t_L g4049 ( 
.A(n_3982),
.B(n_3946),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3991),
.Y(n_4050)
);

OAI21xp5_ASAP7_75t_SL g4051 ( 
.A1(n_3962),
.A2(n_3952),
.B(n_3949),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3974),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3980),
.Y(n_4053)
);

OR2x2_ASAP7_75t_L g4054 ( 
.A(n_4037),
.B(n_3942),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3962),
.B(n_3925),
.Y(n_4055)
);

INVx2_ASAP7_75t_SL g4056 ( 
.A(n_3978),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3998),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_4035),
.B(n_3955),
.Y(n_4058)
);

O2A1O1Ixp33_ASAP7_75t_L g4059 ( 
.A1(n_3963),
.A2(n_3958),
.B(n_3957),
.C(n_3929),
.Y(n_4059)
);

OAI21xp33_ASAP7_75t_L g4060 ( 
.A1(n_3989),
.A2(n_3984),
.B(n_4015),
.Y(n_4060)
);

OAI211xp5_ASAP7_75t_SL g4061 ( 
.A1(n_3966),
.A2(n_3926),
.B(n_3953),
.C(n_121),
.Y(n_4061)
);

OAI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3969),
.A2(n_123),
.B1(n_118),
.B2(n_119),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3967),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_4026),
.B(n_123),
.Y(n_4064)
);

AOI221xp5_ASAP7_75t_L g4065 ( 
.A1(n_3983),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.C(n_129),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_4022),
.Y(n_4066)
);

NAND2xp33_ASAP7_75t_SL g4067 ( 
.A(n_3992),
.B(n_126),
.Y(n_4067)
);

OR2x2_ASAP7_75t_L g4068 ( 
.A(n_4040),
.B(n_127),
.Y(n_4068)
);

AOI21xp33_ASAP7_75t_L g4069 ( 
.A1(n_3970),
.A2(n_129),
.B(n_130),
.Y(n_4069)
);

OR2x2_ASAP7_75t_L g4070 ( 
.A(n_4029),
.B(n_4024),
.Y(n_4070)
);

A2O1A1Ixp33_ASAP7_75t_L g4071 ( 
.A1(n_4016),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3975),
.B(n_131),
.Y(n_4072)
);

NAND4xp25_ASAP7_75t_SL g4073 ( 
.A(n_3965),
.B(n_4001),
.C(n_3988),
.D(n_3973),
.Y(n_4073)
);

OR2x2_ASAP7_75t_L g4074 ( 
.A(n_4030),
.B(n_132),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_4002),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_4075)
);

AOI211xp5_ASAP7_75t_SL g4076 ( 
.A1(n_3979),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_3977),
.B(n_136),
.Y(n_4077)
);

HB1xp67_ASAP7_75t_L g4078 ( 
.A(n_4009),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3999),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_4028),
.Y(n_4080)
);

OAI221xp5_ASAP7_75t_L g4081 ( 
.A1(n_3995),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.C(n_140),
.Y(n_4081)
);

NOR2xp33_ASAP7_75t_L g4082 ( 
.A(n_4031),
.B(n_139),
.Y(n_4082)
);

AOI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_3986),
.A2(n_3997),
.B(n_4008),
.Y(n_4083)
);

O2A1O1Ixp33_ASAP7_75t_L g4084 ( 
.A1(n_4039),
.A2(n_145),
.B(n_140),
.C(n_142),
.Y(n_4084)
);

NAND3xp33_ASAP7_75t_L g4085 ( 
.A(n_3973),
.B(n_145),
.C(n_146),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3999),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3972),
.B(n_146),
.Y(n_4087)
);

OAI211xp5_ASAP7_75t_L g4088 ( 
.A1(n_3976),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_3981),
.B(n_149),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3985),
.B(n_151),
.Y(n_4090)
);

OAI22xp5_ASAP7_75t_L g4091 ( 
.A1(n_3976),
.A2(n_155),
.B1(n_152),
.B2(n_153),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_4019),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4004),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_4003),
.B(n_152),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3990),
.B(n_153),
.Y(n_4095)
);

AOI22xp5_ASAP7_75t_L g4096 ( 
.A1(n_4032),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_4012),
.B(n_156),
.Y(n_4097)
);

OAI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3987),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4034),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_4021),
.B(n_160),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_4027),
.B(n_160),
.Y(n_4101)
);

AOI322xp5_ASAP7_75t_L g4102 ( 
.A1(n_4042),
.A2(n_161),
.A3(n_162),
.B1(n_163),
.B2(n_164),
.C1(n_165),
.C2(n_166),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3968),
.B(n_161),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_3971),
.B(n_164),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_4007),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_4014),
.B(n_166),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4017),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_4013),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_4020),
.B(n_168),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_4025),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_4064),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_4049),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_4044),
.B(n_4036),
.Y(n_4113)
);

AND2x4_ASAP7_75t_L g4114 ( 
.A(n_4050),
.B(n_4056),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_4076),
.B(n_4053),
.Y(n_4115)
);

O2A1O1Ixp5_ASAP7_75t_L g4116 ( 
.A1(n_4075),
.A2(n_4000),
.B(n_3996),
.C(n_4010),
.Y(n_4116)
);

AOI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_4061),
.A2(n_3993),
.B1(n_3987),
.B2(n_4038),
.Y(n_4117)
);

INVx2_ASAP7_75t_SL g4118 ( 
.A(n_4070),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_4076),
.B(n_4018),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_4043),
.B(n_4023),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_4078),
.B(n_4006),
.Y(n_4121)
);

INVx3_ASAP7_75t_L g4122 ( 
.A(n_4079),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_4046),
.B(n_4093),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_4048),
.B(n_4041),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4086),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4047),
.Y(n_4126)
);

INVxp67_ASAP7_75t_SL g4127 ( 
.A(n_4054),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_4058),
.B(n_3994),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_4068),
.Y(n_4129)
);

OAI32xp33_ASAP7_75t_L g4130 ( 
.A1(n_4055),
.A2(n_4033),
.A3(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_4130)
);

AOI22xp5_ASAP7_75t_L g4131 ( 
.A1(n_4073),
.A2(n_173),
.B1(n_170),
.B2(n_172),
.Y(n_4131)
);

AOI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_4075),
.A2(n_175),
.B(n_176),
.Y(n_4132)
);

NOR3xp33_ASAP7_75t_L g4133 ( 
.A(n_4060),
.B(n_176),
.C(n_177),
.Y(n_4133)
);

OAI21xp33_ASAP7_75t_SL g4134 ( 
.A1(n_4062),
.A2(n_177),
.B(n_178),
.Y(n_4134)
);

INVx1_ASAP7_75t_SL g4135 ( 
.A(n_4067),
.Y(n_4135)
);

AOI22xp5_ASAP7_75t_L g4136 ( 
.A1(n_4045),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4077),
.Y(n_4137)
);

OAI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_4083),
.A2(n_179),
.B(n_180),
.Y(n_4138)
);

AOI221xp5_ASAP7_75t_L g4139 ( 
.A1(n_4062),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.C(n_186),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_4074),
.Y(n_4140)
);

AOI21xp33_ASAP7_75t_L g4141 ( 
.A1(n_4059),
.A2(n_186),
.B(n_187),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_4065),
.B(n_189),
.Y(n_4142)
);

OR2x2_ASAP7_75t_L g4143 ( 
.A(n_4087),
.B(n_190),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4094),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4052),
.B(n_190),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4104),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_4057),
.B(n_191),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_4051),
.B(n_191),
.Y(n_4148)
);

AOI21xp5_ASAP7_75t_L g4149 ( 
.A1(n_4098),
.A2(n_192),
.B(n_194),
.Y(n_4149)
);

INVx2_ASAP7_75t_SL g4150 ( 
.A(n_4105),
.Y(n_4150)
);

AOI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_4080),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_4151)
);

AOI32xp33_ASAP7_75t_L g4152 ( 
.A1(n_4098),
.A2(n_195),
.A3(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4089),
.Y(n_4153)
);

OAI22xp33_ASAP7_75t_SL g4154 ( 
.A1(n_4072),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_4063),
.Y(n_4155)
);

AOI221xp5_ASAP7_75t_L g4156 ( 
.A1(n_4051),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.C(n_207),
.Y(n_4156)
);

XNOR2x1_ASAP7_75t_SL g4157 ( 
.A(n_4066),
.B(n_205),
.Y(n_4157)
);

INVx2_ASAP7_75t_SL g4158 ( 
.A(n_4107),
.Y(n_4158)
);

OR2x2_ASAP7_75t_L g4159 ( 
.A(n_4085),
.B(n_206),
.Y(n_4159)
);

INVxp67_ASAP7_75t_L g4160 ( 
.A(n_4082),
.Y(n_4160)
);

AOI221xp5_ASAP7_75t_L g4161 ( 
.A1(n_4081),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.C(n_211),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_4092),
.B(n_208),
.Y(n_4162)
);

NAND2xp33_ASAP7_75t_L g4163 ( 
.A(n_4071),
.B(n_209),
.Y(n_4163)
);

OAI221xp5_ASAP7_75t_L g4164 ( 
.A1(n_4108),
.A2(n_4084),
.B1(n_4088),
.B2(n_4090),
.C(n_4099),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_4110),
.Y(n_4165)
);

OAI21xp5_ASAP7_75t_L g4166 ( 
.A1(n_4091),
.A2(n_211),
.B(n_212),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_4102),
.B(n_213),
.Y(n_4167)
);

INVx1_ASAP7_75t_SL g4168 ( 
.A(n_4097),
.Y(n_4168)
);

OR2x2_ASAP7_75t_L g4169 ( 
.A(n_4095),
.B(n_213),
.Y(n_4169)
);

OAI211xp5_ASAP7_75t_SL g4170 ( 
.A1(n_4069),
.A2(n_214),
.B(n_215),
.C(n_216),
.Y(n_4170)
);

OR2x2_ASAP7_75t_L g4171 ( 
.A(n_4101),
.B(n_214),
.Y(n_4171)
);

OAI221xp5_ASAP7_75t_L g4172 ( 
.A1(n_4091),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.C(n_219),
.Y(n_4172)
);

OAI21xp33_ASAP7_75t_L g4173 ( 
.A1(n_4103),
.A2(n_217),
.B(n_219),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_4096),
.B(n_220),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4157),
.B(n_4100),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_4114),
.B(n_4122),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4114),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_4127),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_SL g4179 ( 
.A(n_4134),
.B(n_4106),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4113),
.Y(n_4180)
);

AOI21xp33_ASAP7_75t_SL g4181 ( 
.A1(n_4118),
.A2(n_4109),
.B(n_220),
.Y(n_4181)
);

NAND4xp25_ASAP7_75t_L g4182 ( 
.A(n_4131),
.B(n_221),
.C(n_222),
.D(n_223),
.Y(n_4182)
);

NOR2xp33_ASAP7_75t_L g4183 ( 
.A(n_4135),
.B(n_223),
.Y(n_4183)
);

NOR2xp33_ASAP7_75t_L g4184 ( 
.A(n_4135),
.B(n_224),
.Y(n_4184)
);

INVx4_ASAP7_75t_SL g4185 ( 
.A(n_4112),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_4122),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4111),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4145),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_L g4189 ( 
.A(n_4119),
.B(n_225),
.Y(n_4189)
);

OAI21xp5_ASAP7_75t_SL g4190 ( 
.A1(n_4131),
.A2(n_227),
.B(n_228),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_4169),
.Y(n_4191)
);

OAI21xp33_ASAP7_75t_L g4192 ( 
.A1(n_4121),
.A2(n_227),
.B(n_228),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4147),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4123),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4125),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4162),
.Y(n_4196)
);

OAI221xp5_ASAP7_75t_L g4197 ( 
.A1(n_4138),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.C(n_233),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_SL g4198 ( 
.A(n_4134),
.B(n_229),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4137),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4171),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4144),
.B(n_233),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4146),
.Y(n_4202)
);

NOR2xp33_ASAP7_75t_SL g4203 ( 
.A(n_4164),
.B(n_234),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_4148),
.B(n_236),
.Y(n_4204)
);

NOR2xp33_ASAP7_75t_SL g4205 ( 
.A(n_4129),
.B(n_237),
.Y(n_4205)
);

NOR3xp33_ASAP7_75t_L g4206 ( 
.A(n_4124),
.B(n_4120),
.C(n_4141),
.Y(n_4206)
);

NOR3x1_ASAP7_75t_L g4207 ( 
.A(n_4115),
.B(n_237),
.C(n_238),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_L g4208 ( 
.A(n_4170),
.B(n_239),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4143),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4159),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_4173),
.B(n_239),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_L g4212 ( 
.A(n_4136),
.B(n_241),
.Y(n_4212)
);

NOR2xp33_ASAP7_75t_SL g4213 ( 
.A(n_4173),
.B(n_241),
.Y(n_4213)
);

NAND3xp33_ASAP7_75t_SL g4214 ( 
.A(n_4136),
.B(n_242),
.C(n_243),
.Y(n_4214)
);

AOI21xp5_ASAP7_75t_L g4215 ( 
.A1(n_4163),
.A2(n_242),
.B(n_244),
.Y(n_4215)
);

XOR2x2_ASAP7_75t_L g4216 ( 
.A(n_4133),
.B(n_245),
.Y(n_4216)
);

AOI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_4132),
.A2(n_245),
.B(n_246),
.Y(n_4217)
);

NOR3x1_ASAP7_75t_L g4218 ( 
.A(n_4167),
.B(n_246),
.C(n_247),
.Y(n_4218)
);

NAND3xp33_ASAP7_75t_SL g4219 ( 
.A(n_4117),
.B(n_247),
.C(n_249),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4139),
.B(n_250),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4140),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_4128),
.B(n_252),
.Y(n_4222)
);

NOR3xp33_ASAP7_75t_SL g4223 ( 
.A(n_4126),
.B(n_252),
.C(n_253),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4150),
.Y(n_4224)
);

OAI21xp33_ASAP7_75t_L g4225 ( 
.A1(n_4168),
.A2(n_254),
.B(n_255),
.Y(n_4225)
);

NOR2xp33_ASAP7_75t_L g4226 ( 
.A(n_4130),
.B(n_254),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_SL g4227 ( 
.A(n_4154),
.B(n_255),
.Y(n_4227)
);

AOI211xp5_ASAP7_75t_L g4228 ( 
.A1(n_4160),
.A2(n_256),
.B(n_257),
.C(n_258),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_4142),
.B(n_257),
.Y(n_4229)
);

XNOR2x2_ASAP7_75t_L g4230 ( 
.A(n_4156),
.B(n_258),
.Y(n_4230)
);

AOI21xp33_ASAP7_75t_SL g4231 ( 
.A1(n_4176),
.A2(n_4158),
.B(n_4166),
.Y(n_4231)
);

AOI211xp5_ASAP7_75t_L g4232 ( 
.A1(n_4181),
.A2(n_4154),
.B(n_4155),
.C(n_4165),
.Y(n_4232)
);

AOI22xp5_ASAP7_75t_L g4233 ( 
.A1(n_4203),
.A2(n_4161),
.B1(n_4153),
.B2(n_4174),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_4177),
.B(n_4152),
.Y(n_4234)
);

AOI221xp5_ASAP7_75t_L g4235 ( 
.A1(n_4219),
.A2(n_4116),
.B1(n_4149),
.B2(n_4172),
.C(n_4151),
.Y(n_4235)
);

NOR3xp33_ASAP7_75t_L g4236 ( 
.A(n_4178),
.B(n_259),
.C(n_260),
.Y(n_4236)
);

AOI221xp5_ASAP7_75t_L g4237 ( 
.A1(n_4189),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.C(n_264),
.Y(n_4237)
);

NAND4xp25_ASAP7_75t_L g4238 ( 
.A(n_4206),
.B(n_265),
.C(n_266),
.D(n_268),
.Y(n_4238)
);

OAI21xp33_ASAP7_75t_L g4239 ( 
.A1(n_4194),
.A2(n_265),
.B(n_266),
.Y(n_4239)
);

NOR2xp33_ASAP7_75t_R g4240 ( 
.A(n_4214),
.B(n_268),
.Y(n_4240)
);

NAND3xp33_ASAP7_75t_L g4241 ( 
.A(n_4213),
.B(n_269),
.C(n_270),
.Y(n_4241)
);

AOI221x1_ASAP7_75t_L g4242 ( 
.A1(n_4192),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.C(n_272),
.Y(n_4242)
);

AOI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_4224),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_4243)
);

NAND3xp33_ASAP7_75t_L g4244 ( 
.A(n_4198),
.B(n_274),
.C(n_277),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4185),
.Y(n_4245)
);

NOR3xp33_ASAP7_75t_L g4246 ( 
.A(n_4175),
.B(n_277),
.C(n_278),
.Y(n_4246)
);

OA33x2_ASAP7_75t_L g4247 ( 
.A1(n_4220),
.A2(n_280),
.A3(n_281),
.B1(n_282),
.B2(n_283),
.B3(n_284),
.Y(n_4247)
);

AOI211xp5_ASAP7_75t_SL g4248 ( 
.A1(n_4186),
.A2(n_4180),
.B(n_4183),
.C(n_4184),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_4185),
.Y(n_4249)
);

OAI21xp33_ASAP7_75t_L g4250 ( 
.A1(n_4221),
.A2(n_280),
.B(n_281),
.Y(n_4250)
);

NAND4xp25_ASAP7_75t_L g4251 ( 
.A(n_4218),
.B(n_282),
.C(n_283),
.D(n_285),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4185),
.B(n_285),
.Y(n_4252)
);

AOI211xp5_ASAP7_75t_SL g4253 ( 
.A1(n_4195),
.A2(n_286),
.B(n_287),
.C(n_290),
.Y(n_4253)
);

AOI221xp5_ASAP7_75t_L g4254 ( 
.A1(n_4227),
.A2(n_286),
.B1(n_287),
.B2(n_291),
.C(n_293),
.Y(n_4254)
);

OAI22xp33_ASAP7_75t_L g4255 ( 
.A1(n_4205),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_4190),
.B(n_295),
.Y(n_4256)
);

NAND5xp2_ASAP7_75t_L g4257 ( 
.A(n_4188),
.B(n_296),
.C(n_298),
.D(n_299),
.E(n_301),
.Y(n_4257)
);

INVxp67_ASAP7_75t_L g4258 ( 
.A(n_4211),
.Y(n_4258)
);

AOI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_4179),
.A2(n_302),
.B(n_303),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_4187),
.A2(n_4199),
.B1(n_4202),
.B2(n_4197),
.Y(n_4260)
);

OAI211xp5_ASAP7_75t_L g4261 ( 
.A1(n_4190),
.A2(n_302),
.B(n_303),
.C(n_304),
.Y(n_4261)
);

AOI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_4208),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_4262)
);

AOI22xp33_ASAP7_75t_L g4263 ( 
.A1(n_4193),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_4263)
);

AOI221xp5_ASAP7_75t_L g4264 ( 
.A1(n_4226),
.A2(n_307),
.B1(n_308),
.B2(n_310),
.C(n_311),
.Y(n_4264)
);

AOI211xp5_ASAP7_75t_L g4265 ( 
.A1(n_4222),
.A2(n_310),
.B(n_311),
.C(n_312),
.Y(n_4265)
);

AOI211xp5_ASAP7_75t_L g4266 ( 
.A1(n_4215),
.A2(n_312),
.B(n_313),
.C(n_314),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4201),
.B(n_313),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4196),
.B(n_314),
.Y(n_4268)
);

AOI221xp5_ASAP7_75t_L g4269 ( 
.A1(n_4210),
.A2(n_4182),
.B1(n_4200),
.B2(n_4209),
.C(n_4229),
.Y(n_4269)
);

OAI221xp5_ASAP7_75t_L g4270 ( 
.A1(n_4225),
.A2(n_315),
.B1(n_316),
.B2(n_332),
.C(n_334),
.Y(n_4270)
);

NAND3xp33_ASAP7_75t_SL g4271 ( 
.A(n_4217),
.B(n_335),
.C(n_336),
.Y(n_4271)
);

AOI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_4212),
.A2(n_339),
.B(n_340),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4204),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4252),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4245),
.Y(n_4275)
);

INVxp67_ASAP7_75t_SL g4276 ( 
.A(n_4249),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4256),
.Y(n_4277)
);

O2A1O1Ixp33_ASAP7_75t_SL g4278 ( 
.A1(n_4253),
.A2(n_4232),
.B(n_4261),
.C(n_4231),
.Y(n_4278)
);

INVxp33_ASAP7_75t_SL g4279 ( 
.A(n_4240),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4267),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4234),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4244),
.Y(n_4282)
);

AOI31xp33_ASAP7_75t_L g4283 ( 
.A1(n_4248),
.A2(n_4228),
.A3(n_4191),
.B(n_4207),
.Y(n_4283)
);

INVx2_ASAP7_75t_SL g4284 ( 
.A(n_4268),
.Y(n_4284)
);

OAI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_4262),
.A2(n_4223),
.B1(n_4230),
.B2(n_4216),
.Y(n_4285)
);

AO22x2_ASAP7_75t_L g4286 ( 
.A1(n_4260),
.A2(n_4182),
.B1(n_343),
.B2(n_345),
.Y(n_4286)
);

OAI22xp5_ASAP7_75t_L g4287 ( 
.A1(n_4233),
.A2(n_956),
.B1(n_946),
.B2(n_941),
.Y(n_4287)
);

BUFx2_ASAP7_75t_L g4288 ( 
.A(n_4251),
.Y(n_4288)
);

HB1xp67_ASAP7_75t_L g4289 ( 
.A(n_4253),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4241),
.Y(n_4290)
);

OAI22x1_ASAP7_75t_L g4291 ( 
.A1(n_4258),
.A2(n_342),
.B1(n_354),
.B2(n_358),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4239),
.Y(n_4292)
);

NAND4xp25_ASAP7_75t_SL g4293 ( 
.A(n_4235),
.B(n_359),
.C(n_362),
.D(n_364),
.Y(n_4293)
);

NOR2x1_ASAP7_75t_L g4294 ( 
.A(n_4238),
.B(n_365),
.Y(n_4294)
);

AOI221xp5_ASAP7_75t_L g4295 ( 
.A1(n_4269),
.A2(n_366),
.B1(n_369),
.B2(n_370),
.C(n_372),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_4273),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4243),
.Y(n_4297)
);

AOI22xp33_ASAP7_75t_SL g4298 ( 
.A1(n_4259),
.A2(n_375),
.B1(n_376),
.B2(n_381),
.Y(n_4298)
);

OAI22xp5_ASAP7_75t_L g4299 ( 
.A1(n_4265),
.A2(n_956),
.B1(n_946),
.B2(n_941),
.Y(n_4299)
);

A2O1A1Ixp33_ASAP7_75t_L g4300 ( 
.A1(n_4276),
.A2(n_4254),
.B(n_4264),
.C(n_4246),
.Y(n_4300)
);

OAI21xp33_ASAP7_75t_L g4301 ( 
.A1(n_4279),
.A2(n_4257),
.B(n_4271),
.Y(n_4301)
);

NOR3xp33_ASAP7_75t_L g4302 ( 
.A(n_4283),
.B(n_4250),
.C(n_4270),
.Y(n_4302)
);

AOI211xp5_ASAP7_75t_SL g4303 ( 
.A1(n_4278),
.A2(n_4255),
.B(n_4272),
.C(n_4266),
.Y(n_4303)
);

NOR2xp33_ASAP7_75t_L g4304 ( 
.A(n_4289),
.B(n_4236),
.Y(n_4304)
);

AOI22xp5_ASAP7_75t_L g4305 ( 
.A1(n_4281),
.A2(n_4237),
.B1(n_4263),
.B2(n_4247),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4286),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_4275),
.B(n_4242),
.Y(n_4307)
);

OAI21xp5_ASAP7_75t_L g4308 ( 
.A1(n_4294),
.A2(n_386),
.B(n_387),
.Y(n_4308)
);

OAI211xp5_ASAP7_75t_SL g4309 ( 
.A1(n_4292),
.A2(n_388),
.B(n_389),
.C(n_392),
.Y(n_4309)
);

OAI31xp33_ASAP7_75t_L g4310 ( 
.A1(n_4285),
.A2(n_4286),
.A3(n_4293),
.B(n_4288),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4294),
.Y(n_4311)
);

AOI211xp5_ASAP7_75t_L g4312 ( 
.A1(n_4290),
.A2(n_393),
.B(n_396),
.C(n_397),
.Y(n_4312)
);

AOI211xp5_ASAP7_75t_L g4313 ( 
.A1(n_4282),
.A2(n_398),
.B(n_401),
.C(n_405),
.Y(n_4313)
);

AOI211x1_ASAP7_75t_SL g4314 ( 
.A1(n_4297),
.A2(n_406),
.B(n_408),
.C(n_410),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4274),
.B(n_415),
.Y(n_4315)
);

AOI21xp5_ASAP7_75t_L g4316 ( 
.A1(n_4307),
.A2(n_4296),
.B(n_4284),
.Y(n_4316)
);

INVx2_ASAP7_75t_SL g4317 ( 
.A(n_4311),
.Y(n_4317)
);

XNOR2xp5_ASAP7_75t_L g4318 ( 
.A(n_4305),
.B(n_4302),
.Y(n_4318)
);

NOR2xp33_ASAP7_75t_SL g4319 ( 
.A(n_4301),
.B(n_4277),
.Y(n_4319)
);

OAI221xp5_ASAP7_75t_L g4320 ( 
.A1(n_4310),
.A2(n_4298),
.B1(n_4295),
.B2(n_4280),
.C(n_4299),
.Y(n_4320)
);

OAI211xp5_ASAP7_75t_SL g4321 ( 
.A1(n_4303),
.A2(n_4287),
.B(n_4291),
.C(n_419),
.Y(n_4321)
);

OAI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_4306),
.A2(n_956),
.B1(n_946),
.B2(n_941),
.Y(n_4322)
);

NOR3xp33_ASAP7_75t_SL g4323 ( 
.A(n_4304),
.B(n_417),
.C(n_418),
.Y(n_4323)
);

OAI221xp5_ASAP7_75t_SL g4324 ( 
.A1(n_4300),
.A2(n_420),
.B1(n_421),
.B2(n_423),
.C(n_424),
.Y(n_4324)
);

OAI21xp5_ASAP7_75t_SL g4325 ( 
.A1(n_4314),
.A2(n_429),
.B(n_431),
.Y(n_4325)
);

O2A1O1Ixp5_ASAP7_75t_L g4326 ( 
.A1(n_4308),
.A2(n_434),
.B(n_436),
.C(n_438),
.Y(n_4326)
);

OAI32xp33_ASAP7_75t_L g4327 ( 
.A1(n_4321),
.A2(n_4315),
.A3(n_4309),
.B1(n_4313),
.B2(n_4312),
.Y(n_4327)
);

AOI22xp5_ASAP7_75t_L g4328 ( 
.A1(n_4319),
.A2(n_938),
.B1(n_946),
.B2(n_956),
.Y(n_4328)
);

AOI221xp5_ASAP7_75t_L g4329 ( 
.A1(n_4317),
.A2(n_439),
.B1(n_440),
.B2(n_442),
.C(n_443),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4318),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4325),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4323),
.B(n_444),
.Y(n_4332)
);

AOI22xp5_ASAP7_75t_L g4333 ( 
.A1(n_4320),
.A2(n_938),
.B1(n_955),
.B2(n_949),
.Y(n_4333)
);

AND3x4_ASAP7_75t_L g4334 ( 
.A(n_4327),
.B(n_4316),
.C(n_4326),
.Y(n_4334)
);

NAND2x1p5_ASAP7_75t_L g4335 ( 
.A(n_4332),
.B(n_4324),
.Y(n_4335)
);

NAND5xp2_ASAP7_75t_L g4336 ( 
.A(n_4330),
.B(n_4331),
.C(n_4333),
.D(n_4328),
.E(n_4329),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4332),
.Y(n_4337)
);

NOR4xp75_ASAP7_75t_SL g4338 ( 
.A(n_4330),
.B(n_4322),
.C(n_447),
.D(n_450),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4332),
.Y(n_4339)
);

NOR3xp33_ASAP7_75t_L g4340 ( 
.A(n_4336),
.B(n_446),
.C(n_451),
.Y(n_4340)
);

CKINVDCx16_ASAP7_75t_R g4341 ( 
.A(n_4337),
.Y(n_4341)
);

AO22x1_ASAP7_75t_L g4342 ( 
.A1(n_4334),
.A2(n_453),
.B1(n_455),
.B2(n_457),
.Y(n_4342)
);

AND3x4_ASAP7_75t_L g4343 ( 
.A(n_4340),
.B(n_4338),
.C(n_4335),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4342),
.Y(n_4344)
);

AND3x1_ASAP7_75t_L g4345 ( 
.A(n_4341),
.B(n_4339),
.C(n_459),
.Y(n_4345)
);

OAI22xp5_ASAP7_75t_L g4346 ( 
.A1(n_4343),
.A2(n_458),
.B1(n_460),
.B2(n_462),
.Y(n_4346)
);

AO22x2_ASAP7_75t_L g4347 ( 
.A1(n_4346),
.A2(n_4344),
.B1(n_4345),
.B2(n_469),
.Y(n_4347)
);

OAI22xp5_ASAP7_75t_SL g4348 ( 
.A1(n_4347),
.A2(n_465),
.B1(n_467),
.B2(n_1268),
.Y(n_4348)
);

AOI31xp33_ASAP7_75t_L g4349 ( 
.A1(n_4348),
.A2(n_1476),
.A3(n_942),
.B(n_938),
.Y(n_4349)
);

OAI22xp5_ASAP7_75t_SL g4350 ( 
.A1(n_4349),
.A2(n_1248),
.B1(n_1175),
.B2(n_1163),
.Y(n_4350)
);

AOI22xp33_ASAP7_75t_L g4351 ( 
.A1(n_4350),
.A2(n_955),
.B1(n_940),
.B2(n_943),
.Y(n_4351)
);

NOR2xp33_ASAP7_75t_L g4352 ( 
.A(n_4351),
.B(n_955),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4352),
.Y(n_4353)
);

OAI221xp5_ASAP7_75t_L g4354 ( 
.A1(n_4353),
.A2(n_955),
.B1(n_940),
.B2(n_943),
.C(n_949),
.Y(n_4354)
);

OR2x6_ASAP7_75t_L g4355 ( 
.A(n_4353),
.B(n_1163),
.Y(n_4355)
);

AOI221xp5_ASAP7_75t_L g4356 ( 
.A1(n_4354),
.A2(n_955),
.B1(n_943),
.B2(n_949),
.C(n_1163),
.Y(n_4356)
);

AOI211xp5_ASAP7_75t_L g4357 ( 
.A1(n_4356),
.A2(n_4355),
.B(n_943),
.C(n_949),
.Y(n_4357)
);


endmodule