module fake_jpeg_5126_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_20),
.CON(n_52),
.SN(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_31),
.B1(n_24),
.B2(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_57),
.B1(n_62),
.B2(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_25),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_50),
.B(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_R g73 ( 
.A(n_52),
.B(n_38),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_31),
.B1(n_24),
.B2(n_29),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_31),
.B1(n_24),
.B2(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_42),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_34),
.B1(n_33),
.B2(n_17),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_17),
.B1(n_19),
.B2(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_44),
.C(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_77),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_9),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_84),
.B(n_79),
.C(n_28),
.Y(n_121)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_39),
.B1(n_59),
.B2(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_35),
.Y(n_113)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_112),
.B1(n_117),
.B2(n_93),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_120),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_69),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_107),
.Y(n_141)
);

INVx2_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_32),
.C(n_27),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_114),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_43),
.B1(n_61),
.B2(n_40),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_40),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_43),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_74),
.C(n_88),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_43),
.B1(n_46),
.B2(n_64),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_94),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_77),
.B1(n_85),
.B2(n_19),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_22),
.Y(n_150)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_78),
.B1(n_70),
.B2(n_51),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_127),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_129),
.B1(n_148),
.B2(n_151),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_60),
.B1(n_96),
.B2(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_144),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_48),
.B1(n_96),
.B2(n_82),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_136),
.B1(n_139),
.B2(n_143),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_96),
.B1(n_82),
.B2(n_80),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_137),
.B(n_140),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_108),
.C(n_121),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_90),
.B1(n_76),
.B2(n_74),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_145),
.C(n_149),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_21),
.B1(n_41),
.B2(n_23),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_34),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_146),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_97),
.A2(n_103),
.B1(n_122),
.B2(n_106),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_88),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_99),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_23),
.B1(n_27),
.B2(n_65),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_98),
.B1(n_118),
.B2(n_115),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_103),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_141),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_157),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_103),
.B(n_105),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_161),
.B(n_130),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_105),
.B(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_105),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_171),
.C(n_180),
.Y(n_199)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_173),
.Y(n_185)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_118),
.C(n_119),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_100),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_143),
.B1(n_147),
.B2(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_65),
.B1(n_18),
.B2(n_26),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_126),
.B1(n_75),
.B2(n_130),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_36),
.C(n_35),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_197),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_184),
.A2(n_207),
.B1(n_177),
.B2(n_170),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_194),
.B(n_203),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_141),
.B(n_134),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_36),
.C(n_95),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_0),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_159),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_201),
.C(n_205),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_36),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_181),
.A2(n_36),
.B(n_95),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_123),
.C(n_86),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_75),
.B1(n_86),
.B2(n_30),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_0),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g212 ( 
.A(n_208),
.B(n_209),
.CI(n_167),
.CON(n_212),
.SN(n_212)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_154),
.B(n_1),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_163),
.B1(n_162),
.B2(n_155),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_123),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_213),
.B(n_222),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_180),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_228),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_195),
.B(n_168),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_9),
.C(n_15),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_189),
.A2(n_197),
.B1(n_204),
.B2(n_203),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_219),
.A2(n_234),
.B1(n_192),
.B2(n_185),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_153),
.B1(n_165),
.B2(n_156),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_189),
.B(n_156),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_227),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_195),
.A2(n_190),
.B1(n_196),
.B2(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_177),
.C(n_166),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_230),
.C(n_231),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_177),
.B1(n_75),
.B2(n_30),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_187),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_30),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_201),
.C(n_205),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_30),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_191),
.A2(n_30),
.B1(n_26),
.B2(n_18),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_26),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_185),
.B(n_208),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_198),
.B(n_202),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_186),
.A2(n_26),
.B1(n_18),
.B2(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

AO221x1_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_187),
.B1(n_192),
.B2(n_26),
.C(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_245),
.B(n_249),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_209),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_188),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_255),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_252),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_184),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_1),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_254),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_233),
.B1(n_220),
.B2(n_219),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_251),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_211),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_230),
.B1(n_212),
.B2(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_212),
.B1(n_214),
.B2(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_218),
.C(n_216),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_266),
.C(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_228),
.C(n_234),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_9),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_241),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_248),
.A2(n_10),
.B1(n_15),
.B2(n_4),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_271),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_2),
.C(n_3),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_244),
.C(n_245),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_242),
.A2(n_16),
.B1(n_8),
.B2(n_4),
.Y(n_271)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_276),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_277),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_242),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_236),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_283),
.C(n_284),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_247),
.B(n_253),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_258),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_255),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_241),
.C(n_249),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_243),
.C(n_235),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_293),
.B1(n_294),
.B2(n_275),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_257),
.B1(n_278),
.B2(n_283),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_6),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_261),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_292),
.B(n_11),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_266),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_3),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_270),
.B1(n_269),
.B2(n_267),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_261),
.B1(n_246),
.B2(n_2),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_11),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_272),
.C(n_5),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_6),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_302),
.C(n_303),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_11),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_299),
.B(n_301),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_5),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_287),
.B(n_290),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_307),
.B(n_308),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_286),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_8),
.C(n_12),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_13),
.C(n_14),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_311),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_312),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_304),
.Y(n_315)
);


endmodule