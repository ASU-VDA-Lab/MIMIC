module fake_jpeg_11299_n_621 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_621);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_621;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_11),
.B(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_64),
.B(n_65),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_17),
.C(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_67),
.B(n_68),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_37),
.B(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_75),
.B(n_90),
.Y(n_197)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_78),
.Y(n_206)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_79),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_12),
.B1(n_11),
.B2(n_9),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_81),
.A2(n_36),
.B1(n_52),
.B2(n_51),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_83),
.B(n_124),
.Y(n_186)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_18),
.B(n_12),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_91),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_93),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_12),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_94),
.B(n_104),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_98),
.Y(n_187)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_11),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_19),
.B(n_9),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_115),
.B(n_126),
.Y(n_202)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_53),
.Y(n_124)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_8),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_60),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_127),
.B(n_132),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_83),
.A2(n_33),
.B(n_30),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_77),
.B(n_20),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_139),
.B(n_148),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_140),
.A2(n_190),
.B1(n_50),
.B2(n_46),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_62),
.B(n_26),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_26),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_161),
.B(n_162),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_102),
.A2(n_36),
.B(n_27),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_48),
.B1(n_28),
.B2(n_52),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_167),
.A2(n_169),
.B1(n_199),
.B2(n_40),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_48),
.B1(n_28),
.B2(n_27),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_82),
.B(n_51),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_170),
.B(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_74),
.Y(n_185)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_82),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_66),
.A2(n_29),
.B1(n_32),
.B2(n_54),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_88),
.B(n_33),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_124),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_89),
.B(n_30),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_193),
.B(n_114),
.Y(n_256)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_105),
.A2(n_54),
.B1(n_29),
.B2(n_50),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_69),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_210),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_211),
.A2(n_133),
.B1(n_137),
.B2(n_69),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_212),
.B(n_218),
.Y(n_288)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_214),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_215),
.Y(n_299)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_216),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_220),
.B(n_256),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_223),
.A2(n_225),
.B1(n_232),
.B2(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_40),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_224),
.B(n_227),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_157),
.A2(n_198),
.B1(n_202),
.B2(n_182),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_91),
.B1(n_85),
.B2(n_92),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_226),
.A2(n_278),
.B1(n_207),
.B2(n_191),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_127),
.B(n_49),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_151),
.A2(n_108),
.B1(n_56),
.B2(n_60),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_134),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_229),
.Y(n_307)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_231),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_119),
.B1(n_113),
.B2(n_112),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_267),
.Y(n_298)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_235),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_166),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_240),
.Y(n_301)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_156),
.Y(n_237)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_130),
.Y(n_238)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_144),
.Y(n_239)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_132),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_241),
.Y(n_315)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_156),
.Y(n_243)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_151),
.A2(n_60),
.B1(n_56),
.B2(n_59),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_246),
.A2(n_248),
.B1(n_265),
.B2(n_268),
.Y(n_305)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_128),
.Y(n_247)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_131),
.A2(n_59),
.B1(n_46),
.B2(n_98),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_165),
.Y(n_250)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_163),
.Y(n_252)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_252),
.Y(n_322)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_254),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_110),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_54),
.C(n_195),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_186),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_257),
.B(n_259),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

INVx11_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_173),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_176),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_260),
.B(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_177),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_263),
.Y(n_311)
);

BUFx4f_ASAP7_75t_L g264 ( 
.A(n_145),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_165),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_197),
.A2(n_111),
.B1(n_107),
.B2(n_29),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_197),
.A2(n_86),
.B(n_96),
.C(n_142),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_135),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_270),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_141),
.A2(n_49),
.B1(n_44),
.B2(n_42),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_271),
.A2(n_273),
.B1(n_0),
.B2(n_2),
.Y(n_333)
);

BUFx4f_ASAP7_75t_SL g272 ( 
.A(n_203),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_272),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_146),
.A2(n_42),
.B1(n_34),
.B2(n_44),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_173),
.A2(n_63),
.B(n_96),
.C(n_58),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_103),
.B(n_172),
.Y(n_285)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_164),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_280),
.Y(n_318)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_171),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_277),
.Y(n_330)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_194),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_147),
.B(n_58),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_279),
.B(n_168),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_136),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_138),
.B(n_34),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_282),
.Y(n_337)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_129),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_211),
.A2(n_149),
.B1(n_154),
.B2(n_178),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_283),
.A2(n_284),
.B1(n_320),
.B2(n_274),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_249),
.A2(n_207),
.B1(n_191),
.B2(n_138),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_285),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_291),
.A2(n_314),
.B1(n_321),
.B2(n_335),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_293),
.B(n_321),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_143),
.C(n_206),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_316),
.C(n_323),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_312),
.B(n_272),
.Y(n_369)
);

OAI22x1_ASAP7_75t_R g313 ( 
.A1(n_262),
.A2(n_79),
.B1(n_184),
.B2(n_187),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g387 ( 
.A1(n_313),
.A2(n_329),
.B(n_309),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_206),
.B1(n_54),
.B2(n_150),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_224),
.B(n_174),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_262),
.A2(n_106),
.B1(n_101),
.B2(n_97),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_262),
.B(n_86),
.C(n_95),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_227),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_325),
.A2(n_326),
.B(n_336),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_220),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_333),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_232),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_267),
.A2(n_0),
.B(n_3),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_213),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_338),
.A2(n_339),
.B1(n_265),
.B2(n_268),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_281),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_242),
.A2(n_5),
.B1(n_6),
.B2(n_234),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_330),
.Y(n_343)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_343),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_295),
.A2(n_230),
.B1(n_216),
.B2(n_269),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_345),
.A2(n_352),
.B1(n_355),
.B2(n_363),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_324),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_349),
.Y(n_395)
);

OAI22xp33_ASAP7_75t_SL g424 ( 
.A1(n_348),
.A2(n_289),
.B1(n_290),
.B2(n_296),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_324),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_247),
.B(n_244),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_350),
.A2(n_313),
.B(n_318),
.Y(n_388)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_295),
.A2(n_221),
.B1(n_233),
.B2(n_217),
.Y(n_352)
);

OAI32xp33_ASAP7_75t_L g354 ( 
.A1(n_298),
.A2(n_209),
.A3(n_231),
.B1(n_210),
.B2(n_214),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_354),
.B(n_357),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_298),
.A2(n_243),
.B1(n_237),
.B2(n_250),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_359),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_254),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_361),
.B(n_377),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_283),
.A2(n_284),
.B1(n_337),
.B2(n_308),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_362),
.A2(n_365),
.B1(n_367),
.B2(n_371),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g364 ( 
.A1(n_297),
.A2(n_260),
.A3(n_276),
.B1(n_277),
.B2(n_222),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_366),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_293),
.A2(n_241),
.B1(n_280),
.B2(n_253),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_316),
.B(n_219),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_285),
.A2(n_253),
.B1(n_215),
.B2(n_218),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_287),
.B(n_5),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_368),
.B(n_370),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_369),
.B(n_379),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_297),
.B(n_229),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_331),
.A2(n_222),
.B1(n_275),
.B2(n_245),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_373),
.B(n_333),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_314),
.A2(n_278),
.B1(n_222),
.B2(n_258),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_374),
.A2(n_376),
.B1(n_378),
.B2(n_381),
.Y(n_394)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_291),
.A2(n_264),
.B1(n_278),
.B2(n_272),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_324),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_331),
.A2(n_264),
.B1(n_340),
.B2(n_305),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_286),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_286),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_380),
.B(n_382),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_335),
.A2(n_301),
.B1(n_339),
.B2(n_326),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_299),
.B(n_312),
.Y(n_382)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_383),
.A2(n_384),
.B1(n_290),
.B2(n_302),
.Y(n_425)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_292),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_325),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_315),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_332),
.A2(n_323),
.B1(n_313),
.B2(n_318),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_386),
.A2(n_329),
.B1(n_311),
.B2(n_315),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_387),
.A2(n_307),
.B(n_334),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_388),
.A2(n_413),
.B(n_421),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_357),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_389),
.B(n_412),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_288),
.C(n_292),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_390),
.B(n_401),
.C(n_405),
.Y(n_438)
);

XNOR2x1_ASAP7_75t_SL g391 ( 
.A(n_358),
.B(n_313),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_386),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_396),
.B(n_381),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_347),
.A2(n_318),
.B1(n_328),
.B2(n_319),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_399),
.A2(n_402),
.B1(n_417),
.B2(n_420),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_358),
.B(n_319),
.C(n_322),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_348),
.A2(n_306),
.B1(n_303),
.B2(n_322),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_403),
.A2(n_408),
.B(n_371),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_311),
.C(n_300),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_300),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_409),
.C(n_410),
.Y(n_447)
);

OAI21xp33_ASAP7_75t_SL g408 ( 
.A1(n_385),
.A2(n_307),
.B(n_289),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_294),
.C(n_304),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_294),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_382),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_360),
.A2(n_304),
.B(n_334),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_369),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_415),
.B(n_419),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_362),
.A2(n_306),
.B1(n_310),
.B2(n_317),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_342),
.A2(n_317),
.B1(n_303),
.B2(n_296),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_352),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_422),
.B(n_354),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_424),
.A2(n_374),
.B1(n_376),
.B2(n_355),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_425),
.Y(n_431)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_427),
.Y(n_463)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_398),
.Y(n_429)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_423),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_430),
.B(n_437),
.Y(n_474)
);

XOR2x1_ASAP7_75t_L g481 ( 
.A(n_432),
.B(n_441),
.Y(n_481)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_434),
.Y(n_484)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_420),
.Y(n_436)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_436),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_439),
.A2(n_426),
.B1(n_435),
.B2(n_403),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_423),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_454),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_343),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_389),
.B(n_418),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_442),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_414),
.A2(n_360),
.B1(n_365),
.B2(n_345),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_456),
.B1(n_400),
.B2(n_414),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_368),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_451),
.C(n_391),
.Y(n_464)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_412),
.B(n_418),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_449),
.B(n_452),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_393),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_450),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_401),
.B(n_377),
.C(n_346),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_413),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_406),
.B(n_349),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_453),
.B(n_457),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_406),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_455),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_394),
.A2(n_350),
.B1(n_344),
.B2(n_367),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_392),
.B(n_364),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_419),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_387),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_459),
.A2(n_460),
.B(n_388),
.Y(n_466)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_393),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_461),
.B(n_395),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_467),
.C(n_446),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_443),
.B(n_459),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_390),
.C(n_409),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_468),
.A2(n_480),
.B1(n_482),
.B2(n_485),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_396),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_469),
.B(n_472),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_396),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_450),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_478),
.B(n_491),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_435),
.A2(n_394),
.B1(n_411),
.B2(n_426),
.Y(n_479)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_479),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_456),
.A2(n_400),
.B1(n_402),
.B2(n_411),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_445),
.A2(n_417),
.B1(n_344),
.B2(n_378),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_458),
.A2(n_408),
.B1(n_410),
.B2(n_399),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_489),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_459),
.A2(n_415),
.B1(n_353),
.B2(n_405),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_488),
.A2(n_493),
.B(n_452),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_438),
.B(n_395),
.Y(n_489)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_490),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_449),
.B(n_416),
.Y(n_491)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_492),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_458),
.A2(n_363),
.B1(n_416),
.B2(n_350),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_494),
.A2(n_498),
.B(n_510),
.Y(n_533)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_473),
.Y(n_497)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_497),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_466),
.A2(n_443),
.B(n_459),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_463),
.Y(n_499)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_499),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_451),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_503),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_467),
.B(n_432),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_505),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_433),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_507),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_433),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_464),
.B(n_444),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_508),
.B(n_521),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_465),
.A2(n_444),
.B(n_431),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_511),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_474),
.A2(n_460),
.B(n_437),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_516),
.Y(n_524)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_471),
.Y(n_513)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_513),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_SL g514 ( 
.A1(n_486),
.A2(n_436),
.B(n_439),
.C(n_431),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_514),
.Y(n_541)
);

A2O1A1Ixp33_ASAP7_75t_SL g515 ( 
.A1(n_486),
.A2(n_441),
.B(n_457),
.C(n_428),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_515),
.A2(n_475),
.B1(n_462),
.B2(n_430),
.Y(n_540)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_518),
.B(n_520),
.Y(n_539)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_477),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_442),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_476),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_522),
.A2(n_484),
.B1(n_461),
.B2(n_429),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_481),
.C(n_488),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_525),
.B(n_530),
.Y(n_547)
);

XNOR2x1_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_481),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_528),
.B(n_543),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_485),
.C(n_493),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_509),
.A2(n_468),
.B1(n_480),
.B2(n_482),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_534),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_521),
.B(n_474),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_542),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_501),
.B(n_505),
.C(n_496),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_538),
.B(n_546),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_540),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_483),
.Y(n_542)
);

XNOR2x1_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_479),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_517),
.A2(n_440),
.B1(n_454),
.B2(n_427),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_544),
.A2(n_512),
.B1(n_509),
.B2(n_500),
.Y(n_549)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_545),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_496),
.B(n_453),
.C(n_470),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_549),
.A2(n_541),
.B1(n_533),
.B2(n_530),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_544),
.A2(n_495),
.B1(n_500),
.B2(n_519),
.Y(n_550)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_550),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_529),
.B(n_507),
.C(n_504),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_551),
.B(n_554),
.Y(n_568)
);

A2O1A1Ixp33_ASAP7_75t_SL g552 ( 
.A1(n_541),
.A2(n_498),
.B(n_494),
.C(n_514),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_552),
.B(n_556),
.C(n_564),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_523),
.B(n_384),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_529),
.B(n_517),
.C(n_510),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_539),
.Y(n_557)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_557),
.Y(n_576)
);

BUFx24_ASAP7_75t_SL g560 ( 
.A(n_537),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_560),
.B(n_546),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_525),
.A2(n_514),
.B1(n_470),
.B2(n_484),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_561),
.B(n_533),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_455),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_562),
.B(n_547),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_538),
.B(n_514),
.C(n_515),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_540),
.Y(n_565)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_565),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_566),
.B(n_571),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_570),
.B(n_552),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_537),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_573),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_532),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_536),
.C(n_532),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_575),
.B(n_580),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_563),
.Y(n_588)
);

INVx11_ASAP7_75t_L g578 ( 
.A(n_553),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_578),
.B(n_526),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_524),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_579),
.A2(n_581),
.B(n_582),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_535),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_558),
.B(n_527),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_551),
.B(n_536),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_574),
.A2(n_548),
.B1(n_552),
.B2(n_543),
.Y(n_584)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_584),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_586),
.B(n_587),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_569),
.A2(n_548),
.B1(n_531),
.B2(n_515),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_588),
.B(n_589),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_574),
.B(n_552),
.C(n_563),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_568),
.B(n_528),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_590),
.B(n_591),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_572),
.B(n_570),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_592),
.B(n_383),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_576),
.A2(n_515),
.B1(n_434),
.B2(n_448),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_594),
.B(n_577),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_SL g597 ( 
.A1(n_595),
.A2(n_579),
.B(n_581),
.C(n_567),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_597),
.B(n_602),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_589),
.A2(n_567),
.B1(n_578),
.B2(n_575),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_599),
.B(n_604),
.Y(n_607)
);

AOI21xp33_ASAP7_75t_L g603 ( 
.A1(n_585),
.A2(n_573),
.B(n_380),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_603),
.A2(n_351),
.B(n_356),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_593),
.B(n_379),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_605),
.B(n_588),
.C(n_583),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_606),
.B(n_610),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_583),
.C(n_592),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_608),
.A2(n_611),
.B(n_600),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_601),
.A2(n_591),
.B1(n_584),
.B2(n_590),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_609),
.A2(n_599),
.B(n_596),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_612),
.A2(n_613),
.B(n_615),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_609),
.A2(n_597),
.B(n_361),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_614),
.B(n_607),
.C(n_375),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_616),
.A2(n_359),
.B(n_372),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_618),
.B(n_617),
.C(n_372),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_619),
.B(n_383),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g621 ( 
.A(n_620),
.B(n_302),
.Y(n_621)
);


endmodule