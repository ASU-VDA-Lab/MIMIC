module fake_ibex_1946_n_677 (n_85, n_84, n_64, n_3, n_73, n_65, n_95, n_55, n_63, n_98, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_97, n_15, n_24, n_52, n_99, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_96, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_677);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_95;
input n_55;
input n_63;
input n_98;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_97;
input n_15;
input n_24;
input n_52;
input n_99;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_96;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_677;

wire n_151;
wire n_599;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_652;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_645;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_105;
wire n_187;
wire n_667;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_673;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_122;
wire n_523;
wire n_116;
wire n_614;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_136;
wire n_261;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_437;
wire n_602;
wire n_355;
wire n_474;
wire n_594;
wire n_636;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_676;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_643;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_672;
wire n_401;
wire n_553;
wire n_554;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_605;
wire n_539;
wire n_100;
wire n_179;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_411;
wire n_135;
wire n_520;
wire n_658;
wire n_512;
wire n_615;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_627;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_650;
wire n_409;
wire n_582;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_633;
wire n_532;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_385;
wire n_233;
wire n_342;
wire n_414;
wire n_430;
wire n_118;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_639;
wire n_303;
wire n_362;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_668;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_631;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_160;
wire n_657;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_45),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_49),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_2),
.B(n_53),
.Y(n_110)
);

BUFx2_ASAP7_75t_SL g111 ( 
.A(n_57),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_54),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_11),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_13),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_12),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_24),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_22),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_0),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_23),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_28),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_79),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_63),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_14),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_26),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_30),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_16),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_14),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_23),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_43),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_86),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_61),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_76),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_40),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_90),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_4),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_22),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_8),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_50),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_27),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_47),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_31),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_32),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_6),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_92),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_11),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_2),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_17),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_44),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_L g165 ( 
.A(n_38),
.B(n_71),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_21),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_36),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_39),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_59),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_52),
.B(n_68),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_93),
.B(n_64),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_8),
.Y(n_173)
);

NOR2xp67_ASAP7_75t_L g174 ( 
.A(n_80),
.B(n_6),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_10),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_65),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_157),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_136),
.B(n_3),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_116),
.A2(n_46),
.B(n_95),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_116),
.B(n_5),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_7),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_121),
.B(n_48),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_112),
.B(n_10),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_113),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g209 ( 
.A(n_123),
.B(n_13),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_115),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_128),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_156),
.B(n_18),
.Y(n_220)
);

OA21x2_ASAP7_75t_L g221 ( 
.A1(n_135),
.A2(n_69),
.B(n_94),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_155),
.A2(n_67),
.B(n_88),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_119),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_103),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_105),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_141),
.B(n_20),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_170),
.B(n_120),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_124),
.B(n_20),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_143),
.B(n_176),
.Y(n_235)
);

AND2x6_ASAP7_75t_L g236 ( 
.A(n_126),
.B(n_62),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_134),
.B(n_21),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_140),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_151),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_164),
.B(n_25),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_167),
.B(n_29),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_169),
.B(n_34),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_111),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_122),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_110),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_128),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_109),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_190),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_191),
.B(n_145),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_182),
.B(n_133),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_190),
.B(n_137),
.C(n_166),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_222),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_185),
.B1(n_191),
.B2(n_195),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_195),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_187),
.B(n_146),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_177),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

CKINVDCx11_ASAP7_75t_R g274 ( 
.A(n_204),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_241),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_241),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_187),
.B(n_173),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_131),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_207),
.B(n_130),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_243),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_207),
.B(n_144),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_207),
.B(n_153),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_150),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_240),
.A2(n_107),
.B1(n_168),
.B2(n_132),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_236),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_225),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_248),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_214),
.B(n_154),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_196),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_214),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_196),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_212),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_214),
.B(n_160),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_236),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_179),
.Y(n_302)
);

NOR2x1p5_ASAP7_75t_L g303 ( 
.A(n_235),
.B(n_149),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_196),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_237),
.B(n_209),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_197),
.B(n_125),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_244),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_209),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_208),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_208),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_245),
.B(n_172),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_215),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_181),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_181),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

OR2x6_ASAP7_75t_L g317 ( 
.A(n_216),
.B(n_171),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_215),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_245),
.B(n_142),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_183),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_183),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_183),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_183),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_193),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_189),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_189),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_217),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_226),
.B(n_138),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_219),
.B(n_161),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_189),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_189),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

AND3x1_ASAP7_75t_L g333 ( 
.A(n_286),
.B(n_203),
.C(n_231),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_L g334 ( 
.A(n_250),
.B(n_236),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_275),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_252),
.B(n_245),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_256),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_283),
.B(n_232),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_329),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_256),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_274),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_257),
.B(n_227),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

AO22x2_ASAP7_75t_L g345 ( 
.A1(n_287),
.A2(n_184),
.B1(n_237),
.B2(n_193),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_299),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_193),
.B(n_213),
.C(n_218),
.Y(n_347)
);

OR2x6_ASAP7_75t_L g348 ( 
.A(n_250),
.B(n_237),
.Y(n_348)
);

OAI221xp5_ASAP7_75t_L g349 ( 
.A1(n_264),
.A2(n_199),
.B1(n_227),
.B2(n_230),
.C(n_239),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_324),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_280),
.B(n_230),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_305),
.A2(n_132),
.B1(n_107),
.B2(n_139),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_265),
.B(n_228),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_267),
.A2(n_194),
.B(n_221),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_328),
.Y(n_357)
);

NAND2x1p5_ASAP7_75t_L g358 ( 
.A(n_275),
.B(n_213),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_168),
.B1(n_139),
.B2(n_239),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_324),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_289),
.B(n_218),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_286),
.B(n_218),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_233),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_213),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_308),
.B(n_234),
.Y(n_365)
);

INVx4_ASAP7_75t_SL g366 ( 
.A(n_275),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_289),
.B(n_220),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_303),
.B(n_224),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_252),
.B(n_242),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_291),
.B(n_305),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_305),
.B(n_229),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_271),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_310),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_295),
.A2(n_297),
.B1(n_306),
.B2(n_304),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_272),
.B(n_165),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_276),
.B(n_192),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_303),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_276),
.B(n_192),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_311),
.B(n_246),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_277),
.B(n_192),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_297),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_306),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_272),
.B(n_288),
.Y(n_386)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_293),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_313),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_263),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_271),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_309),
.B(n_180),
.Y(n_392)
);

AO22x2_ASAP7_75t_L g393 ( 
.A1(n_312),
.A2(n_211),
.B1(n_180),
.B2(n_188),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_282),
.B(n_180),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_258),
.B(n_201),
.Y(n_395)
);

OR2x2_ASAP7_75t_SL g396 ( 
.A(n_317),
.B(n_247),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_317),
.Y(n_399)
);

AO22x2_ASAP7_75t_L g400 ( 
.A1(n_319),
.A2(n_247),
.B1(n_204),
.B2(n_163),
.Y(n_400)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_251),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_267),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_300),
.C(n_294),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_339),
.B(n_296),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_296),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_334),
.A2(n_281),
.B(n_288),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_375),
.A2(n_327),
.B1(n_317),
.B2(n_163),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_356),
.A2(n_194),
.B(n_223),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_375),
.A2(n_327),
.B1(n_254),
.B2(n_279),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_369),
.A2(n_279),
.B(n_253),
.Y(n_411)
);

CKINVDCx10_ASAP7_75t_R g412 ( 
.A(n_341),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_358),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_271),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_346),
.B(n_285),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_384),
.A2(n_254),
.B(n_249),
.C(n_259),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_266),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_366),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_336),
.A2(n_255),
.B(n_262),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_284),
.Y(n_421)
);

BUFx4f_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_35),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_262),
.B1(n_261),
.B2(n_260),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_372),
.B(n_255),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_301),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_377),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_386),
.A2(n_261),
.B(n_194),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_345),
.A2(n_202),
.B1(n_301),
.B2(n_223),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_347),
.A2(n_221),
.B1(n_223),
.B2(n_194),
.Y(n_431)
);

OR2x6_ASAP7_75t_SL g432 ( 
.A(n_357),
.B(n_202),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_358),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

AO21x1_ASAP7_75t_L g435 ( 
.A1(n_376),
.A2(n_290),
.B(n_268),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_345),
.A2(n_202),
.B1(n_223),
.B2(n_221),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_387),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_348),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_362),
.B(n_345),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_360),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_348),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_373),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_347),
.A2(n_348),
.B1(n_342),
.B2(n_352),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_338),
.A2(n_278),
.B(n_269),
.Y(n_446)
);

NOR2x1_ASAP7_75t_L g447 ( 
.A(n_368),
.B(n_273),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_400),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_367),
.A2(n_210),
.B(n_206),
.C(n_200),
.Y(n_450)
);

OA22x2_ASAP7_75t_L g451 ( 
.A1(n_396),
.A2(n_331),
.B1(n_330),
.B2(n_326),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_393),
.A2(n_201),
.B1(n_206),
.B2(n_210),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_365),
.B(n_58),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_392),
.A2(n_298),
.B(n_302),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_379),
.B(n_383),
.Y(n_457)
);

AO31x2_ASAP7_75t_L g458 ( 
.A1(n_431),
.A2(n_382),
.A3(n_398),
.B(n_397),
.Y(n_458)
);

BUFx12f_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_393),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_431),
.A2(n_394),
.B(n_361),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_426),
.B(n_387),
.Y(n_462)
);

AO22x2_ASAP7_75t_L g463 ( 
.A1(n_452),
.A2(n_400),
.B1(n_381),
.B2(n_335),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_422),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_406),
.A2(n_394),
.B(n_343),
.Y(n_465)
);

AO31x2_ASAP7_75t_L g466 ( 
.A1(n_452),
.A2(n_325),
.A3(n_331),
.B(n_330),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_432),
.Y(n_467)
);

NAND3xp33_ASAP7_75t_SL g468 ( 
.A(n_448),
.B(n_400),
.C(n_332),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_408),
.B(n_395),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_332),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_414),
.Y(n_471)
);

AO31x2_ASAP7_75t_L g472 ( 
.A1(n_445),
.A2(n_322),
.A3(n_314),
.B(n_315),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_425),
.A2(n_388),
.B1(n_370),
.B2(n_390),
.Y(n_473)
);

AOI211x1_ASAP7_75t_L g474 ( 
.A1(n_445),
.A2(n_206),
.B(n_200),
.C(n_74),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_354),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_407),
.A2(n_403),
.B1(n_427),
.B2(n_451),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_439),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_453),
.A2(n_424),
.B(n_410),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_449),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_422),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_440),
.B(n_443),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_407),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_415),
.A2(n_405),
.B(n_411),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_404),
.B(n_340),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_416),
.B(n_337),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_456),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_425),
.B(n_200),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_430),
.A2(n_200),
.B(n_326),
.C(n_316),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_428),
.B(n_70),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_421),
.B(n_72),
.Y(n_491)
);

AO31x2_ASAP7_75t_L g492 ( 
.A1(n_450),
.A2(n_316),
.A3(n_323),
.B(n_322),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_436),
.Y(n_493)
);

AND3x4_ASAP7_75t_L g494 ( 
.A(n_401),
.B(n_78),
.C(n_84),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_87),
.Y(n_495)
);

AOI211x1_ASAP7_75t_L g496 ( 
.A1(n_410),
.A2(n_97),
.B(n_321),
.C(n_316),
.Y(n_496)
);

NAND2x1p5_ASAP7_75t_L g497 ( 
.A(n_419),
.B(n_320),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_447),
.Y(n_498)
);

CKINVDCx8_ASAP7_75t_R g499 ( 
.A(n_414),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_433),
.B(n_270),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_433),
.Y(n_501)
);

CKINVDCx6p67_ASAP7_75t_R g502 ( 
.A(n_433),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_438),
.B(n_442),
.Y(n_503)
);

AO31x2_ASAP7_75t_L g504 ( 
.A1(n_417),
.A2(n_420),
.A3(n_446),
.B(n_455),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_454),
.B(n_434),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_423),
.A2(n_444),
.B1(n_454),
.B2(n_434),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_402),
.B(n_339),
.Y(n_507)
);

AO31x2_ASAP7_75t_L g508 ( 
.A1(n_431),
.A2(n_452),
.A3(n_445),
.B(n_435),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_402),
.B(n_339),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_402),
.A2(n_389),
.B1(n_425),
.B2(n_287),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_448),
.A2(n_407),
.B1(n_426),
.B2(n_287),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_402),
.B(n_339),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_419),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_402),
.B(n_339),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_409),
.A2(n_356),
.B(n_437),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_SL g517 ( 
.A1(n_453),
.A2(n_421),
.B(n_365),
.C(n_437),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_402),
.B(n_339),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_426),
.B(n_355),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_402),
.B(n_339),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_482),
.B(n_462),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g523 ( 
.A(n_459),
.B(n_477),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_507),
.B(n_509),
.Y(n_524)
);

OAI222xp33_ASAP7_75t_L g525 ( 
.A1(n_512),
.A2(n_476),
.B1(n_467),
.B2(n_510),
.C1(n_511),
.C2(n_460),
.Y(n_525)
);

AOI332xp33_ASAP7_75t_L g526 ( 
.A1(n_519),
.A2(n_476),
.A3(n_521),
.B1(n_518),
.B2(n_515),
.B3(n_513),
.C1(n_511),
.C2(n_481),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_479),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

O2A1O1Ixp33_ASAP7_75t_SL g529 ( 
.A1(n_517),
.A2(n_491),
.B(n_470),
.C(n_488),
.Y(n_529)
);

OAI22xp33_ASAP7_75t_L g530 ( 
.A1(n_467),
.A2(n_468),
.B1(n_490),
.B2(n_503),
.Y(n_530)
);

INVx4_ASAP7_75t_SL g531 ( 
.A(n_471),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_463),
.A2(n_494),
.B1(n_481),
.B2(n_520),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_463),
.A2(n_495),
.B1(n_506),
.B2(n_514),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_489),
.A2(n_464),
.B1(n_480),
.B2(n_469),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_493),
.B(n_475),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_499),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_478),
.B(n_471),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_502),
.B(n_485),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_474),
.A2(n_461),
.B1(n_496),
.B2(n_484),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_501),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_483),
.B(n_461),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_457),
.A2(n_465),
.B(n_473),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_458),
.B(n_508),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_501),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_458),
.B(n_508),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_498),
.B(n_514),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_505),
.B(n_471),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_514),
.Y(n_549)
);

CKINVDCx6p67_ASAP7_75t_R g550 ( 
.A(n_487),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_516),
.Y(n_551)
);

OR2x4_ASAP7_75t_L g552 ( 
.A(n_474),
.B(n_496),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_500),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_497),
.Y(n_554)
);

AO21x2_ASAP7_75t_L g555 ( 
.A1(n_458),
.A2(n_508),
.B(n_472),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_472),
.A2(n_466),
.B(n_492),
.Y(n_556)
);

O2A1O1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_472),
.A2(n_504),
.B(n_466),
.C(n_492),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_479),
.Y(n_558)
);

AND2x2_ASAP7_75t_SL g559 ( 
.A(n_467),
.B(n_512),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_459),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_459),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_464),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_479),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g564 ( 
.A1(n_482),
.A2(n_287),
.B1(n_353),
.B2(n_467),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_514),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_511),
.B(n_507),
.Y(n_566)
);

AOI221xp5_ASAP7_75t_L g567 ( 
.A1(n_512),
.A2(n_407),
.B1(n_333),
.B2(n_400),
.C(n_345),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_499),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_524),
.B(n_566),
.Y(n_569)
);

INVx4_ASAP7_75t_SL g570 ( 
.A(n_537),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_566),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_553),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_555),
.B(n_546),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_544),
.B(n_546),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_552),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_552),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_550),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_544),
.B(n_542),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_555),
.B(n_559),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_531),
.Y(n_581)
);

AOI222xp33_ASAP7_75t_L g582 ( 
.A1(n_567),
.A2(n_564),
.B1(n_525),
.B2(n_522),
.C1(n_532),
.C2(n_560),
.Y(n_582)
);

AOI21xp33_ASAP7_75t_L g583 ( 
.A1(n_530),
.A2(n_542),
.B(n_540),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_531),
.B(n_543),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_556),
.B(n_558),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_549),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_556),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_533),
.B(n_563),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_573),
.B(n_551),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_573),
.B(n_533),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_574),
.B(n_549),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_587),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_570),
.B(n_531),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_569),
.B(n_567),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_569),
.B(n_564),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_585),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_584),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_585),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_574),
.B(n_548),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_575),
.B(n_557),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_578),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_586),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_602),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_596),
.B(n_580),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_596),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_592),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_598),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_580),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_601),
.B(n_571),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_591),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_591),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_592),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_610),
.B(n_600),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_603),
.B(n_599),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_589),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_612),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_605),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_605),
.Y(n_618)
);

NAND2x1p5_ASAP7_75t_L g619 ( 
.A(n_607),
.B(n_577),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_606),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_600),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_616),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_614),
.B(n_604),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_616),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_620),
.Y(n_625)
);

NAND4xp25_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_582),
.C(n_595),
.D(n_577),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_619),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_617),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_615),
.B(n_608),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_615),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_628),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_622),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_626),
.A2(n_582),
.B1(n_621),
.B2(n_590),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_628),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_627),
.A2(n_590),
.B1(n_607),
.B2(n_608),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_623),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_624),
.Y(n_637)
);

AOI322xp5_ASAP7_75t_L g638 ( 
.A1(n_633),
.A2(n_580),
.A3(n_594),
.B1(n_607),
.B2(n_530),
.C1(n_588),
.C2(n_618),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_630),
.B(n_625),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_631),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_637),
.Y(n_641)
);

OAI21xp33_ASAP7_75t_L g642 ( 
.A1(n_638),
.A2(n_635),
.B(n_634),
.Y(n_642)
);

AOI211xp5_ASAP7_75t_L g643 ( 
.A1(n_641),
.A2(n_523),
.B(n_525),
.C(n_577),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_L g644 ( 
.A1(n_640),
.A2(n_636),
.B(n_630),
.Y(n_644)
);

AOI211xp5_ASAP7_75t_L g645 ( 
.A1(n_643),
.A2(n_577),
.B(n_583),
.C(n_593),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_642),
.A2(n_639),
.B(n_561),
.Y(n_646)
);

OAI211xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_644),
.B(n_526),
.C(n_545),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_645),
.B(n_536),
.C(n_565),
.Y(n_648)
);

NOR3xp33_ASAP7_75t_L g649 ( 
.A(n_647),
.B(n_536),
.C(n_565),
.Y(n_649)
);

AND3x4_ASAP7_75t_L g650 ( 
.A(n_648),
.B(n_593),
.C(n_632),
.Y(n_650)
);

NOR2x1_ASAP7_75t_L g651 ( 
.A(n_650),
.B(n_541),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_649),
.Y(n_652)
);

XNOR2x1_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_568),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_651),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_652),
.B(n_632),
.Y(n_655)
);

XOR2x2_ASAP7_75t_L g656 ( 
.A(n_653),
.B(n_619),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_655),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_655),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_SL g659 ( 
.A1(n_654),
.A2(n_568),
.B1(n_581),
.B2(n_538),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_654),
.A2(n_568),
.B1(n_576),
.B2(n_572),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_654),
.A2(n_539),
.B1(n_593),
.B2(n_534),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_657),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_658),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_656),
.A2(n_554),
.B(n_538),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_659),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_661),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_660),
.B(n_547),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_659),
.A2(n_593),
.B1(n_562),
.B2(n_581),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_657),
.A2(n_554),
.B(n_581),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_662),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_663),
.A2(n_666),
.B1(n_665),
.B2(n_667),
.Y(n_671)
);

AOI22x1_ASAP7_75t_L g672 ( 
.A1(n_664),
.A2(n_562),
.B1(n_586),
.B2(n_528),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_670),
.A2(n_669),
.B1(n_668),
.B2(n_576),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_671),
.A2(n_527),
.B(n_529),
.Y(n_674)
);

AOI21xp33_ASAP7_75t_L g675 ( 
.A1(n_673),
.A2(n_672),
.B(n_569),
.Y(n_675)
);

AO21x2_ASAP7_75t_L g676 ( 
.A1(n_675),
.A2(n_674),
.B(n_609),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_676),
.A2(n_572),
.B1(n_588),
.B2(n_579),
.Y(n_677)
);


endmodule