module fake_netlist_6_2087_n_1902 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1902);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1902;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_67),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_136),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_75),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_179),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_73),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_71),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_30),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_68),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_17),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_86),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_106),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_46),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_74),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_42),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_105),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_124),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_90),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_89),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_137),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_92),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_88),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_116),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_114),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_38),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_112),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_26),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_160),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_32),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_109),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_175),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_194),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_36),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_122),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_78),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_165),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_172),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_135),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_56),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_168),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_91),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_127),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_164),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_33),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_24),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_2),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_50),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_61),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_178),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_6),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_66),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_44),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_0),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_158),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_40),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_5),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_144),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_40),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_22),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_95),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_133),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_103),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_93),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_7),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_2),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_48),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_181),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_101),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_182),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_79),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_49),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_150),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_87),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_156),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_64),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_142),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_54),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_147),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_162),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_188),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_50),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_12),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_65),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_3),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_154),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_83),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_119),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_41),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_189),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_32),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_29),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_36),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_123),
.Y(n_314)
);

BUFx8_ASAP7_75t_SL g315 ( 
.A(n_81),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_102),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_155),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_47),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_184),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_121),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_34),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_113),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_18),
.Y(n_324)
);

BUFx8_ASAP7_75t_SL g325 ( 
.A(n_59),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_190),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_23),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_125),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_104),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_38),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_45),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_55),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_80),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_58),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_12),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_41),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_31),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_25),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_99),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_131),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_51),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_117),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_35),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_22),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_39),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_49),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_118),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_187),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_58),
.Y(n_349)
);

BUFx10_ASAP7_75t_L g350 ( 
.A(n_77),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_52),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_33),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_24),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_39),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_44),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_76),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_23),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_193),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_1),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_176),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_134),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_3),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_140),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_130),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_43),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_143),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_43),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_152),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_37),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_14),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_10),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_96),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_20),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_185),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_31),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_16),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_195),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_151),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_26),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_53),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_47),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_70),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_11),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_7),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_84),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_14),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_9),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_55),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_69),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_51),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_1),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_161),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_25),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_110),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_60),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_35),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_220),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_395),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_325),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_245),
.Y(n_402)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_303),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_269),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_239),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_199),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_241),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_370),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_246),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_247),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_253),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_390),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_345),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_199),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_236),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_260),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_261),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_268),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_263),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_296),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_282),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_264),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_274),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_276),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_277),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_291),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_226),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_305),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_312),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_337),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_299),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_270),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_341),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_344),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_282),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_286),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_378),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_271),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_286),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_300),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_226),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_382),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_300),
.Y(n_458)
);

BUFx2_ASAP7_75t_SL g459 ( 
.A(n_232),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_279),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_208),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_315),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_363),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_283),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_212),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_244),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_363),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_207),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_210),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_215),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_226),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_342),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_208),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_284),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_285),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_251),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_360),
.Y(n_478)
);

BUFx2_ASAP7_75t_SL g479 ( 
.A(n_232),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_214),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_228),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_214),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_297),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_216),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_231),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_206),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_206),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_225),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_218),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_217),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_222),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_298),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_223),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_302),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_229),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_230),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_219),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_225),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_415),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_415),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_290),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_371),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_440),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_456),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_472),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_469),
.B(n_290),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_422),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_397),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_459),
.B(n_371),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_419),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_401),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_440),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_481),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_403),
.A2(n_357),
.B1(n_211),
.B2(n_362),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_419),
.B(n_292),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_440),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_479),
.B(n_248),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_404),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_470),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_448),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_448),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_410),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_450),
.B(n_451),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_454),
.B(n_292),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_411),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_471),
.B(n_492),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_402),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_412),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_474),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_413),
.Y(n_547)
);

OA21x2_ASAP7_75t_L g548 ( 
.A1(n_487),
.A2(n_372),
.B(n_235),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_487),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_482),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_494),
.B(n_198),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_488),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_486),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_496),
.B(n_372),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_499),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_480),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_489),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_499),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_423),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_423),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_480),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_497),
.B(n_198),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_455),
.B(n_234),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_458),
.B(n_237),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_428),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_461),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_428),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_463),
.B(n_200),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_498),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_429),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_429),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_477),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_468),
.B(n_256),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_430),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_424),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_430),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_479),
.B(n_200),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_529),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_522),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_522),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_529),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_532),
.B(n_418),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_532),
.B(n_433),
.Y(n_587)
);

AOI21x1_ASAP7_75t_L g588 ( 
.A1(n_539),
.A2(n_275),
.B(n_272),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_522),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_510),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_534),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_557),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_503),
.B(n_466),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

BUFx8_ASAP7_75t_SL g595 ( 
.A(n_516),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_516),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_568),
.B(n_478),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_539),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_542),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_503),
.B(n_467),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_557),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_510),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_565),
.B(n_434),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_502),
.A2(n_398),
.B1(n_473),
.B2(n_484),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_523),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_581),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_510),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_510),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_542),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_523),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_530),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_502),
.B(n_406),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_520),
.B(n_490),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_563),
.Y(n_618)
);

INVx8_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_504),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_504),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_545),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_509),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_545),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_547),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_547),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_509),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_530),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_530),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_581),
.B(n_406),
.Y(n_631)
);

AO21x2_ASAP7_75t_L g632 ( 
.A1(n_571),
.A2(n_281),
.B(n_280),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_571),
.B(n_438),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_509),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_512),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_510),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_530),
.B(n_226),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_512),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_530),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_527),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_565),
.B(n_434),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_530),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_530),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_531),
.A2(n_313),
.B1(n_398),
.B2(n_309),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_565),
.B(n_425),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_527),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_531),
.B(n_425),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_535),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_566),
.B(n_427),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_568),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_535),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_566),
.B(n_427),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_580),
.Y(n_653)
);

AO21x2_ASAP7_75t_L g654 ( 
.A1(n_551),
.A2(n_294),
.B(n_288),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_512),
.Y(n_655)
);

AND3x1_ASAP7_75t_L g656 ( 
.A(n_526),
.B(n_407),
.C(n_465),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_520),
.B(n_409),
.Y(n_657)
);

AND3x2_ASAP7_75t_L g658 ( 
.A(n_563),
.B(n_332),
.C(n_250),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_572),
.B(n_420),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_517),
.Y(n_660)
);

INVx8_ASAP7_75t_L g661 ( 
.A(n_543),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_580),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_572),
.B(n_420),
.Y(n_663)
);

CKINVDCx16_ASAP7_75t_R g664 ( 
.A(n_544),
.Y(n_664)
);

NOR2x1p5_ASAP7_75t_L g665 ( 
.A(n_575),
.B(n_400),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_575),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_551),
.B(n_421),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_536),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_517),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_548),
.A2(n_307),
.B(n_295),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_535),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_535),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_533),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_533),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_505),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_564),
.B(n_421),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_517),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_518),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_518),
.Y(n_679)
);

INVxp33_ASAP7_75t_L g680 ( 
.A(n_505),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_519),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_519),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_521),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_566),
.B(n_465),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_546),
.B(n_432),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_533),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_511),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_511),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_564),
.B(n_432),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_500),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_543),
.B(n_435),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_521),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_543),
.B(n_435),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_543),
.B(n_445),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_500),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_501),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_543),
.B(n_445),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_536),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_576),
.B(n_226),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_501),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_580),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_506),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_546),
.B(n_453),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_576),
.B(n_453),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_536),
.B(n_460),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_506),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_550),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_550),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_536),
.B(n_460),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_511),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_576),
.B(n_464),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_526),
.A2(n_495),
.B1(n_493),
.B2(n_464),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_507),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_540),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_540),
.B(n_485),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_525),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_540),
.B(n_476),
.C(n_475),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_541),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_541),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_544),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_513),
.B(n_475),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_507),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_514),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_511),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_514),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_554),
.B(n_476),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_554),
.A2(n_439),
.B1(n_441),
.B2(n_449),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_515),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_515),
.Y(n_729)
);

BUFx6f_ASAP7_75t_SL g730 ( 
.A(n_554),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_580),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_650),
.B(n_483),
.Y(n_732)
);

INVx8_ASAP7_75t_L g733 ( 
.A(n_619),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_627),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_608),
.B(n_541),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_582),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_608),
.B(n_580),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_654),
.A2(n_548),
.B1(n_554),
.B2(n_266),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_667),
.A2(n_405),
.B1(n_452),
.B2(n_444),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_583),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_627),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_619),
.B(n_580),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_592),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_619),
.B(n_580),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_650),
.B(n_483),
.Y(n_745)
);

OAI22xp33_ASAP7_75t_L g746 ( 
.A1(n_718),
.A2(n_262),
.B1(n_327),
.B2(n_273),
.Y(n_746)
);

BUFx5_ASAP7_75t_L g747 ( 
.A(n_648),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_619),
.B(n_549),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_583),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_654),
.A2(n_548),
.B1(n_554),
.B2(n_379),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_657),
.B(n_493),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_631),
.B(n_721),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_654),
.A2(n_548),
.B1(n_353),
.B2(n_388),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_708),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_582),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_675),
.B(n_495),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_661),
.B(n_233),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_719),
.B(n_549),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_586),
.B(n_457),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_584),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_585),
.B(n_558),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_675),
.B(n_525),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_640),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_591),
.B(n_558),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_591),
.B(n_596),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_587),
.B(n_400),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_596),
.B(n_558),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_661),
.B(n_238),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_599),
.B(n_558),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_614),
.B(n_201),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_599),
.A2(n_513),
.B(n_358),
.C(n_310),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_705),
.B(n_201),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_668),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_704),
.B(n_202),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_600),
.B(n_558),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_600),
.B(n_569),
.Y(n_776)
);

INVx8_ASAP7_75t_L g777 ( 
.A(n_661),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_708),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_584),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_641),
.B(n_567),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_611),
.B(n_569),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_711),
.B(n_202),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_641),
.B(n_714),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_592),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_676),
.A2(n_348),
.B1(n_306),
.B2(n_293),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_717),
.B(n_553),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_L g787 ( 
.A(n_661),
.B(n_240),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_641),
.B(n_668),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_714),
.A2(n_391),
.B1(n_219),
.B2(n_384),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_663),
.B(n_462),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_606),
.B(n_553),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_646),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_611),
.B(n_569),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_SL g794 ( 
.A(n_716),
.B(n_218),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_622),
.B(n_624),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_622),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_616),
.B(n_203),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_624),
.B(n_569),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_625),
.B(n_569),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_625),
.Y(n_800)
);

AND2x6_ASAP7_75t_L g801 ( 
.A(n_648),
.B(n_287),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_632),
.A2(n_548),
.B1(n_289),
.B2(n_301),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_626),
.A2(n_314),
.B(n_326),
.C(n_347),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_689),
.B(n_203),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_605),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_626),
.B(n_690),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_690),
.B(n_569),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_569),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_699),
.A2(n_556),
.B(n_552),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_695),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_605),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_696),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_680),
.B(n_204),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_589),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_589),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_593),
.B(n_204),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_698),
.B(n_567),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_603),
.B(n_579),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_712),
.B(n_205),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_709),
.B(n_205),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_696),
.Y(n_821)
);

NOR3xp33_ASAP7_75t_L g822 ( 
.A(n_602),
.B(n_693),
.C(n_691),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_700),
.B(n_552),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_647),
.B(n_318),
.C(n_311),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_594),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_700),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_698),
.B(n_209),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_607),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_702),
.B(n_552),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_702),
.B(n_706),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_659),
.B(n_209),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_706),
.B(n_556),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_703),
.B(n_213),
.Y(n_833)
);

NAND2x1_ASAP7_75t_L g834 ( 
.A(n_604),
.B(n_508),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_713),
.B(n_556),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_713),
.B(n_508),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_726),
.B(n_213),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_728),
.B(n_651),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_633),
.A2(n_697),
.B1(n_694),
.B2(n_730),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_645),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_651),
.B(n_508),
.Y(n_841)
);

BUFx5_ASAP7_75t_L g842 ( 
.A(n_671),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_671),
.B(n_508),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_633),
.B(n_221),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_645),
.B(n_221),
.Y(n_845)
);

INVx8_ASAP7_75t_L g846 ( 
.A(n_730),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_649),
.B(n_224),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_672),
.B(n_555),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_633),
.B(n_224),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_649),
.B(n_570),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_652),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_652),
.B(n_227),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_633),
.A2(n_329),
.B1(n_242),
.B2(n_249),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_684),
.B(n_227),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_612),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_612),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_672),
.B(n_555),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_603),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_707),
.B(n_374),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_632),
.B(n_559),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_684),
.B(n_374),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_644),
.B(n_377),
.Y(n_862)
);

O2A1O1Ixp5_ASAP7_75t_L g863 ( 
.A1(n_670),
.A2(n_579),
.B(n_577),
.C(n_574),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_715),
.Y(n_864)
);

BUFx5_ASAP7_75t_L g865 ( 
.A(n_731),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_685),
.B(n_377),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_632),
.B(n_559),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_722),
.B(n_560),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_723),
.B(n_252),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_715),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_615),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_678),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_725),
.B(n_560),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_618),
.B(n_385),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_618),
.B(n_385),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_729),
.B(n_368),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_673),
.B(n_561),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_699),
.A2(n_562),
.B(n_561),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_615),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_647),
.B(n_389),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_673),
.B(n_561),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_715),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_715),
.A2(n_376),
.B1(n_367),
.B2(n_369),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_674),
.B(n_562),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_647),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_647),
.B(n_570),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_658),
.B(n_389),
.Y(n_887)
);

OR2x6_ASAP7_75t_SL g888 ( 
.A(n_824),
.B(n_716),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_736),
.B(n_674),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_734),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_739),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_741),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_747),
.B(n_731),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_736),
.B(n_686),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_752),
.B(n_598),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_755),
.B(n_686),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_755),
.B(n_604),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_753),
.A2(n_730),
.B1(n_692),
.B2(n_683),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_751),
.B(n_759),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_753),
.A2(n_738),
.B1(n_750),
.B2(n_851),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_747),
.B(n_842),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_742),
.A2(n_630),
.B(n_613),
.Y(n_902)
);

NOR2xp67_ASAP7_75t_L g903 ( 
.A(n_745),
.B(n_573),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_743),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_851),
.B(n_604),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_822),
.A2(n_656),
.B1(n_665),
.B2(n_639),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_777),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_732),
.B(n_666),
.Y(n_908)
);

O2A1O1Ixp5_ASAP7_75t_L g909 ( 
.A1(n_860),
.A2(n_588),
.B(n_670),
.C(n_678),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_735),
.B(n_609),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_788),
.B(n_665),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_747),
.B(n_613),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_796),
.B(n_609),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_800),
.B(n_609),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_810),
.B(n_617),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_738),
.A2(n_681),
.B1(n_692),
.B2(n_683),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_743),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_812),
.B(n_617),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_763),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_756),
.B(n_666),
.Y(n_920)
);

BUFx8_ASAP7_75t_L g921 ( 
.A(n_762),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_792),
.Y(n_922)
);

INVx3_ASAP7_75t_SL g923 ( 
.A(n_846),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_818),
.Y(n_924)
);

AND3x1_ASAP7_75t_L g925 ( 
.A(n_791),
.B(n_485),
.C(n_727),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_846),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_840),
.B(n_666),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_747),
.B(n_613),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_733),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_822),
.A2(n_642),
.B1(n_630),
.B2(n_639),
.Y(n_930)
);

BUFx4f_ASAP7_75t_L g931 ( 
.A(n_846),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_773),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_872),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_790),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_747),
.B(n_630),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_788),
.B(n_720),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_740),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_805),
.B(n_811),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_747),
.B(n_639),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_821),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_864),
.B(n_720),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_842),
.B(n_642),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_SL g943 ( 
.A(n_870),
.B(n_287),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_826),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_749),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_886),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_760),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_779),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_874),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_795),
.B(n_617),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_784),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_777),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_780),
.Y(n_953)
);

AND2x6_ASAP7_75t_SL g954 ( 
.A(n_887),
.B(n_442),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_842),
.B(n_642),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_784),
.B(n_597),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_780),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_814),
.Y(n_958)
);

AOI21xp33_ASAP7_75t_L g959 ( 
.A1(n_831),
.A2(n_322),
.B(n_320),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_858),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_882),
.B(n_885),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_773),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_806),
.B(n_636),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_850),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_783),
.A2(n_682),
.B1(n_679),
.B2(n_681),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_815),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_850),
.Y(n_967)
);

NOR2x2_ASAP7_75t_L g968 ( 
.A(n_746),
.B(n_664),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_838),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_817),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_817),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_825),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_875),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_765),
.B(n_724),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_830),
.B(n_724),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_845),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_733),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_847),
.Y(n_978)
);

CKINVDCx11_ASAP7_75t_R g979 ( 
.A(n_746),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_766),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_868),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_733),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_737),
.B(n_750),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_828),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_754),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_777),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_852),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_802),
.A2(n_867),
.B1(n_789),
.B2(n_883),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_837),
.A2(n_682),
.B1(n_679),
.B2(n_653),
.Y(n_989)
);

AO22x1_ASAP7_75t_L g990 ( 
.A1(n_833),
.A2(n_367),
.B1(n_369),
.B2(n_375),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_858),
.B(n_664),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_802),
.A2(n_287),
.B1(n_289),
.B2(n_301),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_873),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_SL g994 ( 
.A(n_819),
.B(n_287),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_758),
.B(n_710),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_855),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_834),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_SL g998 ( 
.A(n_789),
.B(n_376),
.C(n_375),
.Y(n_998)
);

OAI22xp33_ASAP7_75t_L g999 ( 
.A1(n_794),
.A2(n_380),
.B1(n_384),
.B2(n_387),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_839),
.A2(n_394),
.B1(n_688),
.B2(n_687),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_748),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_848),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_842),
.B(n_636),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_857),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_856),
.B(n_653),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_883),
.A2(n_287),
.B1(n_289),
.B2(n_301),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_744),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_871),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_842),
.B(n_590),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_754),
.B(n_573),
.Y(n_1010)
);

AND3x1_ASAP7_75t_L g1011 ( 
.A(n_844),
.B(n_446),
.C(n_443),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_862),
.A2(n_289),
.B1(n_301),
.B2(n_380),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_836),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_778),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_816),
.A2(n_289),
.B1(n_301),
.B2(n_393),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_769),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_842),
.B(n_710),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_772),
.B(n_636),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_865),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_778),
.B(n_574),
.Y(n_1020)
);

OAI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_853),
.A2(n_387),
.B1(n_393),
.B2(n_577),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_L g1022 ( 
.A(n_865),
.B(n_590),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_879),
.B(n_653),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_774),
.A2(n_637),
.B(n_638),
.C(n_628),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_823),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_797),
.B(n_687),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_775),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_865),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_865),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_829),
.A2(n_304),
.B1(n_243),
.B2(n_350),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_865),
.B(n_687),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_832),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_SL g1033 ( 
.A1(n_849),
.A2(n_218),
.B1(n_243),
.B2(n_304),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_835),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_865),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_863),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_761),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_764),
.B(n_688),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_786),
.B(n_447),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_813),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_770),
.B(n_662),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_801),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_L g1043 ( 
.A(n_866),
.B(n_662),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_863),
.A2(n_588),
.B(n_662),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_776),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_854),
.B(n_431),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_781),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_SL g1048 ( 
.A1(n_880),
.A2(n_338),
.B1(n_352),
.B2(n_324),
.Y(n_1048)
);

NOR2x1p5_ASAP7_75t_L g1049 ( 
.A(n_876),
.B(n_595),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_861),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_757),
.A2(n_787),
.B(n_768),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_801),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_767),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_827),
.B(n_820),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_793),
.B(n_701),
.Y(n_1055)
);

OAI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_859),
.A2(n_355),
.B(n_330),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_798),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_799),
.Y(n_1058)
);

NAND2x1p5_ASAP7_75t_L g1059 ( 
.A(n_807),
.B(n_701),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_808),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_841),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_843),
.B(n_877),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_782),
.B(n_436),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_881),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_899),
.B(n_804),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_899),
.A2(n_887),
.B(n_869),
.C(n_878),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_900),
.A2(n_785),
.B1(n_771),
.B2(n_809),
.Y(n_1067)
);

AO22x1_ASAP7_75t_L g1068 ( 
.A1(n_980),
.A2(n_336),
.B1(n_331),
.B2(n_334),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_904),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1040),
.B(n_884),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1019),
.A2(n_643),
.B(n_610),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_R g1072 ( 
.A(n_891),
.B(n_394),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_900),
.A2(n_878),
.B1(n_809),
.B2(n_803),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_949),
.B(n_436),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_917),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_909),
.A2(n_634),
.B(n_677),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_973),
.B(n_335),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_907),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1019),
.A2(n_643),
.B(n_590),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_969),
.B(n_620),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_926),
.Y(n_1081)
);

INVx5_ASAP7_75t_L g1082 ( 
.A(n_907),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_921),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_992),
.A2(n_801),
.B1(n_255),
.B2(n_257),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_890),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_1009),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_892),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_934),
.B(n_343),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1028),
.A2(n_643),
.B(n_590),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_981),
.B(n_620),
.Y(n_1090)
);

INVx5_ASAP7_75t_L g1091 ( 
.A(n_907),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_993),
.B(n_621),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_951),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1028),
.A2(n_643),
.B(n_601),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_926),
.B(n_437),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_932),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_908),
.B(n_437),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_919),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_907),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1025),
.B(n_623),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_952),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_946),
.B(n_911),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_920),
.B(n_537),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1032),
.B(n_623),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_937),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1022),
.A2(n_643),
.B(n_601),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1034),
.B(n_628),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_911),
.B(n_537),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_945),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1002),
.B(n_634),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_977),
.B(n_538),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_956),
.B(n_346),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1002),
.B(n_635),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1004),
.B(n_635),
.Y(n_1114)
);

O2A1O1Ixp5_ASAP7_75t_L g1115 ( 
.A1(n_994),
.A2(n_669),
.B(n_660),
.C(n_655),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_924),
.B(n_349),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_970),
.B(n_254),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_992),
.A2(n_590),
.B(n_601),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_L g1119 ( 
.A(n_1033),
.B(n_396),
.C(n_365),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_985),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1051),
.A2(n_601),
.B(n_610),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_970),
.B(n_258),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_901),
.A2(n_601),
.B(n_610),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_895),
.B(n_259),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_927),
.B(n_354),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_901),
.A2(n_610),
.B(n_629),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_956),
.B(n_359),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_951),
.B(n_265),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_960),
.B(n_267),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_947),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_912),
.A2(n_610),
.B(n_629),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_960),
.B(n_1014),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_948),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_895),
.A2(n_356),
.B(n_328),
.C(n_333),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_988),
.A2(n_1006),
.B1(n_898),
.B2(n_922),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_988),
.A2(n_1012),
.B1(n_979),
.B2(n_1021),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_SL g1137 ( 
.A1(n_1033),
.A2(n_278),
.B1(n_308),
.B2(n_316),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_952),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1012),
.A2(n_979),
.B1(n_1021),
.B2(n_1006),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_976),
.A2(n_366),
.B(n_364),
.C(n_340),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_958),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_1010),
.B(n_562),
.Y(n_1142)
);

CKINVDCx14_ASAP7_75t_R g1143 ( 
.A(n_991),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_983),
.A2(n_898),
.B1(n_889),
.B2(n_896),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_991),
.B(n_317),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_938),
.B(n_319),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_940),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_999),
.A2(n_669),
.B(n_660),
.C(n_655),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_978),
.B(n_321),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_987),
.A2(n_323),
.B(n_339),
.C(n_361),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1050),
.B(n_243),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_L g1152 ( 
.A1(n_994),
.A2(n_638),
.B(n_578),
.C(n_801),
.Y(n_1152)
);

AO22x1_ASAP7_75t_L g1153 ( 
.A1(n_921),
.A2(n_801),
.B1(n_392),
.B2(n_350),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_912),
.A2(n_629),
.B(n_528),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_966),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1056),
.B(n_304),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1041),
.A2(n_578),
.B(n_392),
.C(n_350),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_952),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_999),
.A2(n_578),
.B(n_392),
.C(n_8),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_938),
.B(n_629),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1020),
.B(n_4),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_925),
.A2(n_528),
.B1(n_524),
.B2(n_511),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_944),
.Y(n_1163)
);

CKINVDCx11_ASAP7_75t_R g1164 ( 
.A(n_954),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_928),
.A2(n_629),
.B(n_528),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_977),
.B(n_63),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1026),
.A2(n_629),
.B(n_528),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_998),
.A2(n_4),
.B(n_5),
.C(n_8),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1054),
.B(n_9),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_935),
.A2(n_528),
.B(n_524),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1027),
.B(n_10),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1054),
.B(n_11),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1015),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_903),
.B(n_528),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_971),
.B(n_13),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_935),
.A2(n_524),
.B(n_511),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1064),
.B(n_18),
.Y(n_1177)
);

AOI221x1_ASAP7_75t_L g1178 ( 
.A1(n_943),
.A2(n_524),
.B1(n_511),
.B2(n_21),
.C(n_27),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_964),
.B(n_98),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1053),
.B(n_19),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_941),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_952),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1041),
.A2(n_524),
.B(n_20),
.C(n_21),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1057),
.B(n_19),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_967),
.B(n_27),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_906),
.B(n_108),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_936),
.B(n_28),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_998),
.A2(n_28),
.B(n_29),
.C(n_37),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_972),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_894),
.A2(n_120),
.B1(n_196),
.B2(n_186),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1058),
.B(n_42),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1045),
.B(n_45),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_939),
.A2(n_115),
.B(n_177),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_SL g1194 ( 
.A1(n_1015),
.A2(n_100),
.B(n_174),
.C(n_171),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1030),
.A2(n_46),
.B(n_48),
.C(n_52),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_936),
.B(n_53),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1063),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_932),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_986),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1046),
.B(n_57),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1063),
.A2(n_59),
.B(n_60),
.C(n_62),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_986),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_941),
.Y(n_1203)
);

OA22x2_ASAP7_75t_L g1204 ( 
.A1(n_941),
.A2(n_72),
.B1(n_82),
.B2(n_94),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_953),
.B(n_126),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1047),
.B(n_128),
.Y(n_1206)
);

OA22x2_ASAP7_75t_L g1207 ( 
.A1(n_1046),
.A2(n_961),
.B1(n_957),
.B2(n_1039),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1061),
.B(n_197),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_942),
.A2(n_129),
.B(n_141),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_986),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1016),
.B(n_146),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1082),
.B(n_929),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1121),
.A2(n_1044),
.B(n_909),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1065),
.B(n_1013),
.Y(n_1214)
);

OAI22x1_ASAP7_75t_L g1215 ( 
.A1(n_1135),
.A2(n_968),
.B1(n_1039),
.B2(n_1049),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1069),
.B(n_961),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1069),
.B(n_961),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1087),
.Y(n_1218)
);

NOR2x1_ASAP7_75t_L g1219 ( 
.A(n_1211),
.B(n_929),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1097),
.B(n_1060),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1123),
.A2(n_902),
.B(n_995),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1074),
.B(n_1060),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1076),
.A2(n_1036),
.B(n_1062),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_1066),
.A2(n_1018),
.B(n_905),
.C(n_910),
.Y(n_1224)
);

AOI221x1_ASAP7_75t_L g1225 ( 
.A1(n_1183),
.A2(n_943),
.B1(n_1000),
.B2(n_1001),
.C(n_1007),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1167),
.A2(n_1144),
.B(n_1073),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1112),
.B(n_1127),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1075),
.B(n_990),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1170),
.A2(n_1038),
.B(n_1017),
.Y(n_1229)
);

CKINVDCx11_ASAP7_75t_R g1230 ( 
.A(n_1083),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1120),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1067),
.A2(n_1055),
.A3(n_975),
.B(n_950),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1086),
.A2(n_986),
.B(n_982),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1176),
.A2(n_1003),
.B(n_1031),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1136),
.B(n_1030),
.C(n_1048),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1093),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1103),
.B(n_1145),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1067),
.A2(n_974),
.A3(n_963),
.B(n_1035),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1070),
.B(n_1060),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1126),
.A2(n_1059),
.B(n_893),
.Y(n_1240)
);

BUFx10_ASAP7_75t_L g1241 ( 
.A(n_1088),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1125),
.B(n_1011),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1142),
.B(n_1060),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1131),
.A2(n_1059),
.B(n_893),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1139),
.A2(n_1016),
.B1(n_1037),
.B2(n_984),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1200),
.B(n_1116),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1077),
.B(n_888),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1102),
.B(n_1007),
.Y(n_1248)
);

AO21x2_ASAP7_75t_L g1249 ( 
.A1(n_1162),
.A2(n_1135),
.B(n_1186),
.Y(n_1249)
);

INVx5_ASAP7_75t_L g1250 ( 
.A(n_1099),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1161),
.B(n_1171),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1178),
.A2(n_1029),
.A3(n_897),
.B(n_918),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1115),
.A2(n_1024),
.B(n_989),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1154),
.A2(n_1005),
.B(n_1023),
.Y(n_1254)
);

NAND3xp33_ASAP7_75t_L g1255 ( 
.A(n_1119),
.B(n_965),
.C(n_916),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1165),
.A2(n_1079),
.B(n_1071),
.Y(n_1256)
);

O2A1O1Ixp5_ASAP7_75t_SL g1257 ( 
.A1(n_1173),
.A2(n_962),
.B(n_1042),
.C(n_955),
.Y(n_1257)
);

AOI221xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1173),
.A2(n_916),
.B1(n_915),
.B2(n_913),
.C(n_914),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1147),
.B(n_1037),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1089),
.A2(n_1005),
.B(n_1023),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1094),
.A2(n_955),
.B(n_1043),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1148),
.A2(n_930),
.B(n_933),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1163),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1157),
.A2(n_1052),
.A3(n_996),
.B(n_1008),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1084),
.A2(n_962),
.B1(n_1007),
.B2(n_931),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1106),
.A2(n_1042),
.B(n_1001),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1118),
.A2(n_1007),
.B(n_1001),
.Y(n_1267)
);

AOI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1174),
.A2(n_1001),
.B(n_1052),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1169),
.B(n_931),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1156),
.A2(n_968),
.A3(n_997),
.B(n_170),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1143),
.B(n_923),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1152),
.A2(n_997),
.B(n_166),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1172),
.B(n_997),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1137),
.A2(n_159),
.A3(n_1190),
.B1(n_1188),
.B2(n_1168),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1201),
.A2(n_1208),
.A3(n_1206),
.B(n_1184),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1110),
.A2(n_1114),
.B(n_1113),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1080),
.A2(n_1090),
.B(n_1092),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1082),
.B(n_1091),
.Y(n_1278)
);

AO21x1_ASAP7_75t_L g1279 ( 
.A1(n_1195),
.A2(n_1162),
.B(n_1180),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1082),
.B(n_1091),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1100),
.A2(n_1107),
.B(n_1104),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1203),
.Y(n_1282)
);

AOI221x1_ASAP7_75t_L g1283 ( 
.A1(n_1137),
.A2(n_1197),
.B1(n_1191),
.B2(n_1134),
.C(n_1192),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1098),
.Y(n_1284)
);

OAI22x1_ASAP7_75t_L g1285 ( 
.A1(n_1187),
.A2(n_1196),
.B1(n_1185),
.B2(n_1132),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1081),
.Y(n_1286)
);

NAND3xp33_ASAP7_75t_L g1287 ( 
.A(n_1159),
.B(n_1151),
.C(n_1072),
.Y(n_1287)
);

INVx4_ASAP7_75t_L g1288 ( 
.A(n_1091),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1128),
.B(n_1129),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1084),
.A2(n_1177),
.B(n_1124),
.C(n_1149),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1175),
.A2(n_1207),
.B1(n_1179),
.B2(n_1204),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1117),
.A2(n_1122),
.B(n_1194),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1140),
.A2(n_1150),
.A3(n_1109),
.B(n_1141),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1105),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1160),
.A2(n_1155),
.B(n_1189),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1096),
.A2(n_1198),
.B(n_1133),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1181),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1179),
.B(n_1130),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1210),
.A2(n_1198),
.B(n_1096),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1108),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1108),
.Y(n_1301)
);

O2A1O1Ixp5_ASAP7_75t_L g1302 ( 
.A1(n_1146),
.A2(n_1153),
.B(n_1111),
.C(n_1205),
.Y(n_1302)
);

AO21x2_ASAP7_75t_L g1303 ( 
.A1(n_1111),
.A2(n_1166),
.B(n_1210),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1068),
.B(n_1095),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1166),
.B(n_1095),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1210),
.A2(n_1078),
.B(n_1158),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1078),
.A2(n_1158),
.B(n_1138),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1138),
.A2(n_1099),
.B1(n_1101),
.B2(n_1182),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1101),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1095),
.B(n_1202),
.Y(n_1310)
);

AND2x6_ASAP7_75t_L g1311 ( 
.A(n_1182),
.B(n_1199),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1202),
.B(n_1199),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1164),
.A2(n_1028),
.B(n_1019),
.Y(n_1313)
);

CKINVDCx8_ASAP7_75t_R g1314 ( 
.A(n_1120),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1136),
.A2(n_899),
.B1(n_1065),
.B2(n_1139),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1121),
.A2(n_1123),
.B(n_1076),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1167),
.A2(n_1051),
.B(n_1121),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1065),
.B(n_899),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1065),
.B(n_899),
.Y(n_1319)
);

AO21x2_ASAP7_75t_L g1320 ( 
.A1(n_1167),
.A2(n_1051),
.B(n_1121),
.Y(n_1320)
);

OAI22x1_ASAP7_75t_L g1321 ( 
.A1(n_1065),
.A2(n_899),
.B1(n_980),
.B2(n_934),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1085),
.Y(n_1322)
);

BUFx8_ASAP7_75t_L g1323 ( 
.A(n_1083),
.Y(n_1323)
);

INVx5_ASAP7_75t_L g1324 ( 
.A(n_1099),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_SL g1325 ( 
.A1(n_1211),
.A2(n_1209),
.B(n_1193),
.Y(n_1325)
);

BUFx4_ASAP7_75t_SL g1326 ( 
.A(n_1081),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1078),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1121),
.A2(n_1123),
.B(n_1076),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1065),
.B(n_899),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1082),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1065),
.B(n_899),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1073),
.A2(n_899),
.B(n_1067),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1073),
.A2(n_899),
.B(n_1067),
.Y(n_1333)
);

AO21x2_ASAP7_75t_L g1334 ( 
.A1(n_1167),
.A2(n_1051),
.B(n_1121),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1065),
.A2(n_899),
.B(n_751),
.C(n_895),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1065),
.B(n_1040),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_SL g1337 ( 
.A1(n_1066),
.A2(n_1194),
.B(n_1183),
.C(n_1186),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1121),
.A2(n_1123),
.B(n_1076),
.Y(n_1338)
);

NAND2x1_ASAP7_75t_L g1339 ( 
.A(n_1078),
.B(n_1019),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1073),
.A2(n_899),
.B(n_1067),
.Y(n_1340)
);

NOR2xp67_ASAP7_75t_L g1341 ( 
.A(n_1082),
.B(n_608),
.Y(n_1341)
);

BUFx4_ASAP7_75t_SL g1342 ( 
.A(n_1081),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1073),
.A2(n_899),
.B(n_1067),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1073),
.A2(n_899),
.B(n_1067),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1065),
.B(n_899),
.Y(n_1345)
);

O2A1O1Ixp5_ASAP7_75t_SL g1346 ( 
.A1(n_1173),
.A2(n_752),
.B(n_959),
.C(n_1124),
.Y(n_1346)
);

NAND3x1_ASAP7_75t_L g1347 ( 
.A(n_1119),
.B(n_899),
.C(n_526),
.Y(n_1347)
);

NAND3x1_ASAP7_75t_L g1348 ( 
.A(n_1119),
.B(n_899),
.C(n_526),
.Y(n_1348)
);

NOR2x1_ASAP7_75t_SL g1349 ( 
.A(n_1082),
.B(n_907),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1065),
.A2(n_899),
.B(n_751),
.C(n_895),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1076),
.A2(n_1044),
.B(n_909),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1076),
.A2(n_1044),
.B(n_909),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1073),
.A2(n_899),
.B(n_1067),
.Y(n_1353)
);

AO31x2_ASAP7_75t_L g1354 ( 
.A1(n_1073),
.A2(n_1067),
.A3(n_1144),
.B(n_1178),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1065),
.A2(n_899),
.B(n_752),
.C(n_751),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1074),
.B(n_1097),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1074),
.B(n_1097),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1081),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1314),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1332),
.A2(n_1353),
.B(n_1343),
.C(n_1344),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1227),
.A2(n_1315),
.B1(n_1251),
.B2(n_1329),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1235),
.A2(n_1340),
.B1(n_1353),
.B2(n_1333),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1256),
.A2(n_1221),
.B(n_1254),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1356),
.B(n_1357),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1335),
.A2(n_1350),
.B(n_1355),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1246),
.B(n_1289),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1332),
.A2(n_1340),
.B(n_1333),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1230),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1343),
.A2(n_1344),
.B(n_1226),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1315),
.A2(n_1318),
.B(n_1319),
.C(n_1345),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1235),
.A2(n_1331),
.B1(n_1287),
.B2(n_1321),
.Y(n_1371)
);

AOI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1292),
.A2(n_1268),
.B(n_1225),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1214),
.B(n_1237),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1242),
.B(n_1222),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1213),
.A2(n_1328),
.B(n_1316),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1338),
.A2(n_1258),
.B(n_1253),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1336),
.B(n_1287),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1260),
.A2(n_1261),
.B(n_1244),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1234),
.A2(n_1229),
.B(n_1240),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1279),
.A2(n_1283),
.A3(n_1290),
.B(n_1281),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1267),
.A2(n_1296),
.B(n_1223),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1346),
.A2(n_1347),
.B(n_1348),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1272),
.A2(n_1262),
.B(n_1334),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1325),
.A2(n_1266),
.B(n_1276),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1262),
.A2(n_1257),
.B(n_1277),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1250),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1263),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1337),
.A2(n_1302),
.B(n_1220),
.C(n_1273),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1255),
.A2(n_1291),
.B(n_1258),
.C(n_1272),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1358),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1317),
.A2(n_1334),
.B(n_1320),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1259),
.B(n_1248),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1288),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1322),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1219),
.A2(n_1295),
.B(n_1352),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1285),
.A2(n_1215),
.B1(n_1247),
.B2(n_1255),
.C(n_1304),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1269),
.B(n_1236),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1326),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1351),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1291),
.A2(n_1245),
.B1(n_1228),
.B2(n_1305),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1300),
.B(n_1241),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1342),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1241),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1245),
.A2(n_1243),
.B1(n_1239),
.B2(n_1217),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1298),
.A2(n_1295),
.B(n_1224),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1284),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_SL g1407 ( 
.A1(n_1313),
.A2(n_1299),
.B(n_1265),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1311),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1311),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1216),
.B(n_1301),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1249),
.A2(n_1294),
.B1(n_1303),
.B2(n_1310),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1233),
.B(n_1280),
.Y(n_1412)
);

NAND2x1p5_ASAP7_75t_L g1413 ( 
.A(n_1250),
.B(n_1324),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1323),
.B(n_1297),
.C(n_1271),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1312),
.B(n_1309),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_L g1416 ( 
.A(n_1286),
.B(n_1308),
.C(n_1341),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1339),
.A2(n_1307),
.B(n_1306),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1293),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1250),
.B(n_1324),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1249),
.A2(n_1274),
.B1(n_1323),
.B2(n_1354),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1212),
.A2(n_1327),
.B(n_1278),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1317),
.A2(n_1320),
.B(n_1349),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1293),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1354),
.A2(n_1232),
.B(n_1238),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1232),
.A2(n_1238),
.B(n_1275),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1311),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1232),
.A2(n_1264),
.B(n_1274),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1274),
.A2(n_1288),
.B1(n_1330),
.B2(n_1311),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1275),
.A2(n_1252),
.B(n_1270),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1330),
.A2(n_899),
.B1(n_1227),
.B2(n_980),
.Y(n_1430)
);

OAI21xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1252),
.A2(n_992),
.B(n_900),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1252),
.A2(n_1333),
.B(n_1332),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1332),
.A2(n_1340),
.B(n_1333),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1434)
);

CKINVDCx8_ASAP7_75t_R g1435 ( 
.A(n_1231),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1358),
.Y(n_1436)
);

AND2x6_ASAP7_75t_SL g1437 ( 
.A(n_1271),
.B(n_1088),
.Y(n_1437)
);

AO32x2_ASAP7_75t_L g1438 ( 
.A1(n_1354),
.A2(n_1173),
.A3(n_1137),
.B1(n_1144),
.B2(n_1067),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1250),
.Y(n_1439)
);

AOI21xp33_ASAP7_75t_SL g1440 ( 
.A1(n_1227),
.A2(n_980),
.B(n_934),
.Y(n_1440)
);

AO31x2_ASAP7_75t_L g1441 ( 
.A1(n_1225),
.A2(n_1279),
.A3(n_1178),
.B(n_1283),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1235),
.A2(n_899),
.B1(n_1315),
.B2(n_1227),
.Y(n_1443)
);

O2A1O1Ixp33_ASAP7_75t_L g1444 ( 
.A1(n_1335),
.A2(n_1350),
.B(n_899),
.C(n_1355),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1231),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1282),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1332),
.A2(n_1340),
.B(n_1333),
.Y(n_1447)
);

AO31x2_ASAP7_75t_L g1448 ( 
.A1(n_1225),
.A2(n_1279),
.A3(n_1178),
.B(n_1283),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1256),
.A2(n_1221),
.B(n_1254),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1235),
.A2(n_899),
.B1(n_1315),
.B2(n_1227),
.Y(n_1450)
);

BUFx4f_ASAP7_75t_L g1451 ( 
.A(n_1278),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1288),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1227),
.A2(n_899),
.B1(n_980),
.B2(n_1315),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1326),
.Y(n_1454)
);

AO31x2_ASAP7_75t_L g1455 ( 
.A1(n_1225),
.A2(n_1279),
.A3(n_1178),
.B(n_1283),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1332),
.A2(n_1340),
.B(n_1333),
.Y(n_1456)
);

OAI222xp33_ASAP7_75t_L g1457 ( 
.A1(n_1315),
.A2(n_1136),
.B1(n_1139),
.B2(n_1173),
.C1(n_900),
.C2(n_1227),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1332),
.A2(n_1340),
.B(n_1333),
.Y(n_1458)
);

AO22x1_ASAP7_75t_L g1459 ( 
.A1(n_1227),
.A2(n_899),
.B1(n_980),
.B2(n_934),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1315),
.A2(n_1227),
.B1(n_1319),
.B2(n_1318),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1288),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1282),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1256),
.A2(n_1221),
.B(n_1254),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1358),
.Y(n_1465)
);

CKINVDCx12_ASAP7_75t_R g1466 ( 
.A(n_1271),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1218),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1335),
.A2(n_1350),
.B(n_899),
.C(n_1355),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1218),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_SL g1470 ( 
.A1(n_1335),
.A2(n_1350),
.B(n_1290),
.C(n_1333),
.Y(n_1470)
);

NAND2x1p5_ASAP7_75t_L g1471 ( 
.A(n_1250),
.B(n_1082),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1356),
.B(n_1357),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1218),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1218),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1256),
.A2(n_1221),
.B(n_1254),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1356),
.B(n_1357),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1256),
.A2(n_1221),
.B(n_1254),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1335),
.A2(n_899),
.B1(n_1350),
.B2(n_1227),
.C(n_1319),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1358),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_SL g1480 ( 
.A1(n_1335),
.A2(n_1350),
.B(n_1290),
.C(n_1333),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1227),
.A2(n_899),
.B1(n_980),
.B2(n_934),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1227),
.A2(n_899),
.B(n_1335),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1332),
.A2(n_899),
.B(n_1340),
.C(n_1333),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_SL g1484 ( 
.A(n_1314),
.B(n_716),
.Y(n_1484)
);

BUFx2_ASAP7_75t_SL g1485 ( 
.A(n_1314),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1453),
.A2(n_1482),
.B(n_1468),
.C(n_1444),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1483),
.A2(n_1444),
.B(n_1468),
.C(n_1360),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_SL g1488 ( 
.A(n_1412),
.B(n_1409),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1390),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1359),
.Y(n_1490)
);

NOR4xp25_ASAP7_75t_L g1491 ( 
.A(n_1470),
.B(n_1480),
.C(n_1450),
.D(n_1443),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1483),
.A2(n_1360),
.B(n_1470),
.Y(n_1492)
);

O2A1O1Ixp5_ASAP7_75t_L g1493 ( 
.A1(n_1382),
.A2(n_1365),
.B(n_1459),
.C(n_1389),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1373),
.B(n_1392),
.Y(n_1494)
);

BUFx4f_ASAP7_75t_L g1495 ( 
.A(n_1368),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1362),
.B(n_1461),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1377),
.B(n_1371),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1410),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1397),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1478),
.A2(n_1377),
.B(n_1450),
.C(n_1443),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1481),
.B(n_1430),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1362),
.B(n_1461),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1445),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1371),
.B(n_1410),
.Y(n_1504)
);

O2A1O1Ixp5_ASAP7_75t_L g1505 ( 
.A1(n_1389),
.A2(n_1457),
.B(n_1405),
.C(n_1400),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1415),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1370),
.B(n_1361),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1420),
.A2(n_1434),
.B1(n_1460),
.B2(n_1442),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1446),
.B(n_1463),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1420),
.A2(n_1456),
.B1(n_1458),
.B2(n_1433),
.Y(n_1510)
);

O2A1O1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1457),
.A2(n_1480),
.B(n_1440),
.C(n_1396),
.Y(n_1511)
);

AOI211xp5_ASAP7_75t_L g1512 ( 
.A1(n_1400),
.A2(n_1404),
.B(n_1388),
.C(n_1401),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1466),
.A2(n_1435),
.B1(n_1414),
.B2(n_1485),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1422),
.A2(n_1379),
.B(n_1384),
.Y(n_1514)
);

INVx3_ASAP7_75t_SL g1515 ( 
.A(n_1398),
.Y(n_1515)
);

O2A1O1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1404),
.A2(n_1407),
.B(n_1431),
.C(n_1416),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1394),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1395),
.A2(n_1423),
.B(n_1381),
.Y(n_1518)
);

NOR2xp67_ASAP7_75t_L g1519 ( 
.A(n_1467),
.B(n_1469),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_SL g1520 ( 
.A1(n_1412),
.A2(n_1419),
.B(n_1413),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1367),
.B(n_1447),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1363),
.A2(n_1449),
.B(n_1477),
.Y(n_1522)
);

AOI221x1_ASAP7_75t_SL g1523 ( 
.A1(n_1473),
.A2(n_1474),
.B1(n_1406),
.B2(n_1426),
.C(n_1437),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1433),
.A2(n_1458),
.B1(n_1456),
.B2(n_1428),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1456),
.A2(n_1458),
.B1(n_1428),
.B2(n_1409),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1409),
.A2(n_1432),
.B1(n_1451),
.B2(n_1408),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1416),
.A2(n_1451),
.B(n_1411),
.C(n_1408),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1471),
.A2(n_1386),
.B(n_1439),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1432),
.B(n_1380),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1432),
.B(n_1380),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1380),
.B(n_1369),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1484),
.B(n_1479),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1403),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1380),
.B(n_1369),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1441),
.B(n_1455),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1411),
.A2(n_1454),
.B(n_1465),
.C(n_1436),
.Y(n_1536)
);

CKINVDCx16_ASAP7_75t_R g1537 ( 
.A(n_1436),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1409),
.A2(n_1427),
.B1(n_1438),
.B2(n_1386),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_SL g1539 ( 
.A(n_1383),
.B(n_1372),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1427),
.A2(n_1438),
.B1(n_1386),
.B2(n_1465),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1441),
.B(n_1448),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1448),
.B(n_1455),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1376),
.B(n_1479),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1421),
.A2(n_1462),
.B(n_1452),
.C(n_1393),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1402),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1427),
.A2(n_1439),
.B1(n_1376),
.B2(n_1399),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1376),
.A2(n_1399),
.B1(n_1424),
.B2(n_1418),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1424),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1464),
.A2(n_1475),
.B(n_1417),
.C(n_1378),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1383),
.B(n_1391),
.Y(n_1550)
);

INVxp67_ASAP7_75t_L g1551 ( 
.A(n_1391),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1375),
.A2(n_1483),
.B(n_1333),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1375),
.A2(n_1483),
.B(n_1333),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1375),
.A2(n_899),
.B(n_1350),
.C(n_1335),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1483),
.A2(n_1333),
.B(n_1332),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1385),
.A2(n_1425),
.B(n_1429),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1482),
.A2(n_1335),
.B(n_1350),
.C(n_899),
.Y(n_1557)
);

O2A1O1Ixp5_ASAP7_75t_L g1558 ( 
.A1(n_1382),
.A2(n_899),
.B(n_1333),
.C(n_1332),
.Y(n_1558)
);

AOI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1457),
.A2(n_899),
.B1(n_1480),
.B2(n_1470),
.C(n_1350),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1483),
.A2(n_1333),
.B(n_1332),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1360),
.A2(n_900),
.B1(n_992),
.B2(n_1006),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1385),
.A2(n_1425),
.B(n_1429),
.Y(n_1562)
);

O2A1O1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1453),
.A2(n_899),
.B(n_1350),
.C(n_1335),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1374),
.B(n_1364),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1374),
.B(n_1364),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1483),
.A2(n_1333),
.B(n_1332),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1483),
.A2(n_1333),
.B(n_1332),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1387),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1483),
.A2(n_899),
.B(n_1227),
.C(n_1355),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1362),
.B(n_1461),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1366),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1472),
.B(n_1476),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1453),
.A2(n_899),
.B(n_1350),
.C(n_1335),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1410),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1360),
.A2(n_900),
.B1(n_992),
.B2(n_1006),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1453),
.A2(n_899),
.B(n_1350),
.C(n_1335),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1483),
.A2(n_1333),
.B(n_1332),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1548),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1524),
.B(n_1550),
.Y(n_1579)
);

OR2x6_ASAP7_75t_L g1580 ( 
.A(n_1552),
.B(n_1553),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1498),
.Y(n_1581)
);

OR2x6_ASAP7_75t_L g1582 ( 
.A(n_1555),
.B(n_1560),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1518),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1524),
.B(n_1521),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1534),
.B(n_1531),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1551),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1531),
.B(n_1529),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1556),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1574),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1530),
.B(n_1541),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1510),
.B(n_1542),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1510),
.B(n_1535),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1497),
.B(n_1566),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1549),
.B(n_1488),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1562),
.Y(n_1597)
);

INVx3_ASAP7_75t_SL g1598 ( 
.A(n_1537),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1517),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1568),
.B(n_1539),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1540),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1540),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_L g1603 ( 
.A(n_1501),
.B(n_1500),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1514),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1525),
.B(n_1538),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1514),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1522),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1559),
.A2(n_1502),
.B1(n_1570),
.B2(n_1496),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1538),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1547),
.Y(n_1610)
);

BUFx4f_ASAP7_75t_SL g1611 ( 
.A(n_1515),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1546),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1566),
.A2(n_1577),
.B(n_1567),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1567),
.B(n_1577),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1525),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1507),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1519),
.Y(n_1617)
);

NOR3xp33_ASAP7_75t_L g1618 ( 
.A(n_1563),
.B(n_1576),
.C(n_1573),
.Y(n_1618)
);

AO21x2_ASAP7_75t_L g1619 ( 
.A1(n_1487),
.A2(n_1508),
.B(n_1492),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1558),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1526),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1607),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1579),
.B(n_1605),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1586),
.B(n_1508),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1595),
.B(n_1506),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1578),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1578),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1586),
.B(n_1601),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1588),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1579),
.B(n_1526),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1595),
.B(n_1496),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1596),
.B(n_1544),
.Y(n_1632)
);

BUFx8_ASAP7_75t_L g1633 ( 
.A(n_1621),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1579),
.B(n_1493),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1587),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1619),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1601),
.B(n_1499),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1585),
.B(n_1486),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1596),
.B(n_1600),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1584),
.B(n_1565),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1603),
.A2(n_1559),
.B1(n_1504),
.B2(n_1575),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1584),
.B(n_1564),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1583),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1582),
.B(n_1516),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1582),
.B(n_1491),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1583),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1582),
.B(n_1505),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1647),
.A2(n_1603),
.B(n_1619),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1643),
.A2(n_1618),
.B1(n_1619),
.B2(n_1647),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1623),
.B(n_1621),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1623),
.B(n_1635),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1626),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1643),
.A2(n_1618),
.B1(n_1523),
.B2(n_1608),
.C(n_1614),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1626),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1628),
.B(n_1593),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1647),
.A2(n_1619),
.B1(n_1580),
.B2(n_1582),
.Y(n_1658)
);

NOR4xp25_ASAP7_75t_SL g1659 ( 
.A(n_1629),
.B(n_1621),
.C(n_1533),
.D(n_1617),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1625),
.B(n_1598),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_L g1661 ( 
.A1(n_1639),
.A2(n_1511),
.B(n_1608),
.C(n_1512),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1636),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1622),
.A2(n_1597),
.B(n_1590),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1624),
.A2(n_1580),
.B1(n_1569),
.B2(n_1527),
.Y(n_1664)
);

AOI33xp33_ASAP7_75t_L g1665 ( 
.A1(n_1634),
.A2(n_1581),
.A3(n_1591),
.B1(n_1571),
.B2(n_1594),
.B3(n_1620),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1646),
.A2(n_1619),
.B1(n_1580),
.B2(n_1582),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1626),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_SL g1668 ( 
.A1(n_1624),
.A2(n_1557),
.B1(n_1580),
.B2(n_1615),
.C(n_1536),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1640),
.B(n_1596),
.Y(n_1669)
);

AOI222xp33_ASAP7_75t_L g1670 ( 
.A1(n_1639),
.A2(n_1615),
.B1(n_1609),
.B2(n_1561),
.C1(n_1620),
.C2(n_1513),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1625),
.B(n_1631),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1633),
.A2(n_1580),
.B1(n_1613),
.B2(n_1616),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1636),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1637),
.B(n_1616),
.C(n_1557),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1638),
.Y(n_1676)
);

BUFx3_ASAP7_75t_L g1677 ( 
.A(n_1638),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1641),
.B(n_1581),
.Y(n_1678)
);

AOI222xp33_ASAP7_75t_L g1679 ( 
.A1(n_1634),
.A2(n_1609),
.B1(n_1561),
.B2(n_1620),
.C1(n_1616),
.C2(n_1594),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1638),
.Y(n_1680)
);

OAI332xp33_ASAP7_75t_L g1681 ( 
.A1(n_1624),
.A2(n_1591),
.A3(n_1593),
.B1(n_1612),
.B2(n_1503),
.B3(n_1599),
.C1(n_1494),
.C2(n_1589),
.Y(n_1681)
);

CKINVDCx16_ASAP7_75t_R g1682 ( 
.A(n_1634),
.Y(n_1682)
);

AOI211xp5_ASAP7_75t_L g1683 ( 
.A1(n_1649),
.A2(n_1646),
.B(n_1598),
.C(n_1554),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1646),
.A2(n_1616),
.B1(n_1613),
.B2(n_1598),
.Y(n_1684)
);

AOI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1649),
.A2(n_1613),
.B1(n_1616),
.B2(n_1598),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1630),
.B(n_1592),
.Y(n_1687)
);

OAI31xp33_ASAP7_75t_L g1688 ( 
.A1(n_1649),
.A2(n_1610),
.A3(n_1593),
.B(n_1596),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1654),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1663),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1654),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1682),
.B(n_1653),
.Y(n_1692)
);

AOI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1662),
.A2(n_1648),
.B(n_1645),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1683),
.A2(n_1613),
.B(n_1637),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1656),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1656),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1667),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1676),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1628),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1671),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1662),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1676),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1677),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_SL g1704 ( 
.A1(n_1655),
.A2(n_1632),
.B(n_1637),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1685),
.A2(n_1606),
.B(n_1604),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1672),
.B(n_1641),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1657),
.B(n_1644),
.Y(n_1707)
);

INVx4_ASAP7_75t_SL g1708 ( 
.A(n_1674),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1637),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1710)
);

INVx5_ASAP7_75t_L g1711 ( 
.A(n_1682),
.Y(n_1711)
);

CKINVDCx16_ASAP7_75t_R g1712 ( 
.A(n_1659),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1686),
.B(n_1640),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1674),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1677),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1689),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1689),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1711),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1691),
.Y(n_1719)
);

AOI21xp33_ASAP7_75t_L g1720 ( 
.A1(n_1709),
.A2(n_1670),
.B(n_1683),
.Y(n_1720)
);

NAND4xp25_ASAP7_75t_L g1721 ( 
.A(n_1704),
.B(n_1661),
.C(n_1651),
.D(n_1650),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1706),
.B(n_1679),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1691),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1693),
.Y(n_1724)
);

NOR3xp33_ASAP7_75t_L g1725 ( 
.A(n_1712),
.B(n_1668),
.C(n_1681),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1710),
.A2(n_1658),
.B1(n_1664),
.B2(n_1666),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1698),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1702),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1711),
.B(n_1669),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1715),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1693),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1706),
.B(n_1680),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1711),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1695),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1695),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1704),
.A2(n_1685),
.B(n_1673),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1696),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_L g1738 ( 
.A(n_1709),
.B(n_1703),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1707),
.B(n_1680),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1711),
.B(n_1692),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1703),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1696),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1701),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1707),
.B(n_1699),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1699),
.B(n_1701),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1711),
.B(n_1669),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1711),
.B(n_1669),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1711),
.B(n_1686),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1697),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1700),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1708),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1690),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1692),
.B(n_1652),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1713),
.B(n_1652),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1703),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1713),
.B(n_1687),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1740),
.B(n_1708),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1755),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1740),
.B(n_1708),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1725),
.B(n_1660),
.Y(n_1760)
);

NAND4xp25_ASAP7_75t_L g1761 ( 
.A(n_1720),
.B(n_1694),
.C(n_1684),
.D(n_1688),
.Y(n_1761)
);

INVxp67_ASAP7_75t_SL g1762 ( 
.A(n_1743),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1727),
.B(n_1687),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1716),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1716),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1751),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1712),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1751),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1730),
.B(n_1741),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1753),
.B(n_1708),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1717),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1717),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1732),
.B(n_1739),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1744),
.B(n_1678),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1719),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1721),
.B(n_1694),
.C(n_1637),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1719),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1753),
.B(n_1708),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1745),
.B(n_1701),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1745),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1723),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1723),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1734),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1744),
.B(n_1642),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1734),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1735),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1735),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1722),
.B(n_1642),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1751),
.B(n_1520),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1737),
.Y(n_1790)
);

NOR2x1p5_ASAP7_75t_SL g1791 ( 
.A(n_1724),
.B(n_1690),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1737),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1742),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1779),
.Y(n_1794)
);

AOI22x1_ASAP7_75t_L g1795 ( 
.A1(n_1758),
.A2(n_1736),
.B1(n_1751),
.B2(n_1718),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1760),
.A2(n_1721),
.B1(n_1726),
.B2(n_1738),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1769),
.B(n_1754),
.Y(n_1797)
);

AOI21xp33_ASAP7_75t_SL g1798 ( 
.A1(n_1776),
.A2(n_1490),
.B(n_1532),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1757),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1757),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1779),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1770),
.B(n_1738),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1780),
.B(n_1754),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1759),
.B(n_1748),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1762),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1762),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1761),
.B(n_1705),
.C(n_1742),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1780),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1759),
.B(n_1748),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1770),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1778),
.B(n_1766),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1764),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1778),
.B(n_1729),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1767),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1765),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1788),
.B(n_1756),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1766),
.Y(n_1817)
);

CKINVDCx16_ASAP7_75t_R g1818 ( 
.A(n_1789),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1771),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1773),
.B(n_1756),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1808),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1796),
.A2(n_1789),
.B1(n_1763),
.B2(n_1768),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1796),
.A2(n_1733),
.B(n_1766),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1799),
.B(n_1800),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1802),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1811),
.B(n_1768),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1804),
.Y(n_1827)
);

NAND2x1p5_ASAP7_75t_L g1828 ( 
.A(n_1802),
.B(n_1495),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1804),
.A2(n_1768),
.B1(n_1746),
.B2(n_1747),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1810),
.B(n_1772),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1814),
.B(n_1611),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1802),
.Y(n_1832)
);

NOR2x1_ASAP7_75t_L g1833 ( 
.A(n_1805),
.B(n_1775),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1805),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1803),
.B(n_1774),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1811),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1806),
.Y(n_1837)
);

OAI31xp33_ASAP7_75t_L g1838 ( 
.A1(n_1807),
.A2(n_1793),
.A3(n_1777),
.B(n_1781),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1810),
.B(n_1782),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1809),
.Y(n_1840)
);

NAND2x1_ASAP7_75t_L g1841 ( 
.A(n_1802),
.B(n_1714),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1836),
.B(n_1809),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1827),
.B(n_1813),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1833),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1832),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1836),
.B(n_1817),
.Y(n_1846)
);

NAND2x1_ASAP7_75t_SL g1847 ( 
.A(n_1825),
.B(n_1813),
.Y(n_1847)
);

INVx2_ASAP7_75t_SL g1848 ( 
.A(n_1841),
.Y(n_1848)
);

OAI222xp33_ASAP7_75t_L g1849 ( 
.A1(n_1829),
.A2(n_1795),
.B1(n_1818),
.B2(n_1806),
.C1(n_1794),
.C2(n_1801),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1831),
.B(n_1797),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1840),
.B(n_1821),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1826),
.B(n_1794),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1834),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1849),
.A2(n_1823),
.B1(n_1838),
.B2(n_1822),
.C(n_1837),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_SL g1855 ( 
.A(n_1842),
.B(n_1795),
.Y(n_1855)
);

OAI211xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1850),
.A2(n_1838),
.B(n_1824),
.C(n_1830),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1847),
.Y(n_1857)
);

O2A1O1Ixp5_ASAP7_75t_L g1858 ( 
.A1(n_1844),
.A2(n_1825),
.B(n_1801),
.C(n_1826),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1842),
.Y(n_1859)
);

CKINVDCx20_ASAP7_75t_R g1860 ( 
.A(n_1850),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1852),
.B(n_1828),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1843),
.B(n_1839),
.Y(n_1862)
);

AOI221x1_ASAP7_75t_SL g1863 ( 
.A1(n_1845),
.A2(n_1812),
.B1(n_1815),
.B2(n_1819),
.C(n_1820),
.Y(n_1863)
);

AOI21xp33_ASAP7_75t_L g1864 ( 
.A1(n_1848),
.A2(n_1828),
.B(n_1835),
.Y(n_1864)
);

AOI321xp33_ASAP7_75t_L g1865 ( 
.A1(n_1851),
.A2(n_1798),
.A3(n_1819),
.B1(n_1812),
.B2(n_1815),
.C(n_1816),
.Y(n_1865)
);

AOI221x1_ASAP7_75t_L g1866 ( 
.A1(n_1856),
.A2(n_1853),
.B1(n_1846),
.B2(n_1798),
.C(n_1783),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1860),
.Y(n_1867)
);

OAI21xp33_ASAP7_75t_SL g1868 ( 
.A1(n_1854),
.A2(n_1848),
.B(n_1786),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1859),
.Y(n_1869)
);

NAND4xp75_ASAP7_75t_L g1870 ( 
.A(n_1858),
.B(n_1791),
.C(n_1792),
.D(n_1785),
.Y(n_1870)
);

NAND2xp33_ASAP7_75t_SL g1871 ( 
.A(n_1862),
.B(n_1714),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1863),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1867),
.B(n_1857),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1868),
.B(n_1864),
.Y(n_1874)
);

NAND3xp33_ASAP7_75t_L g1875 ( 
.A(n_1872),
.B(n_1855),
.C(n_1861),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1871),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1869),
.B(n_1818),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1866),
.B(n_1729),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1870),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1872),
.B(n_1746),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1873),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1880),
.Y(n_1882)
);

INVx1_ASAP7_75t_SL g1883 ( 
.A(n_1878),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1877),
.A2(n_1789),
.B1(n_1790),
.B2(n_1787),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_R g1885 ( 
.A(n_1879),
.B(n_1495),
.Y(n_1885)
);

OR2x6_ASAP7_75t_L g1886 ( 
.A(n_1881),
.B(n_1875),
.Y(n_1886)
);

NAND2x1_ASAP7_75t_L g1887 ( 
.A(n_1882),
.B(n_1884),
.Y(n_1887)
);

AND4x2_ASAP7_75t_L g1888 ( 
.A(n_1885),
.B(n_1874),
.C(n_1876),
.D(n_1865),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1887),
.B(n_1883),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1889),
.A2(n_1886),
.B1(n_1888),
.B2(n_1611),
.Y(n_1890)
);

INVx4_ASAP7_75t_L g1891 ( 
.A(n_1890),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1890),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1892),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1891),
.A2(n_1752),
.B1(n_1784),
.B2(n_1545),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1893),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1894),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1895),
.Y(n_1897)
);

AOI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1896),
.B1(n_1752),
.B2(n_1731),
.C(n_1724),
.Y(n_1898)
);

XNOR2xp5_ASAP7_75t_L g1899 ( 
.A(n_1898),
.B(n_1747),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1752),
.B1(n_1714),
.B2(n_1724),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1731),
.B1(n_1750),
.B2(n_1749),
.Y(n_1901)
);

AOI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1901),
.A2(n_1489),
.B(n_1528),
.C(n_1509),
.Y(n_1902)
);


endmodule