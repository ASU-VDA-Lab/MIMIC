module fake_ariane_590_n_170 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_16, n_5, n_12, n_15, n_10, n_170);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_170;

wire n_83;
wire n_56;
wire n_60;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_69;
wire n_95;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_19;
wire n_40;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_111;
wire n_21;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_162;
wire n_112;
wire n_45;
wire n_138;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_121;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_22;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVxp67_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVxp33_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_27),
.B1(n_3),
.B2(n_5),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AO22x2_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_1),
.B1(n_3),
.B2(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2x1p5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_12),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_39),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_53),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2x1p5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_36),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_59),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_41),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_66),
.B(n_63),
.C(n_55),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_62),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_59),
.Y(n_94)
);

OR2x6_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_77),
.Y(n_99)
);

AOI221xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_78),
.B1(n_74),
.B2(n_73),
.C(n_82),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_49),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_82),
.Y(n_103)
);

OR2x6_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_82),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_17),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_18),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_92),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_90),
.Y(n_111)
);

NOR2x1_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_96),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_91),
.B(n_90),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_90),
.B(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_97),
.B(n_98),
.C(n_108),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

OAI21x1_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_109),
.B(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_111),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_116),
.A2(n_105),
.B(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

AO21x2_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_101),
.B(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_117),
.B(n_127),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_125),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_136),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_125),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_R g148 ( 
.A(n_143),
.B(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_129),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_132),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_130),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_129),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_132),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_150),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_135),
.C(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_148),
.C(n_149),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_154),
.Y(n_162)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_158),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_144),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_162),
.A3(n_161),
.B1(n_131),
.B2(n_121),
.C1(n_124),
.C2(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_119),
.B1(n_121),
.B2(n_131),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_138),
.B(n_113),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_166),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_113),
.B1(n_122),
.B2(n_163),
.Y(n_170)
);


endmodule