module fake_jpeg_8535_n_227 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_165;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_45),
.Y(n_70)
);

BUFx3_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_27),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_34),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_28),
.B(n_32),
.C(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_47),
.B(n_54),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_28),
.B1(n_20),
.B2(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_65),
.B1(n_21),
.B2(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_38),
.Y(n_90)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_29),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_41),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_76),
.Y(n_113)
);

AOI211xp5_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_18),
.B(n_31),
.C(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_42),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_92),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_79),
.B(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_85),
.Y(n_108)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_84),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_12),
.B1(n_14),
.B2(n_9),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_98),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_40),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_20),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_48),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_96),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_35),
.B1(n_34),
.B2(n_22),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_100),
.B1(n_56),
.B2(n_38),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_23),
.B(n_16),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_0),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_48),
.A2(n_31),
.B1(n_18),
.B2(n_20),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_99),
.A2(n_31),
.B1(n_23),
.B2(n_38),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_66),
.B1(n_61),
.B2(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_104),
.B1(n_111),
.B2(n_117),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_57),
.B1(n_56),
.B2(n_31),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_99),
.B(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_3),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_80),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_4),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_95),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_123),
.B1(n_119),
.B2(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_97),
.B1(n_94),
.B2(n_87),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_100),
.B(n_73),
.C(n_75),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_140),
.B(n_147),
.Y(n_157)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_129),
.Y(n_154)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

AO221x1_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.C(n_145),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_72),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_147),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_116),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_72),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_143),
.Y(n_151)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_71),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_89),
.B(n_90),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_102),
.C(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_120),
.B1(n_121),
.B2(n_106),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_136),
.B(n_117),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_86),
.C(n_91),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_159),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_111),
.B(n_115),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_157),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_115),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_138),
.B1(n_130),
.B2(n_129),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_182),
.B1(n_153),
.B2(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_110),
.C(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_130),
.B(n_77),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_78),
.B1(n_83),
.B2(n_101),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_176),
.B1(n_177),
.B2(n_180),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_189),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_183),
.B(n_172),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_196),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_192),
.A2(n_169),
.B1(n_184),
.B2(n_152),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_162),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_195),
.C(n_158),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_157),
.C(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_199),
.C(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_204),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_149),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_173),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_173),
.B(n_188),
.C(n_194),
.D(n_167),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_206),
.A2(n_185),
.B1(n_167),
.B2(n_165),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_194),
.B(n_178),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_122),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_206),
.A3(n_201),
.B1(n_202),
.B2(n_197),
.C1(n_205),
.C2(n_76),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_211),
.C(n_76),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_168),
.A3(n_166),
.B1(n_78),
.B2(n_79),
.C1(n_71),
.C2(n_85),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_212),
.C(n_12),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_221),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_10),
.C(n_11),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_215),
.C(n_11),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_222),
.Y(n_227)
);


endmodule