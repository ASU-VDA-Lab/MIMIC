module fake_jpeg_19932_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_58),
.B1(n_57),
.B2(n_42),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_71),
.B1(n_51),
.B2(n_46),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_59),
.B1(n_49),
.B2(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_55),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_53),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_87),
.C(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_47),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_88),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_41),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_98),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_61),
.B1(n_50),
.B2(n_45),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_100),
.B1(n_11),
.B2(n_12),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_40),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_106),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_2),
.B(n_10),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_113),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_111),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.C(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_115),
.A2(n_104),
.B1(n_109),
.B2(n_101),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_114),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_100),
.B(n_110),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_15),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_16),
.C(n_17),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_116),
.A3(n_20),
.B1(n_21),
.B2(n_22),
.C1(n_26),
.C2(n_27),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_108),
.B1(n_28),
.B2(n_30),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_18),
.Y(n_128)
);


endmodule