module fake_netlist_5_1803_n_1682 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1682);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1682;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g156 ( 
.A(n_12),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_38),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_48),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_70),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_67),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_99),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_18),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_54),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_83),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_84),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_77),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_131),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_46),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_75),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_47),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_19),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_152),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_59),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_130),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_7),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_37),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_53),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_85),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_117),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_64),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_28),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_55),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_137),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_145),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_88),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_110),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_80),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_33),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_58),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_22),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_39),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_24),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_34),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_38),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_9),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_111),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_74),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_69),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_73),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_37),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_12),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_122),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_1),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_9),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_90),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_54),
.Y(n_234)
);

BUFx2_ASAP7_75t_SL g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_108),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_78),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_40),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_102),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_126),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_79),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_29),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_1),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_112),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_28),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_93),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_14),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_87),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_129),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_58),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_92),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_139),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_82),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_14),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_57),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_27),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_33),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_45),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_113),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_68),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_49),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_13),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_132),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_81),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_16),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_48),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_42),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_76),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_19),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_10),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_89),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_36),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_123),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_97),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_52),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_66),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_142),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_24),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_133),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_31),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_61),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_44),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_148),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_153),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_91),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_50),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_121),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_18),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_3),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_50),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_53),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_120),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_10),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_65),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_56),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_6),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_114),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_115),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_29),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_25),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_98),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_51),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_40),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_162),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_166),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_171),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_2),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_170),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_172),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_225),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_186),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_174),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_222),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_178),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_254),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_183),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_288),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_187),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_193),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_256),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_177),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_177),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_184),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_194),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_213),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_195),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_213),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_272),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_196),
.Y(n_343)
);

BUFx2_ASAP7_75t_SL g344 ( 
.A(n_219),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_198),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_200),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_201),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_286),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_205),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_167),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_280),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_257),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_206),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_167),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_246),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_156),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_161),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_156),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_219),
.B(n_3),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_163),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_163),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_169),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_182),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_182),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_211),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_249),
.B(n_4),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_169),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_176),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_180),
.B(n_5),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_223),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_182),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_176),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_263),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_224),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_179),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_249),
.B(n_6),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_179),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_263),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_321),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_263),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_368),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_275),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_275),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_334),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_311),
.B(n_293),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_293),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_361),
.B(n_228),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_362),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_364),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_335),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_363),
.B(n_204),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_335),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_344),
.B(n_353),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_311),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_316),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_310),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_344),
.B(n_257),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_312),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_365),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_354),
.B(n_159),
.Y(n_426)
);

AND3x1_ASAP7_75t_L g427 ( 
.A(n_314),
.B(n_274),
.C(n_181),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_354),
.B(n_232),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_336),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_355),
.B(n_236),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_355),
.B(n_240),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_380),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_365),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_338),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_358),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_366),
.B(n_242),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_359),
.B(n_188),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_371),
.B(n_210),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_R g441 ( 
.A(n_313),
.B(n_233),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_371),
.B(n_248),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_319),
.B(n_233),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_316),
.B(n_250),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_372),
.B(n_210),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_385),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_318),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_398),
.Y(n_451)
);

INVx5_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_398),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_396),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_421),
.B(n_322),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_413),
.A2(n_352),
.B1(n_259),
.B2(n_380),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_385),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_325),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_421),
.B(n_327),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_384),
.B(n_426),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_383),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_420),
.B(n_330),
.Y(n_467)
);

BUFx4f_ASAP7_75t_L g468 ( 
.A(n_413),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_413),
.A2(n_259),
.B1(n_274),
.B2(n_309),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_331),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_384),
.B(n_339),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_428),
.B(n_356),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_386),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_SL g479 ( 
.A(n_444),
.B(n_212),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_408),
.B(n_337),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_423),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_413),
.A2(n_260),
.B1(n_192),
.B2(n_191),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_396),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_387),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_412),
.B(n_340),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_418),
.Y(n_489)
);

BUFx8_ASAP7_75t_SL g490 ( 
.A(n_446),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_391),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_443),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_412),
.B(n_343),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_443),
.B(n_346),
.C(n_345),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_422),
.B(n_347),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_422),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_393),
.B(n_204),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_432),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_432),
.B(n_349),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_428),
.B(n_357),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_417),
.B(n_374),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_401),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

CKINVDCx14_ASAP7_75t_R g507 ( 
.A(n_399),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_391),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_417),
.B(n_264),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_444),
.A2(n_235),
.B1(n_309),
.B2(n_191),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_384),
.B(n_339),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_393),
.B(n_204),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_394),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_394),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_396),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_439),
.B(n_369),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_430),
.B(n_378),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_413),
.B(n_204),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_395),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_427),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_430),
.B(n_431),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_417),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_390),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_395),
.Y(n_527)
);

INVx2_ASAP7_75t_SL g528 ( 
.A(n_405),
.Y(n_528)
);

BUFx8_ASAP7_75t_SL g529 ( 
.A(n_399),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_402),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_388),
.B(n_159),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_439),
.B(n_315),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_413),
.A2(n_265),
.B1(n_227),
.B2(n_230),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_426),
.B(n_341),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_389),
.B(n_307),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_427),
.A2(n_373),
.B1(n_221),
.B2(n_234),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_389),
.B(n_405),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_406),
.B(n_320),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_405),
.B(n_267),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_441),
.A2(n_342),
.B1(n_332),
.B2(n_326),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_406),
.B(n_238),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_416),
.B(n_235),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_445),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_402),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_413),
.A2(n_243),
.B1(n_255),
.B2(n_230),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_410),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_405),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_405),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_413),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_441),
.A2(n_245),
.B1(n_308),
.B2(n_231),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_388),
.B(n_277),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_438),
.B(n_250),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_440),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_438),
.B(n_250),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_437),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_437),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_402),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_402),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_402),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_440),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_388),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_413),
.B(n_204),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_414),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_426),
.B(n_341),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_442),
.B(n_323),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_416),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_442),
.B(n_192),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_414),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_388),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_425),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_393),
.B(n_425),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_393),
.B(n_278),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_433),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_440),
.B(n_197),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_390),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_402),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_402),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_433),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_393),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_440),
.B(n_250),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_445),
.A2(n_243),
.B1(n_306),
.B2(n_305),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_392),
.B(n_204),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g586 ( 
.A(n_436),
.B(n_215),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_392),
.B(n_279),
.C(n_158),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_436),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_390),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_403),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_390),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_445),
.B(n_197),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_445),
.B(n_216),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_390),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_544),
.B(n_372),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_448),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_449),
.B(n_419),
.Y(n_597)
);

BUFx5_ASAP7_75t_L g598 ( 
.A(n_493),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_472),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_480),
.B(n_419),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_471),
.A2(n_216),
.B1(n_306),
.B2(n_305),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_468),
.B(n_268),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_540),
.A2(n_445),
.B(n_227),
.C(n_255),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_524),
.A2(n_268),
.B(n_251),
.C(n_173),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_448),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_569),
.B(n_281),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_447),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_481),
.B(n_241),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_472),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_497),
.B(n_218),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_524),
.B(n_464),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_464),
.B(n_419),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_450),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_528),
.B(n_419),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_468),
.B(n_285),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_497),
.B(n_157),
.Y(n_616)
);

INVx8_ASAP7_75t_L g617 ( 
.A(n_545),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_528),
.B(n_419),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_586),
.A2(n_270),
.B1(n_297),
.B2(n_260),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_550),
.B(n_525),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_499),
.B(n_160),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_544),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_450),
.Y(n_623)
);

O2A1O1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_538),
.A2(n_270),
.B(n_261),
.C(n_265),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_447),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_550),
.B(n_429),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_468),
.B(n_289),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_493),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_582),
.Y(n_629)
);

OAI221xp5_ASAP7_75t_L g630 ( 
.A1(n_584),
.A2(n_261),
.B1(n_297),
.B2(n_189),
.C(n_202),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_510),
.A2(n_483),
.B1(n_548),
.B2(n_535),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_510),
.A2(n_189),
.B1(n_253),
.B2(n_251),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_499),
.B(n_168),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_552),
.B(n_290),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_552),
.B(n_291),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_574),
.B(n_429),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_574),
.B(n_429),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_541),
.B(n_190),
.C(n_199),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_475),
.B(n_451),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_476),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_465),
.B(n_429),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_454),
.Y(n_642)
);

BUFx8_ASAP7_75t_L g643 ( 
.A(n_523),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_476),
.B(n_429),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_454),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_501),
.B(n_175),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_501),
.B(n_208),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_511),
.B(n_434),
.Y(n_648)
);

AND2x6_ASAP7_75t_SL g649 ( 
.A(n_534),
.B(n_376),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_458),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_518),
.A2(n_298),
.B1(n_303),
.B2(n_304),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g652 ( 
.A(n_481),
.B(n_484),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_511),
.B(n_434),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_475),
.B(n_376),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_451),
.B(n_434),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_453),
.B(n_434),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_457),
.A2(n_165),
.B1(n_173),
.B2(n_185),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_453),
.B(n_434),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_477),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_495),
.B(n_411),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_533),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_537),
.B(n_379),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_582),
.B(n_533),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_568),
.A2(n_572),
.B1(n_479),
.B2(n_570),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_552),
.B(n_164),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_551),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_456),
.B(n_214),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_536),
.B(n_397),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_536),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_537),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_566),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_458),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_484),
.B(n_244),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_566),
.B(n_397),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_492),
.B(n_218),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_572),
.A2(n_164),
.B1(n_165),
.B2(n_185),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_571),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_587),
.B(n_282),
.C(n_217),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_571),
.B(n_397),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_460),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_460),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_503),
.B(n_397),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_567),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_556),
.B(n_202),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_462),
.B(n_220),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_504),
.B(n_397),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_564),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_505),
.B(n_400),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_564),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_506),
.B(n_400),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_570),
.A2(n_283),
.B1(n_207),
.B2(n_209),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_556),
.B(n_203),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_461),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_532),
.A2(n_522),
.B(n_549),
.C(n_515),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_492),
.B(n_218),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_529),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_519),
.B(n_400),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_531),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_531),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_492),
.B(n_247),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_573),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_567),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_459),
.B(n_203),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_545),
.B(n_218),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_576),
.B(n_400),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_570),
.A2(n_287),
.B1(n_209),
.B2(n_229),
.Y(n_707)
);

AND2x6_ASAP7_75t_L g708 ( 
.A(n_532),
.B(n_207),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_581),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_532),
.A2(n_283),
.B(n_229),
.C(n_300),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_588),
.A2(n_300),
.B(n_237),
.C(n_287),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_479),
.A2(n_570),
.B1(n_517),
.B2(n_542),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_553),
.B(n_545),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_523),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_556),
.B(n_237),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_554),
.A2(n_253),
.B1(n_239),
.B2(n_273),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_478),
.B(n_400),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_563),
.B(n_239),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_545),
.B(n_226),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_510),
.A2(n_271),
.B1(n_284),
.B2(n_302),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_478),
.B(n_435),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_482),
.B(n_435),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_482),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_485),
.B(n_435),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_555),
.A2(n_435),
.B1(n_415),
.B2(n_403),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_485),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_510),
.A2(n_226),
.B1(n_379),
.B2(n_381),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_563),
.B(n_403),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_563),
.B(n_403),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_487),
.B(n_403),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_488),
.B(n_252),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_487),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_514),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_514),
.B(n_435),
.Y(n_734)
);

OR2x6_ASAP7_75t_L g735 ( 
.A(n_577),
.B(n_381),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_526),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_577),
.A2(n_295),
.B1(n_258),
.B2(n_276),
.C(n_266),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_520),
.A2(n_226),
.B1(n_301),
.B2(n_299),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_520),
.A2(n_226),
.B1(n_269),
.B2(n_292),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_494),
.B(n_294),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_526),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_466),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_526),
.B(n_435),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_551),
.B(n_435),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_557),
.A2(n_415),
.B1(n_403),
.B2(n_411),
.Y(n_745)
);

INVxp33_ASAP7_75t_L g746 ( 
.A(n_490),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_578),
.B(n_415),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_578),
.Y(n_748)
);

NOR2x1p5_ASAP7_75t_L g749 ( 
.A(n_489),
.B(n_350),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_531),
.B(n_546),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_578),
.B(n_415),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_531),
.B(n_415),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_466),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_577),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_496),
.B(n_415),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_591),
.B(n_415),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_591),
.B(n_403),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_591),
.B(n_411),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_473),
.B(n_350),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_469),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_502),
.B(n_348),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_469),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_509),
.B(n_348),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_531),
.B(n_154),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_575),
.A2(n_151),
.B1(n_147),
.B2(n_146),
.Y(n_765)
);

NAND2x1p5_ASAP7_75t_L g766 ( 
.A(n_667),
.B(n_546),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_611),
.A2(n_546),
.B1(n_500),
.B2(n_551),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_622),
.B(n_467),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_646),
.B(n_558),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_620),
.A2(n_546),
.B(n_565),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_681),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_658),
.A2(n_565),
.B(n_585),
.C(n_592),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_750),
.A2(n_546),
.B(n_516),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_750),
.A2(n_516),
.B(n_583),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_599),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_682),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_597),
.A2(n_516),
.B(n_579),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_646),
.A2(n_594),
.B(n_589),
.C(n_543),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_640),
.B(n_491),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_699),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_600),
.A2(n_530),
.B(n_560),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_662),
.B(n_491),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_604),
.A2(n_585),
.B(n_593),
.C(n_592),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_670),
.B(n_508),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_728),
.A2(n_530),
.B(n_560),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_672),
.B(n_508),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_728),
.A2(n_547),
.B(n_562),
.Y(n_788)
);

BUFx4f_ASAP7_75t_L g789 ( 
.A(n_617),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_647),
.B(n_558),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_729),
.A2(n_700),
.B(n_612),
.Y(n_791)
);

OAI22xp33_ASAP7_75t_L g792 ( 
.A1(n_712),
.A2(n_593),
.B1(n_592),
.B2(n_577),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_671),
.B(n_592),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_729),
.A2(n_700),
.B(n_690),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_690),
.A2(n_561),
.B(n_547),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_694),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_665),
.B(n_489),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_678),
.B(n_513),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_690),
.A2(n_562),
.B(n_590),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_690),
.A2(n_561),
.B(n_590),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_723),
.B(n_513),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_684),
.B(n_559),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_726),
.B(n_732),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_559),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_760),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_744),
.A2(n_580),
.B(n_579),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_733),
.B(n_521),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_703),
.B(n_521),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_644),
.A2(n_593),
.B(n_527),
.C(n_539),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_595),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_629),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_752),
.A2(n_594),
.B(n_527),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_614),
.A2(n_580),
.B(n_455),
.Y(n_813)
);

NOR2x1_ASAP7_75t_L g814 ( 
.A(n_638),
.B(n_593),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_653),
.B(n_507),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_759),
.B(n_761),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_754),
.B(n_486),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_618),
.A2(n_455),
.B(n_474),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_660),
.B(n_490),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_626),
.A2(n_637),
.B(n_636),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_648),
.A2(n_455),
.B(n_474),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_713),
.A2(n_512),
.B1(n_498),
.B2(n_486),
.Y(n_822)
);

OAI21xp33_ASAP7_75t_L g823 ( 
.A1(n_616),
.A2(n_463),
.B(n_470),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_654),
.A2(n_455),
.B(n_474),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_742),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_639),
.B(n_470),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_762),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_656),
.A2(n_455),
.B(n_474),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_639),
.B(n_486),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_657),
.A2(n_474),
.B(n_470),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_602),
.A2(n_463),
.B(n_498),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_763),
.B(n_463),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_659),
.A2(n_452),
.B(n_512),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_602),
.A2(n_512),
.B(n_498),
.C(n_452),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_610),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_702),
.B(n_512),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_713),
.A2(n_512),
.B(n_498),
.C(n_452),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_664),
.A2(n_452),
.B(n_512),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_709),
.B(n_498),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_668),
.B(n_452),
.Y(n_840)
);

BUFx12f_ASAP7_75t_L g841 ( 
.A(n_643),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_701),
.B(n_714),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_615),
.A2(n_498),
.B(n_144),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_701),
.B(n_529),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_629),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_615),
.A2(n_140),
.B(n_134),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_SL g847 ( 
.A1(n_631),
.A2(n_8),
.B(n_15),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_627),
.A2(n_128),
.B(n_118),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_596),
.B(n_8),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_699),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_627),
.A2(n_116),
.B(n_107),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_616),
.B(n_15),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_753),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_605),
.B(n_17),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_632),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_621),
.B(n_633),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_676),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_631),
.A2(n_104),
.B1(n_101),
.B2(n_100),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_696),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_613),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_634),
.A2(n_96),
.B(n_86),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_621),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_SL g863 ( 
.A1(n_666),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_655),
.B(n_23),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_688),
.A2(n_72),
.B1(n_62),
.B2(n_60),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_606),
.B(n_668),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_623),
.B(n_26),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_663),
.B(n_633),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_736),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_632),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_663),
.B(n_655),
.Y(n_871)
);

O2A1O1Ixp5_ASAP7_75t_L g872 ( 
.A1(n_666),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_741),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_686),
.B(n_32),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_661),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_634),
.A2(n_35),
.B(n_39),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_686),
.B(n_699),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_635),
.A2(n_41),
.B(n_42),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_679),
.B(n_41),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_699),
.B(n_755),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_695),
.A2(n_43),
.B(n_44),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_635),
.A2(n_45),
.B(n_47),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_667),
.B(n_49),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_608),
.B(n_51),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_628),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_752),
.A2(n_743),
.B(n_756),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_619),
.B(n_598),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_747),
.A2(n_757),
.B(n_751),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_705),
.B(n_719),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_748),
.B(n_715),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_641),
.A2(n_758),
.B(n_764),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_755),
.B(n_598),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_607),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_685),
.A2(n_718),
.B(n_693),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_735),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_685),
.A2(n_718),
.B(n_693),
.Y(n_896)
);

CKINVDCx10_ASAP7_75t_R g897 ( 
.A(n_746),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_619),
.B(n_598),
.Y(n_898)
);

AOI21x1_ASAP7_75t_L g899 ( 
.A1(n_721),
.A2(n_722),
.B(n_734),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_715),
.A2(n_730),
.B(n_724),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_598),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_735),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_710),
.A2(n_711),
.B(n_692),
.C(n_707),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_598),
.B(n_727),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_603),
.A2(n_716),
.B(n_630),
.C(n_624),
.Y(n_905)
);

NAND2x1p5_ASAP7_75t_L g906 ( 
.A(n_625),
.B(n_645),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_598),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_642),
.Y(n_908)
);

OR2x6_ASAP7_75t_L g909 ( 
.A(n_617),
.B(n_735),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_727),
.B(n_731),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_731),
.B(n_740),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_740),
.B(n_674),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_669),
.B(n_675),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_680),
.B(n_717),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_749),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_683),
.A2(n_689),
.B(n_687),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_765),
.A2(n_704),
.B(n_706),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_650),
.B(n_673),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_691),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_698),
.A2(n_725),
.B(n_745),
.Y(n_920)
);

OAI21xp33_ASAP7_75t_L g921 ( 
.A1(n_720),
.A2(n_601),
.B(n_739),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_677),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_601),
.A2(n_617),
.B(n_737),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_651),
.A2(n_708),
.B(n_739),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_720),
.A2(n_738),
.B(n_652),
.C(n_708),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_708),
.B(n_738),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_708),
.A2(n_649),
.B(n_697),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_708),
.A2(n_643),
.B(n_647),
.C(n_646),
.Y(n_928)
);

AO21x1_ASAP7_75t_L g929 ( 
.A1(n_666),
.A2(n_602),
.B(n_479),
.Y(n_929)
);

AOI21xp33_ASAP7_75t_L g930 ( 
.A1(n_646),
.A2(n_647),
.B(n_668),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_620),
.A2(n_552),
.B(n_468),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_620),
.A2(n_552),
.B(n_468),
.Y(n_932)
);

AOI21xp33_ASAP7_75t_L g933 ( 
.A1(n_646),
.A2(n_647),
.B(n_668),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_611),
.B(n_622),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_620),
.A2(n_552),
.B(n_468),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_611),
.B(n_569),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_611),
.B(n_569),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_611),
.B(n_569),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_611),
.B(n_569),
.Y(n_939)
);

AND2x2_ASAP7_75t_SL g940 ( 
.A(n_632),
.B(n_727),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_611),
.B(n_665),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_760),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_599),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_620),
.A2(n_552),
.B(n_468),
.Y(n_944)
);

INVx11_ASAP7_75t_L g945 ( 
.A(n_643),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_646),
.A2(n_647),
.B(n_713),
.C(n_686),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_699),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_681),
.Y(n_948)
);

AND2x4_ASAP7_75t_SL g949 ( 
.A(n_599),
.B(n_315),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_612),
.A2(n_620),
.B(n_636),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_620),
.A2(n_552),
.B(n_468),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_617),
.B(n_599),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_690),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_856),
.A2(n_930),
.B(n_933),
.C(n_946),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_897),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_911),
.B(n_856),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_862),
.B(n_936),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_787),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_874),
.A2(n_910),
.B(n_852),
.C(n_912),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_892),
.A2(n_932),
.B(n_931),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_937),
.B(n_938),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_949),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_939),
.B(n_934),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_934),
.B(n_862),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_SL g965 ( 
.A(n_769),
.B(n_804),
.C(n_790),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_943),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_866),
.A2(n_852),
.B(n_921),
.C(n_924),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_850),
.B(n_947),
.Y(n_968)
);

AO21x1_ASAP7_75t_L g969 ( 
.A1(n_881),
.A2(n_941),
.B(n_792),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_850),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_860),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_771),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_776),
.Y(n_973)
);

NOR2x1_ASAP7_75t_SL g974 ( 
.A(n_850),
.B(n_947),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_940),
.B(n_868),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_810),
.B(n_842),
.Y(n_976)
);

XNOR2xp5_ASAP7_75t_L g977 ( 
.A(n_889),
.B(n_797),
.Y(n_977)
);

O2A1O1Ixp5_ASAP7_75t_L g978 ( 
.A1(n_917),
.A2(n_877),
.B(n_929),
.C(n_840),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_835),
.B(n_857),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_816),
.B(n_940),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_943),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_803),
.B(n_835),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_775),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_945),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_855),
.A2(n_870),
.B1(n_858),
.B2(n_887),
.Y(n_985)
);

BUFx2_ASAP7_75t_SL g986 ( 
.A(n_895),
.Y(n_986)
);

CKINVDCx10_ASAP7_75t_R g987 ( 
.A(n_841),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_880),
.A2(n_812),
.B(n_899),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_796),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_871),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_782),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_784),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_792),
.B(n_767),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_935),
.A2(n_944),
.B(n_951),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_894),
.A2(n_896),
.B(n_907),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_901),
.A2(n_907),
.B(n_770),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_901),
.A2(n_950),
.B(n_791),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_915),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_859),
.B(n_768),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_786),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_895),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_815),
.B(n_884),
.Y(n_1002)
);

INVx6_ASAP7_75t_L g1003 ( 
.A(n_895),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_925),
.A2(n_778),
.B(n_849),
.C(n_867),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_798),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_909),
.B(n_895),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_854),
.A2(n_898),
.B(n_885),
.C(n_922),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_904),
.B(n_923),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_779),
.B(n_808),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_919),
.B(n_780),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_850),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_947),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_844),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_947),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_815),
.B(n_802),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_820),
.A2(n_794),
.B(n_891),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_793),
.B(n_902),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_793),
.B(n_811),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_801),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_819),
.Y(n_1020)
);

INVxp33_ASAP7_75t_L g1021 ( 
.A(n_819),
.Y(n_1021)
);

AO32x1_ASAP7_75t_L g1022 ( 
.A1(n_865),
.A2(n_805),
.A3(n_827),
.B1(n_942),
.B2(n_873),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_902),
.B(n_864),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_909),
.B(n_825),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_909),
.B(n_789),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_952),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_953),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_847),
.A2(n_928),
.B(n_863),
.C(n_882),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_780),
.A2(n_870),
.B1(n_855),
.B2(n_926),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_952),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_807),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_876),
.A2(n_878),
.B1(n_875),
.B2(n_879),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_L g1033 ( 
.A1(n_920),
.A2(n_834),
.B(n_916),
.C(n_774),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_883),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_913),
.A2(n_914),
.B(n_900),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_953),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_893),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_773),
.A2(n_888),
.B(n_821),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_SL g1039 ( 
.A(n_927),
.B(n_905),
.C(n_883),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_853),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_948),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_811),
.B(n_845),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_845),
.B(n_817),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_869),
.B(n_817),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_918),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_832),
.B(n_829),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_809),
.A2(n_872),
.B(n_905),
.C(n_903),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_809),
.A2(n_783),
.B(n_903),
.C(n_772),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_766),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_766),
.Y(n_1050)
);

CKINVDCx14_ASAP7_75t_R g1051 ( 
.A(n_789),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_826),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_814),
.B(n_890),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_906),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_906),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_886),
.B(n_890),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_824),
.A2(n_777),
.B(n_818),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_952),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_836),
.Y(n_1059)
);

NAND2x1p5_ASAP7_75t_L g1060 ( 
.A(n_822),
.B(n_851),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_SL g1061 ( 
.A(n_846),
.B(n_861),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_828),
.A2(n_830),
.B(n_813),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_872),
.A2(n_837),
.B(n_783),
.C(n_772),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_781),
.A2(n_795),
.B(n_799),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_823),
.B(n_839),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_785),
.A2(n_788),
.B(n_800),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_831),
.A2(n_843),
.B(n_838),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_806),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_848),
.B(n_834),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_833),
.B(n_930),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_892),
.A2(n_552),
.B(n_468),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_850),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_930),
.B(n_933),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_892),
.A2(n_552),
.B(n_468),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_L g1075 ( 
.A(n_930),
.B(n_933),
.C(n_911),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_930),
.B(n_933),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_856),
.A2(n_930),
.B(n_933),
.C(n_946),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_856),
.A2(n_911),
.B1(n_933),
.B2(n_930),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_946),
.A2(n_911),
.B1(n_856),
.B2(n_910),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_856),
.B(n_936),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_787),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_930),
.B(n_933),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_949),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_856),
.A2(n_911),
.B1(n_933),
.B2(n_930),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_946),
.A2(n_911),
.B1(n_856),
.B2(n_910),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_856),
.B(n_936),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_856),
.B(n_936),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_856),
.B(n_936),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_850),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_930),
.B(n_933),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_892),
.A2(n_552),
.B(n_468),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_892),
.A2(n_552),
.B(n_468),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_892),
.A2(n_552),
.B(n_468),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_787),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_930),
.B(n_933),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_930),
.B(n_933),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_908),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1035),
.A2(n_1016),
.B(n_997),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_965),
.A2(n_1077),
.B(n_1096),
.C(n_1090),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_SL g1100 ( 
.A(n_984),
.B(n_1001),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_971),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_985),
.A2(n_956),
.B1(n_1078),
.B2(n_1084),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_956),
.B(n_1080),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_996),
.A2(n_994),
.B(n_995),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1086),
.B(n_1087),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_960),
.A2(n_1066),
.B(n_1038),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1088),
.B(n_963),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1025),
.B(n_1006),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_961),
.B(n_964),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1082),
.A2(n_1090),
.B(n_1096),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_970),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1082),
.B(n_1075),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1079),
.A2(n_1085),
.B(n_1008),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1057),
.A2(n_1056),
.A3(n_1067),
.B(n_1062),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1075),
.A2(n_1076),
.B1(n_1073),
.B2(n_1095),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_976),
.A2(n_1002),
.B1(n_1015),
.B2(n_1095),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1008),
.A2(n_1071),
.B(n_1074),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1091),
.A2(n_1093),
.B(n_1092),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_959),
.B(n_999),
.C(n_1032),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_980),
.B(n_991),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1033),
.A2(n_1069),
.B(n_1004),
.Y(n_1121)
);

AO21x2_ASAP7_75t_L g1122 ( 
.A1(n_993),
.A2(n_1039),
.B(n_1070),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1064),
.A2(n_988),
.B(n_1068),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1068),
.A2(n_978),
.B(n_1069),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_957),
.B(n_1009),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_981),
.Y(n_1126)
);

CKINVDCx11_ASAP7_75t_R g1127 ( 
.A(n_1083),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_982),
.B(n_958),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_976),
.B(n_1023),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1046),
.A2(n_993),
.B(n_1047),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_992),
.B(n_1000),
.Y(n_1131)
);

NOR3xp33_ASAP7_75t_L g1132 ( 
.A(n_1013),
.B(n_999),
.C(n_1015),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1063),
.A2(n_985),
.B(n_1053),
.Y(n_1133)
);

AOI221x1_ASAP7_75t_L g1134 ( 
.A1(n_1029),
.A2(n_1065),
.B1(n_979),
.B2(n_1005),
.C(n_1031),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1060),
.A2(n_1028),
.B(n_1053),
.Y(n_1135)
);

AO21x1_ASAP7_75t_L g1136 ( 
.A1(n_975),
.A2(n_1007),
.B(n_1060),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1032),
.A2(n_1019),
.B1(n_975),
.B2(n_1010),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1017),
.B(n_990),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_990),
.B(n_979),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_1081),
.B(n_1094),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_966),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1021),
.B(n_977),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1037),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_966),
.B(n_1024),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1020),
.B(n_983),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_968),
.A2(n_1045),
.B(n_974),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_SL g1147 ( 
.A(n_1030),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1034),
.B(n_1044),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1018),
.A2(n_1052),
.B(n_1044),
.C(n_1040),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1052),
.B(n_1059),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_SL g1151 ( 
.A1(n_1043),
.A2(n_1011),
.B(n_1022),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_986),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1042),
.A2(n_1022),
.B(n_1054),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_SL g1154 ( 
.A1(n_1042),
.A2(n_1055),
.B(n_1011),
.C(n_1041),
.Y(n_1154)
);

NOR4xp25_ASAP7_75t_L g1155 ( 
.A(n_972),
.B(n_1097),
.C(n_973),
.D(n_989),
.Y(n_1155)
);

AOI221x1_ASAP7_75t_L g1156 ( 
.A1(n_1022),
.A2(n_1050),
.B1(n_1049),
.B2(n_1061),
.C(n_1014),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1006),
.A2(n_1003),
.B1(n_1058),
.B2(n_1051),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1049),
.A2(n_1050),
.B(n_1014),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1058),
.A2(n_1027),
.B(n_1072),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1058),
.A2(n_998),
.B(n_1027),
.C(n_1036),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1006),
.Y(n_1161)
);

AO21x1_ASAP7_75t_L g1162 ( 
.A1(n_1072),
.A2(n_1089),
.B(n_1027),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_962),
.B(n_955),
.C(n_1036),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1089),
.A2(n_1036),
.B(n_1003),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1026),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_970),
.A2(n_1012),
.B(n_1003),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1012),
.A2(n_969),
.A3(n_1048),
.B(n_967),
.Y(n_1167)
);

AOI221x1_ASAP7_75t_L g1168 ( 
.A1(n_1012),
.A2(n_987),
.B1(n_930),
.B2(n_933),
.C(n_946),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1012),
.A2(n_967),
.B(n_954),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_996),
.A2(n_994),
.B(n_995),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_956),
.B(n_1080),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_971),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_SL g1173 ( 
.A1(n_954),
.A2(n_946),
.B(n_1077),
.C(n_930),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_967),
.A2(n_1077),
.B(n_954),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_996),
.A2(n_994),
.B(n_995),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_956),
.B(n_1080),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_971),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_956),
.A2(n_933),
.B1(n_930),
.B2(n_619),
.C(n_1082),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_971),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_967),
.A2(n_1077),
.B(n_954),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_969),
.A2(n_1048),
.A3(n_967),
.B(n_954),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_961),
.B(n_1080),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_981),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_971),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_965),
.B(n_956),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_987),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_981),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_967),
.A2(n_1077),
.B(n_954),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_956),
.A2(n_933),
.B(n_930),
.C(n_856),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_956),
.A2(n_933),
.B(n_930),
.C(n_856),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_956),
.A2(n_933),
.B(n_930),
.C(n_856),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_996),
.A2(n_994),
.B(n_995),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_969),
.A2(n_1048),
.A3(n_967),
.B(n_954),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_965),
.A2(n_946),
.B(n_933),
.C(n_930),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_971),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_967),
.A2(n_1077),
.B(n_954),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_969),
.A2(n_1048),
.A3(n_967),
.B(n_954),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_985),
.A2(n_956),
.B1(n_940),
.B2(n_855),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_954),
.A2(n_946),
.B(n_1077),
.C(n_930),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_971),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_971),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_966),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_969),
.A2(n_1048),
.A3(n_967),
.B(n_954),
.Y(n_1206)
);

CKINVDCx11_ASAP7_75t_R g1207 ( 
.A(n_1083),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_SL g1208 ( 
.A(n_1082),
.B(n_940),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_SL g1209 ( 
.A1(n_954),
.A2(n_946),
.B(n_1077),
.C(n_930),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_996),
.A2(n_994),
.B(n_995),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_971),
.Y(n_1212)
);

AOI221x1_ASAP7_75t_L g1213 ( 
.A1(n_954),
.A2(n_930),
.B1(n_933),
.B2(n_946),
.C(n_1077),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_961),
.B(n_1080),
.Y(n_1215)
);

INVx3_ASAP7_75t_SL g1216 ( 
.A(n_984),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1082),
.A2(n_856),
.B1(n_1096),
.B2(n_1090),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1078),
.A2(n_911),
.B1(n_608),
.B2(n_586),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_966),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_985),
.A2(n_956),
.B1(n_940),
.B2(n_855),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_971),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_956),
.B(n_1080),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_969),
.A2(n_1048),
.A3(n_967),
.B(n_954),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1035),
.A2(n_552),
.B(n_468),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_956),
.B(n_1080),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_965),
.B(n_956),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_956),
.A2(n_933),
.B(n_930),
.C(n_856),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1219),
.B2(n_1102),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1200),
.A2(n_1223),
.B1(n_1208),
.B2(n_1231),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1167),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1110),
.A2(n_1102),
.B1(n_1200),
.B2(n_1223),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1171),
.B(n_1177),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1230),
.A2(n_1232),
.B1(n_1190),
.B2(n_1191),
.Y(n_1238)
);

BUFx10_ASAP7_75t_L g1239 ( 
.A(n_1145),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1129),
.B(n_1138),
.Y(n_1240)
);

BUFx2_ASAP7_75t_SL g1241 ( 
.A(n_1147),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1186),
.A2(n_1112),
.B1(n_1208),
.B2(n_1119),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1202),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1192),
.A2(n_1116),
.B1(n_1227),
.B2(n_1105),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1220),
.A2(n_1181),
.B1(n_1189),
.B2(n_1174),
.Y(n_1245)
);

INVxp67_ASAP7_75t_SL g1246 ( 
.A(n_1205),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1174),
.A2(n_1189),
.B1(n_1198),
.B2(n_1181),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1198),
.A2(n_1227),
.B1(n_1113),
.B2(n_1142),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1183),
.B(n_1215),
.Y(n_1249)
);

BUFx2_ASAP7_75t_SL g1250 ( 
.A(n_1147),
.Y(n_1250)
);

INVx6_ASAP7_75t_L g1251 ( 
.A(n_1108),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1115),
.A2(n_1113),
.B1(n_1133),
.B2(n_1132),
.Y(n_1252)
);

CKINVDCx8_ASAP7_75t_R g1253 ( 
.A(n_1187),
.Y(n_1253)
);

BUFx10_ASAP7_75t_L g1254 ( 
.A(n_1221),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_1140),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1130),
.A2(n_1109),
.B1(n_1136),
.B2(n_1120),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1163),
.A2(n_1108),
.B1(n_1188),
.B2(n_1126),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1139),
.A2(n_1148),
.B1(n_1169),
.B2(n_1157),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1101),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1126),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_SL g1261 ( 
.A(n_1111),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1207),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1120),
.B(n_1125),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1169),
.A2(n_1157),
.B1(n_1131),
.B2(n_1161),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1188),
.A2(n_1165),
.B1(n_1152),
.B2(n_1128),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1111),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_1172),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1216),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1213),
.A2(n_1168),
.B1(n_1150),
.B2(n_1134),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1122),
.A2(n_1137),
.B1(n_1152),
.B2(n_1141),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1184),
.Y(n_1271)
);

AOI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1137),
.A2(n_1173),
.B1(n_1209),
.B2(n_1201),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1178),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1122),
.A2(n_1143),
.B1(n_1197),
.B2(n_1203),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1180),
.A2(n_1224),
.B1(n_1212),
.B2(n_1144),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1121),
.A2(n_1099),
.B1(n_1135),
.B2(n_1195),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1149),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1154),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1158),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1162),
.Y(n_1280)
);

BUFx2_ASAP7_75t_SL g1281 ( 
.A(n_1166),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1164),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_1100),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1146),
.A2(n_1153),
.B1(n_1098),
.B2(n_1117),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_SL g1285 ( 
.A1(n_1164),
.A2(n_1160),
.B1(n_1228),
.B2(n_1199),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1182),
.A2(n_1194),
.B1(n_1228),
.B2(n_1206),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1155),
.Y(n_1287)
);

OAI22x1_ASAP7_75t_SL g1288 ( 
.A1(n_1159),
.A2(n_1155),
.B1(n_1151),
.B2(n_1199),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1156),
.A2(n_1206),
.B1(n_1228),
.B2(n_1199),
.Y(n_1289)
);

AOI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1124),
.A2(n_1104),
.B(n_1210),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1114),
.B(n_1123),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1176),
.A2(n_1204),
.B1(n_1226),
.B2(n_1225),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1114),
.B(n_1170),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1175),
.B(n_1193),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1196),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1211),
.A2(n_1214),
.B1(n_1217),
.B2(n_1218),
.Y(n_1296)
);

OAI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1222),
.A2(n_1229),
.B1(n_1118),
.B2(n_1106),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1103),
.A2(n_956),
.B1(n_985),
.B2(n_911),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1112),
.B(n_1183),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1219),
.A2(n_965),
.B1(n_769),
.B2(n_804),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1219),
.A2(n_1223),
.B1(n_1200),
.B2(n_1208),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1185),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1127),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1111),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1103),
.B(n_1107),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1082),
.B2(n_1096),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1127),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1186),
.A2(n_884),
.B1(n_790),
.B2(n_804),
.Y(n_1308)
);

BUFx4_ASAP7_75t_SL g1309 ( 
.A(n_1187),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1082),
.B2(n_1096),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1219),
.A2(n_1223),
.B1(n_1200),
.B2(n_1208),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1219),
.A2(n_1223),
.B1(n_1200),
.B2(n_1208),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1111),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1082),
.B2(n_1096),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1082),
.B2(n_1096),
.Y(n_1315)
);

OAI22x1_ASAP7_75t_L g1316 ( 
.A1(n_1219),
.A2(n_1082),
.B1(n_1096),
.B2(n_1090),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1082),
.B2(n_1096),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1127),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1200),
.A2(n_911),
.B1(n_790),
.B2(n_804),
.Y(n_1319)
);

BUFx2_ASAP7_75t_SL g1320 ( 
.A(n_1147),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1103),
.A2(n_956),
.B1(n_985),
.B2(n_911),
.Y(n_1321)
);

BUFx8_ASAP7_75t_L g1322 ( 
.A(n_1147),
.Y(n_1322)
);

INVx8_ASAP7_75t_L g1323 ( 
.A(n_1147),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1179),
.A2(n_1110),
.B1(n_1082),
.B2(n_1096),
.Y(n_1324)
);

CKINVDCx14_ASAP7_75t_R g1325 ( 
.A(n_1187),
.Y(n_1325)
);

BUFx12f_ASAP7_75t_L g1326 ( 
.A(n_1127),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1129),
.B(n_1138),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1127),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_1205),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1185),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1200),
.A2(n_911),
.B1(n_790),
.B2(n_804),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1127),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1103),
.A2(n_956),
.B1(n_985),
.B2(n_911),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1219),
.A2(n_965),
.B1(n_769),
.B2(n_804),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1306),
.A2(n_1317),
.B1(n_1315),
.B2(n_1310),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1235),
.Y(n_1336)
);

NOR2x1_ASAP7_75t_SL g1337 ( 
.A(n_1277),
.B(n_1278),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1306),
.B(n_1310),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1319),
.A2(n_1331),
.B(n_1300),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1235),
.Y(n_1340)
);

BUFx8_ASAP7_75t_SL g1341 ( 
.A(n_1307),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1295),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1279),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1297),
.A2(n_1292),
.B(n_1290),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1284),
.A2(n_1296),
.B(n_1294),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1246),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1314),
.B(n_1315),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1286),
.B(n_1236),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1291),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1259),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1259),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1323),
.Y(n_1352)
);

CKINVDCx8_ASAP7_75t_R g1353 ( 
.A(n_1241),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1314),
.B(n_1317),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1308),
.B(n_1255),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1297),
.A2(n_1292),
.B(n_1293),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1289),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1289),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1288),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1324),
.B(n_1233),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1280),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1286),
.B(n_1238),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1236),
.B(n_1247),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1267),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1247),
.B(n_1234),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1276),
.B(n_1245),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1309),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1260),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1267),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1329),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1323),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1253),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1282),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1285),
.B(n_1272),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1273),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1301),
.A2(n_1311),
.B(n_1312),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1284),
.A2(n_1296),
.B(n_1276),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1243),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1274),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1316),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1301),
.A2(n_1312),
.B(n_1311),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1302),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1324),
.A2(n_1233),
.B1(n_1242),
.B2(n_1321),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1256),
.A2(n_1252),
.B(n_1244),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1299),
.B(n_1287),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1265),
.Y(n_1387)
);

AOI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1298),
.A2(n_1333),
.B(n_1263),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1323),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1275),
.A2(n_1334),
.B(n_1330),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1281),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1269),
.A2(n_1264),
.B(n_1305),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1269),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1257),
.A2(n_1249),
.B1(n_1237),
.B2(n_1240),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1270),
.A2(n_1327),
.B(n_1258),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1271),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1251),
.B(n_1313),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1339),
.A2(n_1385),
.B(n_1384),
.C(n_1383),
.Y(n_1398)
);

AO32x2_ASAP7_75t_L g1399 ( 
.A1(n_1343),
.A2(n_1304),
.A3(n_1266),
.B1(n_1254),
.B2(n_1261),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1361),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1341),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1380),
.B(n_1254),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1386),
.B(n_1239),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1383),
.A2(n_1283),
.B1(n_1268),
.B2(n_1318),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1385),
.B(n_1374),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1386),
.B(n_1250),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1373),
.B(n_1320),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_L g1408 ( 
.A(n_1335),
.B(n_1262),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1384),
.B(n_1322),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1384),
.A2(n_1335),
.B1(n_1376),
.B2(n_1381),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1387),
.A2(n_1328),
.B1(n_1325),
.B2(n_1326),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_R g1412 ( 
.A(n_1395),
.B(n_1322),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1385),
.A2(n_1325),
.B(n_1332),
.Y(n_1413)
);

AO21x1_ASAP7_75t_L g1414 ( 
.A1(n_1392),
.A2(n_1303),
.B(n_1374),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1368),
.B(n_1375),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1359),
.B(n_1395),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1376),
.A2(n_1381),
.B1(n_1365),
.B2(n_1360),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1392),
.A2(n_1347),
.B(n_1354),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1337),
.A2(n_1345),
.B(n_1344),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1372),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1365),
.A2(n_1366),
.B(n_1363),
.C(n_1360),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1346),
.B(n_1370),
.Y(n_1423)
);

OAI211xp5_ASAP7_75t_L g1424 ( 
.A1(n_1394),
.A2(n_1387),
.B(n_1365),
.C(n_1338),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1340),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1370),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1350),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1388),
.A2(n_1355),
.B(n_1377),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1351),
.Y(n_1430)
);

AND2x6_ASAP7_75t_L g1431 ( 
.A(n_1366),
.B(n_1363),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1394),
.B(n_1342),
.Y(n_1432)
);

OR2x6_ASAP7_75t_L g1433 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1362),
.A2(n_1377),
.B(n_1348),
.C(n_1393),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1342),
.B(n_1388),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1391),
.A2(n_1374),
.B(n_1345),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1379),
.B(n_1362),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1345),
.A2(n_1358),
.B(n_1357),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1367),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1378),
.B(n_1382),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1342),
.B(n_1390),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1378),
.B(n_1382),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1433),
.B(n_1356),
.Y(n_1444)
);

BUFx2_ASAP7_75t_SL g1445 ( 
.A(n_1431),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1427),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1417),
.B(n_1379),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1433),
.B(n_1420),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1414),
.B(n_1369),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1428),
.B(n_1356),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_1431),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1436),
.B(n_1344),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1430),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1405),
.B(n_1349),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1399),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1410),
.A2(n_1362),
.B1(n_1348),
.B2(n_1353),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1431),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1435),
.B(n_1364),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1439),
.B(n_1336),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1439),
.B(n_1349),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1437),
.B(n_1419),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1441),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1443),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1400),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1400),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1364),
.Y(n_1466)
);

OAI211xp5_ASAP7_75t_L g1467 ( 
.A1(n_1447),
.A2(n_1424),
.B(n_1398),
.C(n_1418),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1460),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1462),
.B(n_1434),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1448),
.B(n_1442),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1462),
.B(n_1434),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1455),
.B(n_1423),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1458),
.B(n_1402),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1448),
.B(n_1416),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1446),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1462),
.B(n_1426),
.Y(n_1476)
);

INVx5_ASAP7_75t_L g1477 ( 
.A(n_1451),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1448),
.B(n_1429),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1450),
.B(n_1452),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1450),
.B(n_1452),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1463),
.B(n_1425),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1453),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1461),
.Y(n_1483)
);

OAI211xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1447),
.A2(n_1408),
.B(n_1404),
.C(n_1398),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1457),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1455),
.B(n_1425),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1455),
.B(n_1438),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1445),
.B(n_1413),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1459),
.B(n_1415),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1485),
.Y(n_1490)
);

AOI211xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1467),
.A2(n_1408),
.B(n_1456),
.C(n_1432),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1475),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1479),
.B(n_1450),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1480),
.B(n_1450),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1468),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1480),
.B(n_1483),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1469),
.B(n_1463),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1477),
.B(n_1457),
.Y(n_1498)
);

INVxp33_ASAP7_75t_L g1499 ( 
.A(n_1473),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1469),
.B(n_1464),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1471),
.B(n_1464),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1468),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1486),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1471),
.B(n_1464),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1480),
.B(n_1444),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1475),
.Y(n_1506)
);

AND2x4_ASAP7_75t_SL g1507 ( 
.A(n_1488),
.B(n_1454),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1482),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1489),
.B(n_1465),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1486),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1481),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_L g1512 ( 
.A(n_1485),
.B(n_1449),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1485),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1497),
.B(n_1487),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1503),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1503),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1490),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1512),
.B(n_1498),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1512),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1510),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1499),
.B(n_1401),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1495),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1498),
.B(n_1505),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1478),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1495),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1495),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1510),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1497),
.B(n_1481),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1498),
.B(n_1478),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1492),
.Y(n_1530)
);

NOR2x1_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1484),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1495),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1502),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1513),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1513),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1500),
.B(n_1501),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1500),
.B(n_1476),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1492),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1501),
.B(n_1476),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1498),
.B(n_1477),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1502),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1504),
.B(n_1472),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1499),
.B(n_1401),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1506),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1508),
.Y(n_1547)
);

AOI31xp33_ASAP7_75t_L g1548 ( 
.A1(n_1491),
.A2(n_1467),
.A3(n_1409),
.B(n_1432),
.Y(n_1548)
);

INVxp67_ASAP7_75t_SL g1549 ( 
.A(n_1504),
.Y(n_1549)
);

OAI21xp33_ASAP7_75t_L g1550 ( 
.A1(n_1491),
.A2(n_1484),
.B(n_1422),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1496),
.B(n_1477),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1515),
.Y(n_1552)
);

NAND3xp33_ASAP7_75t_L g1553 ( 
.A(n_1550),
.B(n_1456),
.C(n_1422),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1531),
.B(n_1445),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1521),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1531),
.B(n_1511),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1516),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1522),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1550),
.B(n_1548),
.Y(n_1560)
);

INVx5_ASAP7_75t_L g1561 ( 
.A(n_1518),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1516),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1548),
.B(n_1473),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1520),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1520),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1523),
.B(n_1493),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1522),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_L g1568 ( 
.A(n_1551),
.B(n_1541),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1522),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1537),
.B(n_1474),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1523),
.B(n_1493),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1537),
.B(n_1509),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.B(n_1493),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1540),
.B(n_1474),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1519),
.B(n_1409),
.C(n_1411),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1540),
.B(n_1509),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1518),
.B(n_1507),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1527),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1528),
.B(n_1474),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1525),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1525),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1494),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1544),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1527),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1528),
.B(n_1470),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1494),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1557),
.B(n_1536),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1560),
.B(n_1517),
.Y(n_1588)
);

AOI21xp33_ASAP7_75t_L g1589 ( 
.A1(n_1554),
.A2(n_1519),
.B(n_1534),
.Y(n_1589)
);

OAI31xp33_ASAP7_75t_L g1590 ( 
.A1(n_1553),
.A2(n_1551),
.A3(n_1534),
.B(n_1535),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1554),
.B(n_1524),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1556),
.B(n_1549),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1561),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1583),
.B(n_1549),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1572),
.B(n_1536),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1552),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1535),
.Y(n_1598)
);

A2O1A1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1553),
.A2(n_1466),
.B(n_1458),
.C(n_1406),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1575),
.A2(n_1554),
.B(n_1568),
.Y(n_1600)
);

OAI21xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1554),
.A2(n_1529),
.B(n_1524),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1552),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1555),
.Y(n_1603)
);

OAI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1575),
.A2(n_1529),
.B1(n_1514),
.B2(n_1530),
.C(n_1538),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1555),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1577),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1554),
.A2(n_1461),
.B(n_1530),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1561),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_SL g1609 ( 
.A(n_1586),
.B(n_1353),
.C(n_1543),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1558),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1577),
.A2(n_1412),
.B1(n_1507),
.B2(n_1488),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1606),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1613)
);

OAI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1600),
.A2(n_1561),
.B1(n_1412),
.B2(n_1451),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1606),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1610),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1570),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1610),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1597),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1604),
.A2(n_1598),
.B1(n_1589),
.B2(n_1592),
.C(n_1595),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1609),
.A2(n_1577),
.B(n_1586),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1599),
.B(n_1558),
.Y(n_1622)
);

AOI321xp33_ASAP7_75t_L g1623 ( 
.A1(n_1599),
.A2(n_1577),
.A3(n_1578),
.B1(n_1565),
.B2(n_1564),
.C(n_1584),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1606),
.B(n_1562),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1587),
.A2(n_1561),
.B1(n_1451),
.B2(n_1562),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1591),
.Y(n_1626)
);

AOI211xp5_ASAP7_75t_L g1627 ( 
.A1(n_1601),
.A2(n_1565),
.B(n_1578),
.C(n_1564),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1573),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1611),
.A2(n_1584),
.B1(n_1572),
.B2(n_1576),
.C(n_1582),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1593),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1602),
.Y(n_1631)
);

AOI221x1_ASAP7_75t_L g1632 ( 
.A1(n_1612),
.A2(n_1608),
.B1(n_1594),
.B2(n_1605),
.C(n_1603),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1613),
.A2(n_1591),
.B1(n_1608),
.B2(n_1594),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1620),
.A2(n_1613),
.B1(n_1622),
.B2(n_1625),
.C(n_1614),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1626),
.B(n_1587),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1617),
.B(n_1421),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1628),
.B(n_1566),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1628),
.B(n_1566),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1624),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1615),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1630),
.B(n_1596),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1637),
.B(n_1638),
.Y(n_1642)
);

OAI211xp5_ASAP7_75t_L g1643 ( 
.A1(n_1634),
.A2(n_1623),
.B(n_1621),
.C(n_1627),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1633),
.B(n_1630),
.Y(n_1644)
);

AND4x1_ASAP7_75t_L g1645 ( 
.A(n_1636),
.B(n_1631),
.C(n_1619),
.D(n_1616),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1640),
.A2(n_1614),
.B1(n_1629),
.B2(n_1625),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1641),
.A2(n_1618),
.B(n_1607),
.C(n_1596),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1635),
.A2(n_1639),
.B(n_1641),
.Y(n_1648)
);

AOI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1632),
.A2(n_1582),
.B(n_1573),
.C(n_1576),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1637),
.Y(n_1650)
);

NOR4xp25_ASAP7_75t_L g1651 ( 
.A(n_1643),
.B(n_1559),
.C(n_1580),
.D(n_1567),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1650),
.A2(n_1547),
.B1(n_1545),
.B2(n_1546),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1647),
.A2(n_1545),
.B(n_1538),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1644),
.A2(n_1648),
.B1(n_1646),
.B2(n_1649),
.C(n_1650),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1642),
.Y(n_1655)
);

O2A1O1Ixp5_ASAP7_75t_L g1656 ( 
.A1(n_1653),
.A2(n_1581),
.B(n_1569),
.C(n_1580),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1655),
.Y(n_1657)
);

AOI221xp5_ASAP7_75t_L g1658 ( 
.A1(n_1651),
.A2(n_1645),
.B1(n_1559),
.B2(n_1567),
.C(n_1569),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1654),
.A2(n_1581),
.B1(n_1569),
.B2(n_1546),
.C(n_1547),
.Y(n_1659)
);

OAI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1652),
.A2(n_1353),
.B(n_1352),
.C(n_1371),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1654),
.A2(n_1396),
.B(n_1581),
.Y(n_1661)
);

XNOR2xp5_ASAP7_75t_L g1662 ( 
.A(n_1657),
.B(n_1352),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1661),
.Y(n_1663)
);

CKINVDCx12_ASAP7_75t_R g1664 ( 
.A(n_1659),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1656),
.Y(n_1665)
);

XNOR2xp5_ASAP7_75t_L g1666 ( 
.A(n_1658),
.B(n_1352),
.Y(n_1666)
);

OR3x2_ASAP7_75t_L g1667 ( 
.A(n_1663),
.B(n_1660),
.C(n_1440),
.Y(n_1667)
);

OAI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1665),
.A2(n_1371),
.B(n_1396),
.C(n_1389),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1662),
.B(n_1571),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1667),
.A2(n_1666),
.B1(n_1668),
.B2(n_1669),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1670),
.A2(n_1664),
.B1(n_1440),
.B2(n_1571),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1671),
.A2(n_1664),
.B1(n_1389),
.B2(n_1533),
.Y(n_1672)
);

AO211x2_ASAP7_75t_L g1673 ( 
.A1(n_1672),
.A2(n_1585),
.B(n_1514),
.C(n_1407),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1673),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1542),
.B1(n_1525),
.B2(n_1526),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1674),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1574),
.B(n_1579),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1675),
.A2(n_1532),
.B(n_1526),
.Y(n_1678)
);

XOR2xp5_ASAP7_75t_L g1679 ( 
.A(n_1677),
.B(n_1371),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1678),
.A2(n_1526),
.B1(n_1532),
.B2(n_1533),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1679),
.A2(n_1532),
.B1(n_1533),
.B2(n_1539),
.C(n_1542),
.Y(n_1681)
);

AOI211xp5_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1680),
.B(n_1403),
.C(n_1539),
.Y(n_1682)
);


endmodule