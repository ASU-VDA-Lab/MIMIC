module fake_jpeg_20549_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_50),
.Y(n_64)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_42),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_38),
.C(n_45),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_4),
.C(n_5),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_41),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_37),
.B1(n_35),
.B2(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_40),
.B1(n_42),
.B2(n_3),
.Y(n_71)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_1),
.C(n_2),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_79),
.C(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_1),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_86)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_67),
.B1(n_5),
.B2(n_4),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_87),
.B1(n_89),
.B2(n_70),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_93),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_100)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_92),
.B1(n_98),
.B2(n_82),
.C(n_83),
.Y(n_99)
);

XOR2x1_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_20),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_25),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_30),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_33),
.Y(n_108)
);


endmodule