module real_aes_8446_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g113 ( .A(n_0), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_1), .A2(n_150), .B(n_153), .C(n_156), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_2), .A2(n_176), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g536 ( .A(n_3), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_4), .B(n_199), .Y(n_222) );
AOI21xp33_ASAP7_75t_L g463 ( .A1(n_5), .A2(n_176), .B(n_464), .Y(n_463) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g183 ( .A(n_7), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_8), .B(n_41), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_9), .A2(n_230), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_10), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g468 ( .A(n_11), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_12), .B(n_205), .Y(n_507) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
INVx1_ASAP7_75t_L g519 ( .A(n_14), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_15), .A2(n_184), .B(n_194), .C(n_197), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_16), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_17), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_18), .B(n_475), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_19), .B(n_176), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_20), .B(n_240), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_21), .A2(n_205), .B(n_206), .C(n_208), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_22), .B(n_199), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_23), .B(n_162), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_24), .A2(n_196), .B(n_197), .C(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_25), .B(n_162), .Y(n_249) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_26), .Y(n_258) );
INVx1_ASAP7_75t_L g248 ( .A(n_27), .Y(n_248) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_29), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_30), .B(n_162), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_31), .A2(n_65), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_31), .Y(n_127) );
INVx1_ASAP7_75t_L g235 ( .A(n_32), .Y(n_235) );
INVx1_ASAP7_75t_L g457 ( .A(n_33), .Y(n_457) );
INVx2_ASAP7_75t_L g148 ( .A(n_34), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_35), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_36), .A2(n_205), .B(n_218), .C(n_220), .Y(n_217) );
INVxp67_ASAP7_75t_L g237 ( .A(n_37), .Y(n_237) );
CKINVDCx14_ASAP7_75t_R g216 ( .A(n_38), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_39), .A2(n_153), .B(n_247), .C(n_251), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_40), .A2(n_150), .B(n_153), .C(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g456 ( .A(n_42), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_43), .A2(n_164), .B(n_181), .C(n_182), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_44), .B(n_162), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_45), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_46), .Y(n_232) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_47), .A2(n_445), .B1(n_721), .B2(n_724), .C1(n_725), .C2(n_727), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_48), .A2(n_102), .B1(n_115), .B2(n_731), .Y(n_101) );
INVx1_ASAP7_75t_L g203 ( .A(n_49), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g458 ( .A(n_50), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_51), .B(n_176), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_52), .A2(n_153), .B1(n_208), .B2(n_455), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_53), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_54), .Y(n_533) );
CKINVDCx14_ASAP7_75t_R g178 ( .A(n_55), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_56), .A2(n_181), .B(n_220), .C(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_57), .Y(n_499) );
INVx1_ASAP7_75t_L g465 ( .A(n_58), .Y(n_465) );
INVx1_ASAP7_75t_L g151 ( .A(n_59), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_60), .A2(n_78), .B1(n_722), .B2(n_723), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_60), .Y(n_723) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
INVx1_ASAP7_75t_SL g219 ( .A(n_62), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_63), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_64), .B(n_199), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_65), .Y(n_126) );
INVx1_ASAP7_75t_L g261 ( .A(n_66), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_SL g474 ( .A1(n_67), .A2(n_220), .B(n_475), .C(n_476), .Y(n_474) );
INVxp67_ASAP7_75t_L g477 ( .A(n_68), .Y(n_477) );
INVx1_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_70), .A2(n_176), .B(n_177), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_71), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_72), .A2(n_176), .B(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_73), .Y(n_460) );
INVx1_ASAP7_75t_L g493 ( .A(n_74), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_75), .A2(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g192 ( .A(n_76), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_77), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_78), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_79), .A2(n_150), .B(n_153), .C(n_495), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_80), .A2(n_176), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g195 ( .A(n_81), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_82), .B(n_236), .Y(n_487) );
INVx2_ASAP7_75t_L g139 ( .A(n_83), .Y(n_139) );
INVx1_ASAP7_75t_L g157 ( .A(n_84), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_85), .B(n_475), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_86), .A2(n_150), .B(n_153), .C(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g110 ( .A(n_87), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g717 ( .A(n_87), .Y(n_717) );
OR2x2_ASAP7_75t_L g720 ( .A(n_87), .B(n_112), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_88), .A2(n_153), .B(n_260), .C(n_263), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_89), .B(n_138), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_90), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_91), .A2(n_150), .B(n_153), .C(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_92), .Y(n_511) );
INVx1_ASAP7_75t_L g473 ( .A(n_93), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_94), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_95), .B(n_236), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_96), .B(n_169), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_97), .B(n_169), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_98), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g207 ( .A(n_99), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_100), .A2(n_176), .B(n_472), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g732 ( .A(n_105), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g122 ( .A(n_110), .Y(n_122) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_110), .Y(n_442) );
NOR2x2_ASAP7_75t_L g729 ( .A(n_111), .B(n_717), .Y(n_729) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g716 ( .A(n_112), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_443), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g730 ( .A(n_120), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B(n_440), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_128), .B2(n_129), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_128), .A2(n_446), .B1(n_714), .B2(n_718), .Y(n_445) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_129), .A2(n_714), .B1(n_720), .B2(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_395), .Y(n_129) );
NAND5xp2_ASAP7_75t_L g130 ( .A(n_131), .B(n_307), .C(n_345), .D(n_366), .E(n_383), .Y(n_130) );
NOR3xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_279), .C(n_300), .Y(n_131) );
OAI221xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_211), .B1(n_242), .B2(n_266), .C(n_270), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_171), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_135), .B(n_268), .Y(n_287) );
OR2x2_ASAP7_75t_L g314 ( .A(n_135), .B(n_188), .Y(n_314) );
AND2x2_ASAP7_75t_L g328 ( .A(n_135), .B(n_188), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_135), .B(n_174), .Y(n_342) );
AND2x2_ASAP7_75t_L g380 ( .A(n_135), .B(n_344), .Y(n_380) );
AND2x2_ASAP7_75t_L g409 ( .A(n_135), .B(n_319), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_135), .B(n_291), .Y(n_426) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g306 ( .A(n_136), .B(n_187), .Y(n_306) );
BUFx3_ASAP7_75t_L g331 ( .A(n_136), .Y(n_331) );
AND2x2_ASAP7_75t_L g360 ( .A(n_136), .B(n_188), .Y(n_360) );
AND3x2_ASAP7_75t_L g373 ( .A(n_136), .B(n_374), .C(n_375), .Y(n_373) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_166), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_137), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_137), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_137), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_138), .A2(n_175), .B(n_186), .Y(n_174) );
INVx2_ASAP7_75t_L g241 ( .A(n_138), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_138), .A2(n_145), .B(n_245), .C(n_246), .Y(n_244) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_138), .A2(n_514), .B(n_520), .Y(n_513) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_L g170 ( .A(n_139), .B(n_140), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_152), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_145), .A2(n_258), .B(n_259), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g453 ( .A1(n_145), .A2(n_185), .B1(n_454), .B2(n_458), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_145), .A2(n_493), .B(n_494), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_145), .A2(n_533), .B(n_534), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
AND2x4_ASAP7_75t_L g176 ( .A(n_146), .B(n_150), .Y(n_176) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g238 ( .A(n_147), .Y(n_238) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
INVx3_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
INVx1_ASAP7_75t_L g475 ( .A(n_149), .Y(n_475) );
INVx4_ASAP7_75t_SL g185 ( .A(n_150), .Y(n_185) );
BUFx3_ASAP7_75t_L g251 ( .A(n_150), .Y(n_251) );
INVx5_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx3_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_154), .Y(n_221) );
O2A1O1Ixp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_161), .C(n_163), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g260 ( .A1(n_158), .A2(n_163), .B(n_261), .C(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_159), .A2(n_160), .B1(n_456), .B2(n_457), .Y(n_455) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx4_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
INVx2_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
INVx4_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_163), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_163), .A2(n_496), .B(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g197 ( .A(n_165), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx3_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_168), .B(n_253), .Y(n_252) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_168), .A2(n_257), .B(n_264), .Y(n_256) );
NOR2xp33_ASAP7_75t_SL g489 ( .A(n_168), .B(n_490), .Y(n_489) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_169), .Y(n_189) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_169), .A2(n_471), .B(n_478), .Y(n_470) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
INVx1_ASAP7_75t_L g296 ( .A(n_171), .Y(n_296) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_187), .Y(n_171) );
AOI32xp33_ASAP7_75t_L g351 ( .A1(n_172), .A2(n_303), .A3(n_352), .B1(n_355), .B2(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g278 ( .A(n_173), .B(n_187), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_173), .B(n_306), .Y(n_349) );
AND2x2_ASAP7_75t_L g356 ( .A(n_173), .B(n_328), .Y(n_356) );
OR2x2_ASAP7_75t_L g362 ( .A(n_173), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_173), .B(n_317), .Y(n_387) );
OR2x2_ASAP7_75t_L g405 ( .A(n_173), .B(n_224), .Y(n_405) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g269 ( .A(n_174), .B(n_200), .Y(n_269) );
INVx2_ASAP7_75t_L g291 ( .A(n_174), .Y(n_291) );
OR2x2_ASAP7_75t_L g313 ( .A(n_174), .B(n_200), .Y(n_313) );
AND2x2_ASAP7_75t_L g318 ( .A(n_174), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_174), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g374 ( .A(n_174), .B(n_268), .Y(n_374) );
BUFx2_ASAP7_75t_L g230 ( .A(n_176), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B(n_180), .C(n_185), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g191 ( .A1(n_179), .A2(n_185), .B(n_192), .C(n_193), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_SL g202 ( .A1(n_179), .A2(n_185), .B(n_203), .C(n_204), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_179), .A2(n_185), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_179), .A2(n_185), .B(n_232), .C(n_233), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_179), .A2(n_185), .B(n_465), .C(n_466), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_179), .A2(n_185), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_179), .A2(n_185), .B(n_516), .C(n_517), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
INVx5_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_184), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_184), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g263 ( .A(n_185), .Y(n_263) );
INVx1_ASAP7_75t_SL g425 ( .A(n_187), .Y(n_425) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_200), .Y(n_187) );
INVx1_ASAP7_75t_SL g268 ( .A(n_188), .Y(n_268) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_188), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_188), .B(n_354), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_188), .B(n_291), .C(n_409), .Y(n_420) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_198), .Y(n_188) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_189), .A2(n_201), .B(n_210), .Y(n_200) );
OA21x2_ASAP7_75t_L g213 ( .A1(n_189), .A2(n_214), .B(n_222), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_196), .B(n_207), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_196), .A2(n_235), .B1(n_236), .B2(n_237), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_196), .B(n_519), .Y(n_518) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_199), .A2(n_463), .B(n_469), .Y(n_462) );
INVx2_ASAP7_75t_L g319 ( .A(n_200), .Y(n_319) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_200), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_205), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g538 ( .A(n_208), .Y(n_538) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
INVx1_ASAP7_75t_L g355 ( .A(n_212), .Y(n_355) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g273 ( .A(n_213), .B(n_255), .Y(n_273) );
INVx2_ASAP7_75t_L g290 ( .A(n_213), .Y(n_290) );
AND2x2_ASAP7_75t_L g295 ( .A(n_213), .B(n_256), .Y(n_295) );
AND2x2_ASAP7_75t_L g310 ( .A(n_213), .B(n_243), .Y(n_310) );
AND2x2_ASAP7_75t_L g322 ( .A(n_213), .B(n_294), .Y(n_322) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_221), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_223), .B(n_338), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g394 ( .A(n_223), .B(n_295), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_223), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_223), .B(n_289), .Y(n_417) );
BUFx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g254 ( .A(n_224), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_224), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g299 ( .A(n_224), .B(n_243), .Y(n_299) );
AND2x2_ASAP7_75t_L g325 ( .A(n_224), .B(n_255), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_224), .B(n_365), .Y(n_364) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_229), .B(n_239), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_226), .A2(n_284), .B(n_285), .Y(n_283) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_226), .A2(n_492), .B(n_498), .Y(n_491) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_SL g483 ( .A1(n_227), .A2(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_228), .A2(n_453), .B(n_459), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_228), .B(n_460), .Y(n_459) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_228), .A2(n_532), .B(n_539), .Y(n_531) );
INVx1_ASAP7_75t_L g284 ( .A(n_229), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_234), .B(n_238), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_236), .A2(n_248), .B(n_249), .C(n_250), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_236), .A2(n_536), .B(n_537), .C(n_538), .Y(n_535) );
INVx2_ASAP7_75t_L g250 ( .A(n_238), .Y(n_250) );
INVx1_ASAP7_75t_L g285 ( .A(n_239), .Y(n_285) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_241), .B(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_241), .A2(n_503), .B(n_510), .Y(n_502) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_254), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_243), .B(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g289 ( .A(n_243), .B(n_290), .Y(n_289) );
INVx3_ASAP7_75t_SL g294 ( .A(n_243), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_243), .B(n_281), .Y(n_347) );
OR2x2_ASAP7_75t_L g357 ( .A(n_243), .B(n_283), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_243), .B(n_325), .Y(n_385) );
OR2x2_ASAP7_75t_L g415 ( .A(n_243), .B(n_255), .Y(n_415) );
AND2x2_ASAP7_75t_L g419 ( .A(n_243), .B(n_256), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_243), .B(n_295), .Y(n_432) );
AND2x2_ASAP7_75t_L g439 ( .A(n_243), .B(n_321), .Y(n_439) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_252), .Y(n_243) );
INVx1_ASAP7_75t_SL g382 ( .A(n_254), .Y(n_382) );
AND2x2_ASAP7_75t_L g321 ( .A(n_255), .B(n_283), .Y(n_321) );
AND2x2_ASAP7_75t_L g335 ( .A(n_255), .B(n_290), .Y(n_335) );
AND2x2_ASAP7_75t_L g338 ( .A(n_255), .B(n_294), .Y(n_338) );
INVx1_ASAP7_75t_L g365 ( .A(n_255), .Y(n_365) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
BUFx2_ASAP7_75t_L g277 ( .A(n_256), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g436 ( .A1(n_267), .A2(n_313), .B(n_437), .C(n_438), .Y(n_436) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g343 ( .A(n_268), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_269), .B(n_286), .Y(n_301) );
AND2x2_ASAP7_75t_L g327 ( .A(n_269), .B(n_328), .Y(n_327) );
OAI21xp5_ASAP7_75t_SL g270 ( .A1(n_271), .A2(n_274), .B(n_278), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_272), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g298 ( .A(n_273), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_273), .B(n_294), .Y(n_339) );
AND2x2_ASAP7_75t_L g430 ( .A(n_273), .B(n_281), .Y(n_430) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g303 ( .A(n_277), .B(n_290), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_288), .Y(n_304) );
OAI322xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_287), .A3(n_288), .B1(n_291), .B2(n_292), .C1(n_296), .C2(n_297), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_286), .Y(n_280) );
AND2x2_ASAP7_75t_L g391 ( .A(n_281), .B(n_303), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_281), .B(n_355), .Y(n_437) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g334 ( .A(n_283), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g400 ( .A(n_287), .B(n_313), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_288), .B(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_289), .B(n_321), .Y(n_378) );
AND2x2_ASAP7_75t_L g324 ( .A(n_290), .B(n_294), .Y(n_324) );
AND2x2_ASAP7_75t_L g332 ( .A(n_291), .B(n_333), .Y(n_332) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_291), .A2(n_370), .B(n_430), .C(n_431), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_292), .A2(n_305), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_294), .B(n_321), .Y(n_361) );
AND2x2_ASAP7_75t_L g367 ( .A(n_294), .B(n_335), .Y(n_367) );
AND2x2_ASAP7_75t_L g401 ( .A(n_294), .B(n_303), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_295), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_SL g411 ( .A(n_295), .Y(n_411) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_299), .A2(n_327), .B1(n_329), .B2(n_334), .Y(n_326) );
OAI22xp5_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_302), .B1(n_304), .B2(n_305), .Y(n_300) );
OAI22xp33_ASAP7_75t_L g336 ( .A1(n_301), .A2(n_337), .B1(n_339), .B2(n_340), .Y(n_336) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_306), .A2(n_408), .B1(n_410), .B2(n_412), .C(n_416), .Y(n_407) );
AOI211xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B(n_315), .C(n_336), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
OR2x2_ASAP7_75t_L g377 ( .A(n_313), .B(n_330), .Y(n_377) );
INVx1_ASAP7_75t_L g428 ( .A(n_313), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_314), .A2(n_316), .B1(n_320), .B2(n_323), .C(n_326), .Y(n_315) );
INVx2_ASAP7_75t_SL g370 ( .A(n_314), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g435 ( .A(n_317), .Y(n_435) );
AND2x2_ASAP7_75t_L g359 ( .A(n_318), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g344 ( .A(n_319), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g406 ( .A(n_322), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_330), .B(n_432), .Y(n_431) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_331), .Y(n_330) );
INVxp67_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g345 ( .A1(n_334), .A2(n_346), .B(n_348), .C(n_350), .Y(n_345) );
INVx1_ASAP7_75t_L g423 ( .A(n_337), .Y(n_423) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_341), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx2_ASAP7_75t_L g354 ( .A(n_344), .Y(n_354) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI222xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_357), .B1(n_358), .B2(n_361), .C1(n_362), .C2(n_364), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g390 ( .A(n_354), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_357), .B(n_411), .Y(n_410) );
NAND2xp33_ASAP7_75t_SL g388 ( .A(n_358), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g363 ( .A(n_360), .Y(n_363) );
AND2x2_ASAP7_75t_L g427 ( .A(n_360), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g393 ( .A(n_363), .B(n_390), .Y(n_393) );
INVx1_ASAP7_75t_L g422 ( .A(n_364), .Y(n_422) );
AOI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B(n_371), .C(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_370), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_373), .A2(n_401), .A3(n_406), .B1(n_422), .B2(n_423), .C1(n_424), .C2(n_427), .Y(n_421) );
AND2x2_ASAP7_75t_L g408 ( .A(n_374), .B(n_409), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B1(n_379), .B2(n_381), .Y(n_376) );
INVxp33_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B1(n_388), .B2(n_391), .C(n_392), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
NAND5xp2_ASAP7_75t_L g395 ( .A(n_396), .B(n_407), .C(n_421), .D(n_429), .E(n_433), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_401), .B(n_402), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp33_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_409), .A2(n_434), .B(n_435), .C(n_436), .Y(n_433) );
AOI31xp33_ASAP7_75t_L g416 ( .A1(n_411), .A2(n_417), .A3(n_418), .B(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g434 ( .A(n_432), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_440), .B(n_444), .C(n_730), .Y(n_443) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g726 ( .A(n_446), .Y(n_726) );
AND3x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_639), .C(n_688), .Y(n_446) );
NOR3xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_546), .C(n_584), .Y(n_447) );
OAI222xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_479), .B1(n_521), .B2(n_527), .C1(n_541), .C2(n_544), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_461), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_450), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_450), .B(n_589), .Y(n_680) );
BUFx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g557 ( .A(n_451), .B(n_470), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_451), .B(n_462), .Y(n_565) );
AND2x2_ASAP7_75t_L g600 ( .A(n_451), .B(n_577), .Y(n_600) );
OR2x2_ASAP7_75t_L g624 ( .A(n_451), .B(n_462), .Y(n_624) );
OR2x2_ASAP7_75t_L g632 ( .A(n_451), .B(n_531), .Y(n_632) );
AND2x2_ASAP7_75t_L g635 ( .A(n_451), .B(n_470), .Y(n_635) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g529 ( .A(n_452), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g543 ( .A(n_452), .B(n_470), .Y(n_543) );
AND2x2_ASAP7_75t_L g593 ( .A(n_452), .B(n_531), .Y(n_593) );
AND2x2_ASAP7_75t_L g606 ( .A(n_452), .B(n_462), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_452), .B(n_692), .Y(n_713) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_461), .A2(n_632), .B(n_633), .C(n_636), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_461), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_461), .B(n_576), .Y(n_698) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_470), .Y(n_461) );
AND2x2_ASAP7_75t_SL g542 ( .A(n_462), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g556 ( .A(n_462), .Y(n_556) );
AND2x2_ASAP7_75t_L g583 ( .A(n_462), .B(n_577), .Y(n_583) );
INVx1_ASAP7_75t_SL g591 ( .A(n_462), .Y(n_591) );
AND2x2_ASAP7_75t_L g614 ( .A(n_462), .B(n_615), .Y(n_614) );
BUFx2_ASAP7_75t_L g692 ( .A(n_462), .Y(n_692) );
BUFx2_ASAP7_75t_L g528 ( .A(n_470), .Y(n_528) );
INVx1_ASAP7_75t_L g590 ( .A(n_470), .Y(n_590) );
INVx3_ASAP7_75t_L g615 ( .A(n_470), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_479), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_500), .Y(n_479) );
INVx1_ASAP7_75t_L g611 ( .A(n_480), .Y(n_611) );
OAI32xp33_ASAP7_75t_L g617 ( .A1(n_480), .A2(n_556), .A3(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_480), .A2(n_622), .B1(n_625), .B2(n_630), .Y(n_621) );
INVx4_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g559 ( .A(n_481), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g637 ( .A(n_481), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g707 ( .A(n_481), .B(n_653), .Y(n_707) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_491), .Y(n_481) );
AND2x2_ASAP7_75t_L g522 ( .A(n_482), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g552 ( .A(n_482), .Y(n_552) );
INVx1_ASAP7_75t_L g571 ( .A(n_482), .Y(n_571) );
OR2x2_ASAP7_75t_L g579 ( .A(n_482), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g586 ( .A(n_482), .B(n_560), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_482), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g607 ( .A(n_482), .B(n_525), .Y(n_607) );
INVx3_ASAP7_75t_L g629 ( .A(n_482), .Y(n_629) );
AND2x2_ASAP7_75t_L g654 ( .A(n_482), .B(n_526), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_482), .B(n_619), .Y(n_702) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .Y(n_482) );
INVx2_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
AND2x2_ASAP7_75t_L g658 ( .A(n_491), .B(n_501), .Y(n_658) );
INVx2_ASAP7_75t_L g700 ( .A(n_500), .Y(n_700) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
INVx1_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
AND2x2_ASAP7_75t_L g572 ( .A(n_501), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_501), .B(n_526), .Y(n_580) );
AND2x2_ASAP7_75t_L g638 ( .A(n_501), .B(n_561), .Y(n_638) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g524 ( .A(n_502), .Y(n_524) );
AND2x2_ASAP7_75t_L g551 ( .A(n_502), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g560 ( .A(n_502), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_502), .B(n_526), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B(n_508), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_512), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g573 ( .A(n_512), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_512), .B(n_526), .Y(n_619) );
AND2x2_ASAP7_75t_L g628 ( .A(n_512), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g653 ( .A(n_512), .Y(n_653) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g525 ( .A(n_513), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g561 ( .A(n_513), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_521), .A2(n_531), .B1(n_690), .B2(n_693), .Y(n_689) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
OAI21xp5_ASAP7_75t_SL g712 ( .A1(n_523), .A2(n_634), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_524), .B(n_629), .Y(n_646) );
INVx1_ASAP7_75t_L g671 ( .A(n_524), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_525), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g598 ( .A(n_525), .B(n_551), .Y(n_598) );
INVx2_ASAP7_75t_L g554 ( .A(n_526), .Y(n_554) );
INVx1_ASAP7_75t_L g604 ( .A(n_526), .Y(n_604) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_527), .A2(n_679), .B1(n_696), .B2(n_699), .C(n_701), .Y(n_695) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g566 ( .A(n_528), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_528), .B(n_577), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_529), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g620 ( .A(n_529), .B(n_566), .Y(n_620) );
INVx3_ASAP7_75t_SL g661 ( .A(n_529), .Y(n_661) );
AND2x2_ASAP7_75t_L g605 ( .A(n_530), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g634 ( .A(n_530), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_530), .B(n_543), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_530), .B(n_589), .Y(n_675) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g577 ( .A(n_531), .Y(n_577) );
OAI322xp33_ASAP7_75t_L g672 ( .A1(n_531), .A2(n_603), .A3(n_625), .B1(n_673), .B2(n_675), .C1(n_676), .C2(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_542), .A2(n_545), .B(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_SL g622 ( .A(n_543), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g644 ( .A(n_543), .B(n_556), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_543), .B(n_583), .Y(n_659) );
INVxp67_ASAP7_75t_L g610 ( .A(n_545), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g616 ( .A1(n_545), .A2(n_617), .B(n_621), .C(n_631), .Y(n_616) );
OAI221xp5_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_555), .B1(n_558), .B2(n_562), .C(n_567), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g570 ( .A(n_554), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g687 ( .A(n_554), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_555), .A2(n_704), .B1(n_709), .B2(n_710), .C(n_712), .Y(n_703) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_556), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g603 ( .A(n_556), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_556), .B(n_634), .Y(n_641) );
AND2x2_ASAP7_75t_L g683 ( .A(n_556), .B(n_661), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_557), .B(n_582), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g678 ( .A1(n_557), .A2(n_569), .B1(n_679), .B2(n_680), .Y(n_678) );
OR2x2_ASAP7_75t_L g709 ( .A(n_557), .B(n_577), .Y(n_709) );
CKINVDCx16_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g686 ( .A(n_560), .Y(n_686) );
AND2x2_ASAP7_75t_L g711 ( .A(n_560), .B(n_654), .Y(n_711) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_SL g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g575 ( .A(n_565), .B(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_574), .B1(n_578), .B2(n_581), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx1_ASAP7_75t_L g642 ( .A(n_570), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_570), .B(n_610), .Y(n_677) );
AOI322xp5_ASAP7_75t_L g601 ( .A1(n_572), .A2(n_602), .A3(n_604), .B1(n_605), .B2(n_607), .C1(n_608), .C2(n_612), .Y(n_601) );
INVxp67_ASAP7_75t_L g595 ( .A(n_573), .Y(n_595) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_575), .A2(n_580), .B1(n_597), .B2(n_599), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_576), .B(n_589), .Y(n_676) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_577), .B(n_615), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_577), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g673 ( .A(n_579), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
NAND3xp33_ASAP7_75t_SL g584 ( .A(n_585), .B(n_601), .C(n_616), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_592), .B2(n_594), .C(n_596), .Y(n_585) );
AND2x2_ASAP7_75t_L g592 ( .A(n_588), .B(n_593), .Y(n_592) );
INVx3_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g602 ( .A(n_593), .B(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_595), .Y(n_674) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_600), .B(n_614), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_603), .B(n_661), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_604), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g679 ( .A(n_607), .Y(n_679) );
AND2x2_ASAP7_75t_L g694 ( .A(n_607), .B(n_671), .Y(n_694) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_618), .A2(n_689), .B(n_695), .C(n_703), .Y(n_688) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g657 ( .A(n_628), .B(n_658), .Y(n_657) );
NAND2x1_ASAP7_75t_SL g699 ( .A(n_629), .B(n_700), .Y(n_699) );
CKINVDCx16_ASAP7_75t_R g669 ( .A(n_632), .Y(n_669) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g664 ( .A(n_638), .Y(n_664) );
AND2x2_ASAP7_75t_L g668 ( .A(n_638), .B(n_654), .Y(n_668) );
NOR5xp2_ASAP7_75t_L g639 ( .A(n_640), .B(n_655), .C(n_672), .D(n_678), .E(n_681), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_645), .C(n_647), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_644), .B(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g670 ( .A(n_654), .B(n_671), .Y(n_670) );
OAI221xp5_ASAP7_75t_SL g655 ( .A1(n_656), .A2(n_659), .B1(n_660), .B2(n_662), .C(n_665), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g708 ( .A(n_668), .Y(n_708) );
AOI211xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_684), .B(n_686), .C(n_687), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
CKINVDCx14_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx14_ASAP7_75t_R g724 ( .A(n_721), .Y(n_724) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx3_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
endmodule