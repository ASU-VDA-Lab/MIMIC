module fake_jpeg_17649_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_0),
.C(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_39),
.B(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_42),
.B(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_1),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_49),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_21),
.A2(n_3),
.B(n_5),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_58),
.B(n_10),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_3),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_60),
.Y(n_75)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_21),
.B(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_24),
.B(n_6),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_25),
.B(n_7),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_11),
.Y(n_97)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_20),
.B1(n_37),
.B2(n_29),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_70),
.B1(n_73),
.B2(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_20),
.B1(n_37),
.B2(n_29),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_98),
.B1(n_99),
.B2(n_83),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_74),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_36),
.B1(n_31),
.B2(n_22),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_25),
.B1(n_35),
.B2(n_28),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_36),
.B(n_31),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_92),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_35),
.B1(n_28),
.B2(n_27),
.Y(n_84)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_27),
.B1(n_36),
.B2(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_95),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_38),
.A2(n_36),
.B1(n_27),
.B2(n_22),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_27),
.B1(n_12),
.B2(n_11),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_88),
.B1(n_69),
.B2(n_66),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_77),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_12),
.B1(n_19),
.B2(n_56),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_41),
.A2(n_19),
.B1(n_20),
.B2(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_19),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_105),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_72),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_107),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_99),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_110),
.A2(n_124),
.B(n_64),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_80),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_114),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_79),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_78),
.B(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_68),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_104),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_85),
.C(n_89),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_145),
.C(n_149),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_66),
.B1(n_64),
.B2(n_63),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_147),
.B1(n_146),
.B2(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_124),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_89),
.Y(n_144)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_146),
.B1(n_116),
.B2(n_124),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_64),
.B(n_89),
.Y(n_145)
);

AO22x2_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_64),
.B1(n_93),
.B2(n_123),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_125),
.B1(n_117),
.B2(n_101),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_111),
.C(n_105),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_170),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_167),
.B(n_175),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_172),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_125),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_161),
.C(n_168),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_111),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_106),
.C(n_102),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_113),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_173),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_139),
.B1(n_146),
.B2(n_153),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_186),
.B1(n_189),
.B2(n_169),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_154),
.C(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.C(n_188),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_146),
.C(n_132),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_146),
.B(n_137),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_189),
.B(n_139),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_179),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_132),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_145),
.B(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_192),
.Y(n_203)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_167),
.B(n_159),
.C(n_130),
.D(n_168),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_166),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_170),
.C(n_137),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_182),
.C(n_188),
.Y(n_198)
);

AO221x1_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_156),
.B1(n_163),
.B2(n_165),
.C(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_143),
.C(n_174),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_184),
.C(n_102),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_209),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_194),
.C(n_193),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_158),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_193),
.C(n_198),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_112),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_203),
.B(n_208),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_217),
.A3(n_218),
.B1(n_202),
.B2(n_215),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_220),
.A2(n_219),
.B(n_109),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_108),
.Y(n_222)
);


endmodule