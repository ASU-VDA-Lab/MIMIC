module fake_jpeg_32147_n_97 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_97);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_1),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_0),
.B1(n_7),
.B2(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_35),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_14),
.B(n_22),
.C(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_52),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_33),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_16),
.Y(n_45)
);

NOR2x1p5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_27),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_54),
.B(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_31),
.C(n_30),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_53),
.C(n_8),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_32),
.A2(n_30),
.B1(n_27),
.B2(n_13),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_19),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_24),
.B(n_19),
.C(n_13),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_52),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_46),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_48),
.B1(n_41),
.B2(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_10),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_79),
.C(n_62),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_55),
.C(n_64),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_70),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_88),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_90),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g96 ( 
.A(n_95),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_93),
.Y(n_97)
);


endmodule