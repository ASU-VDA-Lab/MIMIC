module real_jpeg_5498_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_45),
.B1(n_76),
.B2(n_80),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_45),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_45),
.B1(n_174),
.B2(n_176),
.Y(n_210)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_3),
.A2(n_21),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_6),
.Y(n_160)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_8),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_10),
.A2(n_54),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_10),
.A2(n_54),
.B1(n_70),
.B2(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_10),
.B(n_132),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_10),
.A2(n_254),
.B(n_256),
.C(n_264),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_10),
.B(n_281),
.C(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_10),
.B(n_83),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_10),
.B(n_154),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_10),
.B(n_68),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_11),
.A2(n_118),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_11),
.A2(n_139),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_11),
.A2(n_51),
.B1(n_139),
.B2(n_260),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_11),
.A2(n_139),
.B1(n_291),
.B2(n_295),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_221),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_219),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_198),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_16),
.B(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.C(n_177),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_17),
.B(n_177),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_81),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_18),
.B(n_115),
.C(n_144),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_19),
.B(n_47),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_30),
.B(n_37),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_20),
.A2(n_152),
.B(n_155),
.Y(n_151)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_31),
.B(n_40),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_31),
.A2(n_181),
.B(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_31),
.B(n_184),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_31),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_32),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_33),
.Y(n_294)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_37),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_37),
.B(n_289),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_44),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_44),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_74),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_48),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_52),
.Y(n_196)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_53),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_54),
.B(n_120),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_54),
.A2(n_165),
.B(n_207),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_54),
.A2(n_257),
.B(n_260),
.Y(n_256)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_56),
.B(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_56),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_56),
.B(n_271),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_64),
.Y(n_282)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_68),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_68),
.B(n_271),
.Y(n_285)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_74),
.A2(n_190),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_74),
.B(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_79),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_115),
.B1(n_144),
.B2(n_145),
.Y(n_81)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_95),
.B(n_109),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_83),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_83),
.B(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_91),
.B2(n_93),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_87),
.Y(n_259)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_92),
.Y(n_192)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_95),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_95),
.B(n_109),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_96),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_99),
.Y(n_255)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_109),
.Y(n_171)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_114),
.Y(n_265)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_137),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_132),
.Y(n_148)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_122),
.B(n_206),
.Y(n_237)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_132),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_132),
.B(n_206),
.Y(n_205)
);

AO22x1_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_137),
.B(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_146),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_168),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_147),
.B(n_168),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_149),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_150),
.B(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_151),
.B(n_156),
.Y(n_234)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_154),
.Y(n_308)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.A3(n_161),
.B1(n_164),
.B2(n_166),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_209),
.Y(n_228)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_187),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_179),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_187),
.B(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B(n_197),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_216),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_189),
.B(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_197),
.B(n_285),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_198),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_212),
.CI(n_218),
.CON(n_198),
.SN(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_211),
.B(n_243),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_213),
.A2(n_217),
.B1(n_253),
.B2(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_339),
.B(n_350),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_272),
.B(n_338),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_248),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_224),
.B(n_248),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_227),
.B(n_233),
.C(n_235),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_232),
.B(n_307),
.Y(n_315)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_236),
.B(n_239),
.C(n_245),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_266),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_249),
.B(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_252),
.A2(n_266),
.B1(n_267),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_332),
.B(n_337),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_322),
.B(n_331),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_301),
.B(n_321),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_286),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_284),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_278),
.B1(n_284),
.B2(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_308),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_299),
.C(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_309),
.B(n_320),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_305),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_316),
.B(n_319),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_325),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_336),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_336),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_347),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_342),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_342),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_348),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.CI(n_345),
.CON(n_342),
.SN(n_342)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_351),
.B(n_352),
.Y(n_350)
);


endmodule