module fake_aes_463_n_57 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_57);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_57;
wire n_53;
wire n_45;
wire n_38;
wire n_20;
wire n_44;
wire n_54;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_48;
wire n_31;
wire n_22;
wire n_46;
wire n_30;
wire n_16;
wire n_26;
wire n_25;
wire n_33;
wire n_50;
wire n_52;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_55;
wire n_17;
wire n_15;
wire n_56;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_51;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
AND2x2_ASAP7_75t_L g15 ( .A(n_14), .B(n_2), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
OA21x2_ASAP7_75t_L g19 ( .A1(n_9), .A2(n_0), .B(n_12), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_1), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_0), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_6), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_10), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_16), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_16), .B(n_5), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_17), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_17), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_18), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_26), .B(n_21), .Y(n_30) );
OAI21x1_ASAP7_75t_L g31 ( .A1(n_26), .A2(n_18), .B(n_24), .Y(n_31) );
HB1xp67_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_28), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_30), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
BUFx3_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
INVx2_ASAP7_75t_L g38 ( .A(n_34), .Y(n_38) );
INVx2_ASAP7_75t_L g39 ( .A(n_34), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_37), .Y(n_40) );
OR2x2_ASAP7_75t_L g41 ( .A(n_37), .B(n_36), .Y(n_41) );
AOI32xp33_ASAP7_75t_L g42 ( .A1(n_38), .A2(n_35), .A3(n_20), .B1(n_25), .B2(n_21), .Y(n_42) );
AOI21xp33_ASAP7_75t_L g43 ( .A1(n_39), .A2(n_31), .B(n_29), .Y(n_43) );
NAND5xp2_ASAP7_75t_L g44 ( .A(n_42), .B(n_40), .C(n_43), .D(n_28), .E(n_27), .Y(n_44) );
INVxp67_ASAP7_75t_L g45 ( .A(n_41), .Y(n_45) );
AND2x2_ASAP7_75t_L g46 ( .A(n_41), .B(n_19), .Y(n_46) );
O2A1O1Ixp33_ASAP7_75t_L g47 ( .A1(n_41), .A2(n_29), .B(n_23), .C(n_15), .Y(n_47) );
INVx2_ASAP7_75t_L g48 ( .A(n_40), .Y(n_48) );
NOR3xp33_ASAP7_75t_L g49 ( .A(n_47), .B(n_22), .C(n_19), .Y(n_49) );
NOR3xp33_ASAP7_75t_L g50 ( .A(n_44), .B(n_45), .C(n_48), .Y(n_50) );
NOR2x1_ASAP7_75t_L g51 ( .A(n_48), .B(n_22), .Y(n_51) );
XNOR2x1_ASAP7_75t_L g52 ( .A(n_46), .B(n_5), .Y(n_52) );
INVx1_ASAP7_75t_L g53 ( .A(n_50), .Y(n_53) );
AO22x2_ASAP7_75t_L g54 ( .A1(n_52), .A2(n_46), .B1(n_7), .B2(n_8), .Y(n_54) );
AOI22x1_ASAP7_75t_L g55 ( .A1(n_49), .A2(n_22), .B1(n_7), .B2(n_8), .Y(n_55) );
AOI221xp5_ASAP7_75t_L g56 ( .A1(n_54), .A2(n_6), .B1(n_9), .B2(n_51), .C(n_13), .Y(n_56) );
AOI22xp33_ASAP7_75t_L g57 ( .A1(n_56), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_57) );
endmodule