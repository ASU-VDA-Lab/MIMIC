module real_jpeg_24934_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_2),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_15),
.B1(n_19),
.B2(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_2),
.A2(n_24),
.B1(n_32),
.B2(n_35),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_6),
.A2(n_21),
.B1(n_23),
.B2(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_15),
.B1(n_19),
.B2(n_29),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_15),
.C(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_6),
.B(n_32),
.C(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_6),
.B(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_6),
.B(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_6),
.B(n_79),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_44),
.B1(n_73),
.B2(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_84),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_82),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_56),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_12),
.B(n_56),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_30),
.C(n_42),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_13),
.A2(n_30),
.B1(n_91),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_20),
.B(n_25),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

OA22x2_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

INVx5_ASAP7_75t_SL g19 ( 
.A(n_15),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_15),
.A2(n_19),
.B1(n_33),
.B2(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_15),
.B(n_90),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_27)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_21),
.Y(n_23)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_21),
.A2(n_23),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_26),
.A2(n_28),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_30),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_30),
.B(n_92),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_36),
.B(n_38),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_32),
.B(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_42),
.B(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_55),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_63),
.B1(n_64),
.B2(n_81),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_60),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_99),
.C(n_108),
.Y(n_113)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_77),
.B2(n_80),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_76),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_76),
.B(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_112),
.B(n_117),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_103),
.B(n_111),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_93),
.B(n_102),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B(n_101),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_106),
.B1(n_107),
.B2(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);


endmodule