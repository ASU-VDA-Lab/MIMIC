module fake_ariane_1226_n_881 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_881);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_881;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_677;
wire n_614;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_612;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g185 ( 
.A(n_25),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g186 ( 
.A(n_71),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

BUFx8_ASAP7_75t_SL g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_51),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_72),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_143),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_27),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_10),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_78),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_10),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_46),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_158),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_142),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_36),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_99),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_136),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_23),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_92),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_57),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_81),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_120),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_86),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_122),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_6),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_119),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_130),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_2),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_1),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_125),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_144),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_33),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_109),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_14),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_15),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_124),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_79),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_121),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_162),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_47),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_53),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_154),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_20),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_182),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_87),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_129),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_123),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_151),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_103),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_69),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_62),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_176),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_108),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_64),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_1),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_45),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_0),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_0),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_2),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_3),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_188),
.B(n_3),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_197),
.B(n_4),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g278 ( 
.A(n_196),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_196),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_195),
.Y(n_281)
);

BUFx8_ASAP7_75t_SL g282 ( 
.A(n_222),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_202),
.B(n_4),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_5),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_219),
.B(n_5),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_223),
.B(n_6),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_191),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_235),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_202),
.B(n_7),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_189),
.B(n_248),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_7),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_241),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_204),
.B(n_8),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_8),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_212),
.B(n_9),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_187),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_212),
.B(n_9),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_195),
.B(n_200),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_227),
.B(n_11),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_233),
.B(n_193),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_252),
.B(n_254),
.Y(n_307)
);

NAND2x1p5_ASAP7_75t_L g308 ( 
.A(n_217),
.B(n_28),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_239),
.B(n_11),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_225),
.B(n_12),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

OA22x2_ASAP7_75t_L g312 ( 
.A1(n_281),
.A2(n_222),
.B1(n_228),
.B2(n_234),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_306),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_248),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_281),
.A2(n_228),
.B1(n_234),
.B2(n_257),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_261),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_257),
.B1(n_186),
.B2(n_247),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_261),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_269),
.A2(n_186),
.B1(n_246),
.B2(n_245),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_272),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_268),
.A2(n_259),
.B1(n_243),
.B2(n_242),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_265),
.A2(n_240),
.B1(n_236),
.B2(n_232),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_308),
.A2(n_231),
.B1(n_230),
.B2(n_229),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_192),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_289),
.A2(n_270),
.B1(n_266),
.B2(n_274),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_226),
.B1(n_224),
.B2(n_221),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_306),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_268),
.A2(n_215),
.B1(n_214),
.B2(n_211),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_209),
.B1(n_208),
.B2(n_205),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_194),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

AO22x2_ASAP7_75t_L g344 ( 
.A1(n_299),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_291),
.B(n_198),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_277),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_309),
.A2(n_203),
.B1(n_199),
.B2(n_17),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_304),
.B(n_13),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_16),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_308),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_277),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_309),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_283),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_277),
.Y(n_357)
);

AO22x2_ASAP7_75t_L g358 ( 
.A1(n_283),
.A2(n_296),
.B1(n_263),
.B2(n_302),
.Y(n_358)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

AO22x2_ASAP7_75t_L g360 ( 
.A1(n_283),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_283),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_266),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_31),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_293),
.Y(n_364)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_296),
.B(n_32),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_293),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_304),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_314),
.B(n_304),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

XOR2x2_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_282),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_365),
.B(n_296),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

AND2x6_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_304),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_315),
.Y(n_378)
);

NAND2x1_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_291),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_334),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_300),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_304),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_300),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_270),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_317),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_274),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

AND2x2_ASAP7_75t_SL g394 ( 
.A(n_355),
.B(n_263),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_267),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_305),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_330),
.B(n_302),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_326),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_326),
.B(n_278),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_352),
.B(n_260),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_339),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_321),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

NAND2x1p5_ASAP7_75t_L g409 ( 
.A(n_349),
.B(n_263),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_332),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_339),
.B(n_260),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_364),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_358),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_319),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_312),
.B(n_305),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_361),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_361),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_360),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_321),
.B(n_278),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_344),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_363),
.B(n_293),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_351),
.Y(n_428)
);

XNOR2x1_ASAP7_75t_L g429 ( 
.A(n_348),
.B(n_263),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_348),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_359),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_341),
.B(n_267),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_362),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_336),
.B(n_280),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_327),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_371),
.B(n_307),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_413),
.B(n_381),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_279),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_371),
.B(n_290),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_394),
.B(n_279),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_372),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_379),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_390),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_290),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_295),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_394),
.B(n_295),
.Y(n_455)
);

AND2x2_ASAP7_75t_SL g456 ( 
.A(n_423),
.B(n_271),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_383),
.B(n_301),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_301),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_368),
.B(n_293),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_293),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_403),
.B(n_297),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_400),
.B(n_273),
.Y(n_465)
);

AND2x2_ASAP7_75t_SL g466 ( 
.A(n_419),
.B(n_284),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_396),
.B(n_273),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_396),
.B(n_286),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_376),
.Y(n_471)
);

BUFx8_ASAP7_75t_L g472 ( 
.A(n_373),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_392),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_399),
.A2(n_287),
.B(n_285),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_387),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_381),
.B(n_297),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_399),
.A2(n_298),
.B(n_367),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_384),
.B(n_428),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_432),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_421),
.B(n_286),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_406),
.Y(n_487)
);

AND2x2_ASAP7_75t_SL g488 ( 
.A(n_425),
.B(n_275),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_288),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_424),
.B(n_435),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_373),
.B(n_288),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_431),
.B(n_262),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_384),
.B(n_297),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_359),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_395),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_373),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_397),
.B(n_262),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_397),
.B(n_280),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_437),
.B(n_260),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_401),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_409),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_373),
.B(n_264),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_377),
.B(n_264),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_430),
.B(n_297),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_408),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_462),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_459),
.B(n_438),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_443),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_459),
.B(n_438),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_405),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_491),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_476),
.B(n_434),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_491),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_439),
.B(n_409),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_482),
.B(n_405),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_487),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_439),
.B(n_427),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g526 ( 
.A(n_472),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_462),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_477),
.B(n_418),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_427),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_476),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_476),
.B(n_410),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_491),
.B(n_411),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_412),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_450),
.B(n_414),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_444),
.B(n_404),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_462),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_464),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_506),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_446),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_465),
.B(n_382),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_444),
.B(n_415),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_446),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_483),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_455),
.B(n_433),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_448),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_465),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_477),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_498),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_502),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_455),
.B(n_466),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_500),
.B(n_264),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_482),
.B(n_398),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_495),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_464),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_466),
.B(n_297),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_466),
.B(n_297),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_442),
.B(n_294),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_490),
.B(n_370),
.Y(n_560)
);

BUFx8_ASAP7_75t_L g561 ( 
.A(n_502),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_451),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_501),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

NAND2x1_ASAP7_75t_SL g565 ( 
.A(n_503),
.B(n_362),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_474),
.A2(n_310),
.B(n_420),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_450),
.B(n_420),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_523),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_512),
.Y(n_569)
);

CKINVDCx14_ASAP7_75t_R g570 ( 
.A(n_555),
.Y(n_570)
);

BUFx6f_ASAP7_75t_SL g571 ( 
.A(n_543),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_549),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_561),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_561),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_522),
.B(n_490),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_530),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_540),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_550),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_551),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_510),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_564),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_516),
.A2(n_481),
.B1(n_452),
.B2(n_480),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_539),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_563),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_522),
.B(n_503),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_548),
.B(n_492),
.Y(n_592)
);

BUFx12f_ASAP7_75t_L g593 ( 
.A(n_560),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_515),
.B(n_500),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_554),
.B(n_514),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_518),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_528),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_550),
.Y(n_598)
);

INVx6_ASAP7_75t_L g599 ( 
.A(n_518),
.Y(n_599)
);

CKINVDCx11_ASAP7_75t_R g600 ( 
.A(n_518),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_519),
.B(n_472),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_SL g602 ( 
.A1(n_548),
.A2(n_473),
.B1(n_480),
.B2(n_452),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_563),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_524),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_527),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_521),
.Y(n_606)
);

BUFx4f_ASAP7_75t_SL g607 ( 
.A(n_524),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_521),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_SL g609 ( 
.A1(n_514),
.A2(n_472),
.B1(n_488),
.B2(n_473),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_532),
.Y(n_610)
);

INVx8_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_546),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_544),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_544),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_511),
.B(n_501),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_536),
.Y(n_617)
);

BUFx2_ASAP7_75t_SL g618 ( 
.A(n_544),
.Y(n_618)
);

CKINVDCx11_ASAP7_75t_R g619 ( 
.A(n_574),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_611),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_572),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_611),
.Y(n_622)
);

BUFx8_ASAP7_75t_SL g623 ( 
.A(n_574),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_610),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_569),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_595),
.B(n_511),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_595),
.A2(n_472),
.B1(n_546),
.B2(n_538),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_583),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_584),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_586),
.A2(n_516),
.B1(n_552),
.B2(n_520),
.Y(n_630)
);

CKINVDCx14_ASAP7_75t_R g631 ( 
.A(n_570),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_592),
.A2(n_552),
.B1(n_520),
.B2(n_565),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_582),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_587),
.Y(n_634)
);

INVx8_ASAP7_75t_L g635 ( 
.A(n_611),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_571),
.Y(n_636)
);

NAND2x1p5_ASAP7_75t_L g637 ( 
.A(n_596),
.B(n_547),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_588),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_583),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_591),
.A2(n_488),
.B1(n_513),
.B2(n_529),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_616),
.A2(n_603),
.B1(n_576),
.B2(n_559),
.Y(n_641)
);

BUFx4_ASAP7_75t_R g642 ( 
.A(n_580),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_568),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_593),
.A2(n_488),
.B1(n_513),
.B2(n_529),
.Y(n_644)
);

INVx6_ASAP7_75t_L g645 ( 
.A(n_585),
.Y(n_645)
);

AOI22x1_ASAP7_75t_SL g646 ( 
.A1(n_568),
.A2(n_505),
.B1(n_471),
.B2(n_475),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_589),
.Y(n_647)
);

BUFx2_ASAP7_75t_SL g648 ( 
.A(n_571),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_590),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_597),
.A2(n_493),
.B1(n_486),
.B2(n_532),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_600),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_613),
.B(n_457),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_579),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_597),
.A2(n_493),
.B1(n_486),
.B2(n_535),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_609),
.A2(n_594),
.B1(n_468),
.B2(n_593),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_575),
.A2(n_442),
.B1(n_559),
.B2(n_535),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_L g658 ( 
.A1(n_602),
.A2(n_474),
.B(n_525),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_605),
.Y(n_659)
);

CKINVDCx11_ASAP7_75t_R g660 ( 
.A(n_580),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_611),
.Y(n_661)
);

INVx6_ASAP7_75t_L g662 ( 
.A(n_585),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_601),
.A2(n_541),
.B1(n_537),
.B2(n_556),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_SL g664 ( 
.A1(n_646),
.A2(n_570),
.B1(n_529),
.B2(n_601),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_625),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_629),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_655),
.A2(n_601),
.B1(n_504),
.B2(n_479),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_642),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_640),
.A2(n_479),
.B1(n_475),
.B2(n_504),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_634),
.Y(n_670)
);

OAI22x1_ASAP7_75t_SL g671 ( 
.A1(n_619),
.A2(n_499),
.B1(n_484),
.B2(n_571),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_644),
.A2(n_499),
.B1(n_484),
.B2(n_594),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_659),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_626),
.B(n_457),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_641),
.A2(n_529),
.B1(n_594),
.B2(n_456),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_657),
.A2(n_525),
.B1(n_607),
.B2(n_606),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_650),
.A2(n_541),
.B1(n_529),
.B2(n_617),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_645),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_627),
.A2(n_607),
.B1(n_606),
.B2(n_608),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_623),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_628),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_653),
.B(n_467),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_639),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_632),
.A2(n_606),
.B1(n_608),
.B2(n_577),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_635),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_656),
.A2(n_608),
.B1(n_578),
.B2(n_577),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_630),
.A2(n_467),
.B1(n_470),
.B2(n_456),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_645),
.Y(n_688)
);

BUFx12f_ASAP7_75t_L g689 ( 
.A(n_660),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_SL g690 ( 
.A1(n_648),
.A2(n_456),
.B1(n_533),
.B2(n_558),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_633),
.A2(n_578),
.B1(n_577),
.B2(n_557),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_638),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_647),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_643),
.B(n_599),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_633),
.B(n_631),
.Y(n_695)
);

AO22x1_ASAP7_75t_L g696 ( 
.A1(n_651),
.A2(n_652),
.B1(n_624),
.B2(n_654),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_621),
.B(n_651),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_658),
.A2(n_485),
.B1(n_464),
.B2(n_497),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_621),
.B(n_470),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_649),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_658),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_663),
.A2(n_497),
.B1(n_485),
.B2(n_509),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_651),
.A2(n_497),
.B1(n_485),
.B2(n_509),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_637),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_637),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_652),
.B(n_596),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_662),
.B(n_604),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_652),
.A2(n_509),
.B1(n_454),
.B2(n_489),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_662),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_636),
.A2(n_454),
.B1(n_489),
.B2(n_531),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_SL g711 ( 
.A1(n_620),
.A2(n_489),
.B1(n_599),
.B2(n_661),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_636),
.A2(n_454),
.B1(n_489),
.B2(n_531),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_635),
.A2(n_454),
.B1(n_441),
.B2(n_533),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_635),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_661),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_620),
.B(n_604),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_622),
.A2(n_441),
.B1(n_460),
.B2(n_447),
.Y(n_717)
);

OA21x2_ASAP7_75t_L g718 ( 
.A1(n_701),
.A2(n_461),
.B(n_460),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_675),
.A2(n_453),
.B1(n_447),
.B2(n_553),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_669),
.A2(n_622),
.B1(n_578),
.B2(n_562),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_693),
.B(n_612),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_700),
.B(n_612),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_677),
.A2(n_447),
.B1(n_453),
.B2(n_553),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_669),
.A2(n_687),
.B1(n_667),
.B2(n_672),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_676),
.B(n_615),
.C(n_614),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_SL g726 ( 
.A1(n_668),
.A2(n_566),
.B1(n_618),
.B2(n_557),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_665),
.B(n_566),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_SL g728 ( 
.A1(n_668),
.A2(n_558),
.B1(n_599),
.B2(n_547),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_666),
.B(n_614),
.Y(n_729)
);

AOI221xp5_ASAP7_75t_L g730 ( 
.A1(n_674),
.A2(n_483),
.B1(n_461),
.B2(n_507),
.C(n_508),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_667),
.A2(n_450),
.B1(n_507),
.B2(n_562),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_677),
.A2(n_453),
.B1(n_547),
.B2(n_448),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_672),
.A2(n_494),
.B1(n_478),
.B2(n_598),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_670),
.B(n_614),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_664),
.A2(n_448),
.B1(n_508),
.B2(n_615),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_682),
.A2(n_690),
.B1(n_702),
.B2(n_673),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_702),
.A2(n_615),
.B1(n_614),
.B2(n_534),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_681),
.A2(n_615),
.B1(n_534),
.B2(n_494),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_683),
.A2(n_478),
.B1(n_463),
.B2(n_581),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_SL g740 ( 
.A1(n_684),
.A2(n_573),
.B1(n_581),
.B2(n_598),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_699),
.A2(n_463),
.B1(n_451),
.B2(n_469),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_708),
.A2(n_710),
.B1(n_712),
.B2(n_703),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_708),
.A2(n_469),
.B1(n_451),
.B2(n_573),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_710),
.A2(n_469),
.B1(n_573),
.B2(n_598),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_712),
.A2(n_573),
.B1(n_498),
.B2(n_458),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_692),
.B(n_449),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_SL g747 ( 
.A1(n_679),
.A2(n_567),
.B1(n_458),
.B2(n_449),
.Y(n_747)
);

OAI211xp5_ASAP7_75t_SL g748 ( 
.A1(n_694),
.A2(n_458),
.B(n_449),
.C(n_40),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_671),
.A2(n_458),
.B1(n_449),
.B2(n_567),
.Y(n_749)
);

OAI222xp33_ASAP7_75t_L g750 ( 
.A1(n_703),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.C1(n_43),
.C2(n_48),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_691),
.A2(n_498),
.B1(n_496),
.B2(n_420),
.Y(n_751)
);

OAI222xp33_ASAP7_75t_L g752 ( 
.A1(n_706),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.C1(n_54),
.C2(n_55),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_697),
.A2(n_713),
.B1(n_695),
.B2(n_698),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_698),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_L g755 ( 
.A1(n_678),
.A2(n_498),
.B1(n_496),
.B2(n_59),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_713),
.A2(n_498),
.B1(n_58),
.B2(n_60),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_696),
.B(n_498),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_734),
.B(n_727),
.Y(n_758)
);

OAI221xp5_ASAP7_75t_SL g759 ( 
.A1(n_736),
.A2(n_688),
.B1(n_717),
.B2(n_709),
.C(n_707),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_724),
.A2(n_686),
.B1(n_689),
.B2(n_711),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_SL g761 ( 
.A1(n_725),
.A2(n_752),
.B(n_753),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_734),
.B(n_716),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_727),
.B(n_722),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_729),
.B(n_717),
.C(n_705),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_721),
.B(n_715),
.Y(n_765)
);

NAND4xp25_ASAP7_75t_L g766 ( 
.A(n_746),
.B(n_730),
.C(n_748),
.D(n_731),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_757),
.B(n_704),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_726),
.B(n_714),
.C(n_685),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_757),
.B(n_685),
.Y(n_769)
);

AOI221xp5_ASAP7_75t_L g770 ( 
.A1(n_733),
.A2(n_754),
.B1(n_755),
.B2(n_750),
.C(n_741),
.Y(n_770)
);

AOI221xp5_ASAP7_75t_L g771 ( 
.A1(n_742),
.A2(n_680),
.B1(n_61),
.B2(n_63),
.C(n_65),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_718),
.Y(n_772)
);

AND2x2_ASAP7_75t_SL g773 ( 
.A(n_718),
.B(n_56),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_718),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_731),
.B(n_66),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_740),
.B(n_184),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_747),
.B(n_67),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_728),
.B(n_183),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_749),
.B(n_68),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_720),
.B(n_180),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_735),
.B(n_73),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_SL g782 ( 
.A(n_744),
.B(n_74),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_738),
.B(n_75),
.C(n_77),
.Y(n_783)
);

AOI221xp5_ASAP7_75t_L g784 ( 
.A1(n_756),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.C(n_85),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_737),
.B(n_745),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_751),
.B(n_88),
.C(n_89),
.Y(n_786)
);

NAND4xp25_ASAP7_75t_L g787 ( 
.A(n_732),
.B(n_90),
.C(n_91),
.D(n_93),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_SL g788 ( 
.A1(n_719),
.A2(n_94),
.B(n_95),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_739),
.B(n_177),
.Y(n_789)
);

NOR3xp33_ASAP7_75t_L g790 ( 
.A(n_760),
.B(n_723),
.C(n_743),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_758),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_763),
.B(n_97),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_769),
.B(n_98),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_765),
.B(n_100),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_762),
.B(n_101),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_766),
.B(n_760),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_767),
.B(n_102),
.Y(n_797)
);

OAI221xp5_ASAP7_75t_SL g798 ( 
.A1(n_761),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.C(n_107),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_764),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_772),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_768),
.B(n_110),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_774),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_785),
.B(n_111),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_SL g804 ( 
.A(n_771),
.B(n_112),
.C(n_113),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_773),
.B(n_114),
.Y(n_805)
);

NOR2x1_ASAP7_75t_L g806 ( 
.A(n_780),
.B(n_115),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_770),
.B(n_116),
.C(n_117),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_800),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_800),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_802),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_802),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_791),
.Y(n_812)
);

NAND4xp75_ASAP7_75t_SL g813 ( 
.A(n_796),
.B(n_778),
.C(n_781),
.D(n_773),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_SL g814 ( 
.A(n_803),
.B(n_801),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_799),
.B(n_775),
.Y(n_815)
);

OAI22x1_ASAP7_75t_L g816 ( 
.A1(n_796),
.A2(n_779),
.B1(n_783),
.B2(n_786),
.Y(n_816)
);

NOR4xp25_ASAP7_75t_L g817 ( 
.A(n_798),
.B(n_759),
.C(n_787),
.D(n_788),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_815),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_815),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_812),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_808),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_810),
.Y(n_822)
);

XNOR2xp5_ASAP7_75t_L g823 ( 
.A(n_818),
.B(n_813),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_819),
.Y(n_824)
);

XNOR2x1_ASAP7_75t_L g825 ( 
.A(n_820),
.B(n_816),
.Y(n_825)
);

AO22x2_ASAP7_75t_L g826 ( 
.A1(n_822),
.A2(n_801),
.B1(n_809),
.B2(n_811),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_824),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_825),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_826),
.Y(n_829)
);

AOI322xp5_ASAP7_75t_L g830 ( 
.A1(n_823),
.A2(n_814),
.A3(n_801),
.B1(n_790),
.B2(n_822),
.C1(n_805),
.C2(n_806),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_827),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_828),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_831),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_831),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_832),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_835),
.B(n_828),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_833),
.B(n_834),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_834),
.A2(n_829),
.B1(n_826),
.B2(n_817),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_835),
.A2(n_816),
.B1(n_807),
.B2(n_830),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_835),
.A2(n_804),
.B1(n_793),
.B2(n_821),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_835),
.B(n_793),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_836),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_837),
.B(n_795),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_838),
.A2(n_795),
.B1(n_794),
.B2(n_792),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_839),
.A2(n_782),
.B1(n_797),
.B2(n_809),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_840),
.A2(n_811),
.B1(n_789),
.B2(n_776),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_841),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_837),
.B(n_784),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_842),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_843),
.Y(n_850)
);

AND4x1_ASAP7_75t_L g851 ( 
.A(n_845),
.B(n_777),
.C(n_759),
.D(n_127),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_847),
.B(n_118),
.Y(n_852)
);

OA22x2_ASAP7_75t_L g853 ( 
.A1(n_848),
.A2(n_844),
.B1(n_846),
.B2(n_131),
.Y(n_853)
);

NOR2x1_ASAP7_75t_L g854 ( 
.A(n_842),
.B(n_126),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_849),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_854),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_850),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_852),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_853),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_851),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_849),
.Y(n_861)
);

OA22x2_ASAP7_75t_L g862 ( 
.A1(n_855),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_862)
);

AOI22x1_ASAP7_75t_L g863 ( 
.A1(n_861),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_863)
);

AO22x2_ASAP7_75t_L g864 ( 
.A1(n_856),
.A2(n_139),
.B1(n_141),
.B2(n_145),
.Y(n_864)
);

AO22x2_ASAP7_75t_L g865 ( 
.A1(n_857),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_858),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_860),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_858),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_866),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_863),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_868),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_862),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_869),
.A2(n_859),
.B1(n_865),
.B2(n_864),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_872),
.A2(n_867),
.B1(n_156),
.B2(n_157),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_871),
.A2(n_155),
.B1(n_160),
.B2(n_164),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_873),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_875),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_876),
.A2(n_870),
.B1(n_874),
.B2(n_167),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_878),
.Y(n_879)
);

AOI221xp5_ASAP7_75t_L g880 ( 
.A1(n_879),
.A2(n_877),
.B1(n_166),
.B2(n_168),
.C(n_169),
.Y(n_880)
);

AOI211xp5_ASAP7_75t_L g881 ( 
.A1(n_880),
.A2(n_165),
.B(n_170),
.C(n_172),
.Y(n_881)
);


endmodule