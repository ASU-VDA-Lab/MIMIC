module fake_jpeg_1710_n_73 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_23),
.B(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_27),
.B1(n_22),
.B2(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_10),
.Y(n_44)
);

NAND2x1_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_27),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_31),
.C(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_46),
.Y(n_49)
);

OA21x2_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_39),
.B(n_34),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_36),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_12),
.C(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_59),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_35),
.B1(n_5),
.B2(n_6),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_58),
.B(n_49),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_35),
.B1(n_5),
.B2(n_7),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_11),
.C(n_17),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_62),
.B(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_4),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_7),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_60),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_60),
.C(n_13),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_16),
.B(n_18),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_68),
.C(n_9),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_66),
.C(n_64),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_8),
.Y(n_73)
);


endmodule