module real_aes_7491_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_1067;
wire n_518;
wire n_673;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_551;
wire n_666;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_1021;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_1040;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_743;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_994;
wire n_495;
wire n_1072;
wire n_892;
wire n_1078;
wire n_938;
wire n_744;
wire n_384;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_746;
wire n_532;
wire n_656;
wire n_1025;
wire n_1148;
wire n_409;
wire n_860;
wire n_748;
wire n_909;
wire n_523;
wire n_781;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_1006;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1037;
wire n_1031;
wire n_1131;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_1079;
wire n_843;
wire n_810;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_972;
wire n_1127;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_1068;
wire n_492;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_1150;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_710;
wire n_823;
wire n_393;
wire n_652;
wire n_1097;
wire n_703;
wire n_601;
wire n_1101;
wire n_500;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_0), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_1), .A2(n_298), .B1(n_456), .B2(n_625), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_2), .A2(n_158), .B1(n_518), .B2(n_521), .Y(n_1056) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_3), .Y(n_450) );
INVx1_ASAP7_75t_L g1051 ( .A(n_4), .Y(n_1051) );
AOI22xp33_ASAP7_75t_SL g754 ( .A1(n_5), .A2(n_347), .B1(n_714), .B2(n_755), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g942 ( .A1(n_6), .A2(n_132), .B1(n_521), .B2(n_808), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_7), .Y(n_697) );
AOI222xp33_ASAP7_75t_L g730 ( .A1(n_8), .A2(n_186), .B1(n_303), .B2(n_534), .C1(n_568), .C2(n_577), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_9), .A2(n_100), .B1(n_520), .B2(n_923), .Y(n_1038) );
AO22x2_ASAP7_75t_L g415 ( .A1(n_10), .A2(n_219), .B1(n_407), .B2(n_412), .Y(n_415) );
INVx1_ASAP7_75t_L g1080 ( .A(n_10), .Y(n_1080) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_11), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_12), .A2(n_147), .B1(n_507), .B2(n_601), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g946 ( .A1(n_13), .A2(n_326), .B1(n_334), .B2(n_580), .C1(n_581), .C2(n_774), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g1066 ( .A(n_14), .Y(n_1066) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_15), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_16), .A2(n_212), .B1(n_520), .B2(n_782), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_17), .A2(n_49), .B1(n_795), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_18), .A2(n_118), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_19), .A2(n_290), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g1020 ( .A1(n_20), .A2(n_245), .B1(n_594), .B2(n_1021), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_21), .A2(n_228), .B1(n_506), .B2(n_1146), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_22), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_23), .A2(n_263), .B1(n_506), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_24), .A2(n_362), .B1(n_621), .B2(n_955), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_25), .A2(n_91), .B1(n_580), .B2(n_581), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_26), .A2(n_201), .B1(n_594), .B2(n_1021), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_27), .A2(n_318), .B1(n_530), .B2(n_719), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g1052 ( .A1(n_28), .A2(n_190), .B1(n_533), .B2(n_535), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_29), .A2(n_110), .B1(n_591), .B2(n_713), .C(n_715), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_30), .A2(n_154), .B1(n_447), .B2(n_898), .Y(n_945) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_31), .A2(n_136), .B1(n_504), .B2(n_896), .Y(n_1040) );
AOI22xp33_ASAP7_75t_SL g614 ( .A1(n_32), .A2(n_83), .B1(n_516), .B2(n_553), .Y(n_614) );
AO22x2_ASAP7_75t_L g417 ( .A1(n_33), .A2(n_117), .B1(n_407), .B2(n_408), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g750 ( .A1(n_34), .A2(n_270), .B1(n_507), .B2(n_672), .Y(n_750) );
INVx1_ASAP7_75t_L g1126 ( .A(n_35), .Y(n_1126) );
AOI222xp33_ASAP7_75t_L g812 ( .A1(n_36), .A2(n_188), .B1(n_302), .B2(n_535), .C1(n_553), .C2(n_609), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_37), .B(n_1037), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_38), .A2(n_74), .B1(n_672), .B2(n_720), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_39), .A2(n_262), .B1(n_705), .B2(n_898), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_40), .A2(n_197), .B1(n_551), .B2(n_616), .C(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_41), .B(n_569), .Y(n_1009) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_42), .A2(n_119), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_43), .A2(n_366), .B1(n_420), .B2(n_447), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_44), .A2(n_126), .B1(n_553), .B2(n_782), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_45), .A2(n_77), .B1(n_669), .B2(n_787), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_46), .A2(n_321), .B1(n_563), .B2(n_590), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_47), .A2(n_96), .B1(n_672), .B2(n_757), .Y(n_987) );
AOI222xp33_ASAP7_75t_L g480 ( .A1(n_48), .A2(n_79), .B1(n_135), .B2(n_481), .C1(n_485), .C2(n_489), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_50), .A2(n_142), .B1(n_501), .B2(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g559 ( .A(n_51), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_52), .B(n_485), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_53), .A2(n_120), .B1(n_624), .B2(n_625), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_54), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_55), .A2(n_284), .B1(n_540), .B2(n_837), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_56), .A2(n_226), .B1(n_566), .B2(n_672), .Y(n_1063) );
AOI222xp33_ASAP7_75t_L g844 ( .A1(n_57), .A2(n_171), .B1(n_343), .B2(n_484), .C1(n_612), .C2(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_58), .A2(n_92), .B1(n_702), .B2(n_938), .Y(n_937) );
CKINVDCx20_ASAP7_75t_R g1003 ( .A(n_59), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_60), .Y(n_866) );
INVx1_ASAP7_75t_L g724 ( .A(n_61), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_62), .A2(n_181), .B1(n_516), .B2(n_520), .Y(n_515) );
INVx1_ASAP7_75t_L g759 ( .A(n_63), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_64), .B(n_462), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_65), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g1043 ( .A1(n_66), .A2(n_380), .B1(n_713), .B2(n_1044), .Y(n_1043) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_67), .A2(n_159), .B1(n_895), .B2(n_896), .Y(n_894) );
AOI22xp33_ASAP7_75t_SL g756 ( .A1(n_68), .A2(n_222), .B1(n_757), .B2(n_758), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_69), .A2(n_301), .B1(n_757), .B2(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g1130 ( .A(n_70), .Y(n_1130) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_71), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_72), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_73), .A2(n_337), .B1(n_834), .B2(n_837), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_75), .A2(n_375), .B1(n_516), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_76), .A2(n_353), .B1(n_566), .B2(n_1141), .Y(n_1140) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_78), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_80), .A2(n_259), .B1(n_591), .B2(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_81), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_82), .A2(n_202), .B1(n_792), .B2(n_793), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_84), .A2(n_194), .B1(n_594), .B2(n_1021), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_85), .A2(n_255), .B1(n_447), .B2(n_672), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_86), .A2(n_108), .B1(n_719), .B2(n_720), .C(n_722), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_87), .Y(n_826) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_88), .A2(n_261), .B1(n_407), .B2(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g1077 ( .A(n_88), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_89), .A2(n_145), .B1(n_485), .B2(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_90), .A2(n_233), .B1(n_591), .B2(n_1019), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_93), .A2(n_285), .B1(n_442), .B2(n_566), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_94), .A2(n_127), .B1(n_465), .B2(n_551), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g1002 ( .A(n_95), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g747 ( .A1(n_97), .A2(n_272), .B1(n_518), .B2(n_533), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_98), .A2(n_183), .B1(n_461), .B2(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_99), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_101), .A2(n_820), .B1(n_846), .B2(n_847), .Y(n_819) );
CKINVDCx16_ASAP7_75t_R g846 ( .A(n_101), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g1089 ( .A(n_102), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_103), .A2(n_373), .B1(n_568), .B2(n_808), .Y(n_807) );
AOI222xp33_ASAP7_75t_L g989 ( .A1(n_104), .A2(n_114), .B1(n_173), .B2(n_577), .C1(n_581), .C2(n_587), .Y(n_989) );
AOI22xp5_ASAP7_75t_L g998 ( .A1(n_105), .A2(n_999), .B1(n_1022), .B2(n_1023), .Y(n_998) );
INVx1_ASAP7_75t_L g1022 ( .A(n_105), .Y(n_1022) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_106), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_107), .A2(n_265), .B1(n_758), .B2(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g728 ( .A(n_109), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_111), .Y(n_957) );
XOR2x2_ASAP7_75t_L g908 ( .A(n_112), .B(n_909), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_113), .A2(n_130), .B1(n_1019), .B2(n_1144), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_115), .A2(n_279), .B1(n_421), .B2(n_590), .Y(n_944) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_116), .Y(n_740) );
INVx1_ASAP7_75t_L g1081 ( .A(n_117), .Y(n_1081) );
XOR2x2_ASAP7_75t_L g572 ( .A(n_121), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_122), .B(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_123), .A2(n_275), .B1(n_705), .B2(n_706), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_124), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g969 ( .A(n_125), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_128), .B(n_919), .Y(n_918) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_129), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g1137 ( .A1(n_131), .A2(n_242), .B1(n_674), .B2(n_1138), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_133), .A2(n_348), .B1(n_442), .B2(n_714), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_134), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_137), .A2(n_140), .B1(n_421), .B2(n_590), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g964 ( .A(n_138), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_139), .A2(n_711), .B1(n_731), .B2(n_732), .Y(n_710) );
INVx1_ASAP7_75t_L g731 ( .A(n_139), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_141), .A2(n_283), .B1(n_433), .B2(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g723 ( .A(n_143), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_144), .A2(n_345), .B1(n_506), .B2(n_510), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_146), .A2(n_358), .B1(n_628), .B2(n_837), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_148), .A2(n_193), .B1(n_533), .B2(n_612), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g1087 ( .A(n_149), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_150), .A2(n_200), .B1(n_553), .B2(n_808), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_151), .A2(n_307), .B1(n_526), .B2(n_626), .Y(n_936) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_152), .A2(n_341), .B1(n_456), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_153), .A2(n_252), .B1(n_506), .B2(n_702), .Y(n_701) );
AND2x6_ASAP7_75t_L g385 ( .A(n_155), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1074 ( .A(n_155), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_156), .A2(n_288), .B1(n_510), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g1031 ( .A1(n_157), .A2(n_266), .B1(n_569), .B2(n_1032), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_160), .A2(n_325), .B1(n_542), .B2(n_669), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_161), .A2(n_239), .B1(n_258), .B2(n_484), .C1(n_568), .C2(n_569), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g947 ( .A(n_162), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_163), .A2(n_315), .B1(n_501), .B2(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g570 ( .A(n_164), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_165), .A2(n_339), .B1(n_706), .B2(n_825), .Y(n_1046) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_166), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_167), .A2(n_360), .B1(n_621), .B2(n_752), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_168), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g1008 ( .A(n_169), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_170), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_172), .A2(n_249), .B1(n_530), .B2(n_542), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g972 ( .A(n_174), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_175), .Y(n_861) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_176), .A2(n_250), .B1(n_407), .B2(n_408), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g1078 ( .A(n_176), .B(n_1079), .Y(n_1078) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_177), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_178), .A2(n_210), .B1(n_510), .B2(n_931), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g940 ( .A(n_179), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g666 ( .A(n_180), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_182), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_184), .A2(n_370), .B1(n_528), .B2(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g1030 ( .A(n_185), .Y(n_1030) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_187), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_189), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_191), .A2(n_254), .B1(n_524), .B2(n_526), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_192), .A2(n_342), .B1(n_433), .B2(n_620), .Y(n_619) );
XOR2x2_ASAP7_75t_L g976 ( .A(n_195), .B(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_196), .A2(n_276), .B1(n_551), .B2(n_616), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_198), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_199), .Y(n_842) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_203), .A2(n_204), .B1(n_625), .B2(n_757), .Y(n_785) );
INVx1_ASAP7_75t_L g561 ( .A(n_205), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g1083 ( .A1(n_206), .A2(n_1084), .B1(n_1107), .B2(n_1108), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g1107 ( .A(n_206), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_207), .A2(n_305), .B1(n_744), .B2(n_746), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_208), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_209), .B(n_612), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_211), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_213), .A2(n_267), .B1(n_621), .B2(n_714), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_214), .B(n_513), .Y(n_1035) );
INVx1_ASAP7_75t_L g975 ( .A(n_215), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_216), .A2(n_297), .B1(n_591), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1128 ( .A(n_217), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_218), .A2(n_247), .B1(n_490), .B2(n_520), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_220), .A2(n_287), .B1(n_504), .B2(n_752), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_221), .A2(n_299), .B1(n_516), .B2(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_223), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_224), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_225), .A2(n_289), .B1(n_563), .B2(n_758), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_227), .A2(n_369), .B1(n_434), .B2(n_755), .Y(n_982) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_229), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_230), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_231), .Y(n_876) );
INVx1_ASAP7_75t_L g556 ( .A(n_232), .Y(n_556) );
INVx1_ASAP7_75t_L g729 ( .A(n_234), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_235), .A2(n_333), .B1(n_568), .B2(n_808), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g1092 ( .A(n_236), .Y(n_1092) );
INVx1_ASAP7_75t_L g1117 ( .A(n_237), .Y(n_1117) );
AOI22xp5_ASAP7_75t_SL g1121 ( .A1(n_237), .A2(n_1117), .B1(n_1122), .B2(n_1147), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_238), .A2(n_264), .B1(n_434), .B2(n_621), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_240), .A2(n_381), .B1(n_461), .B2(n_465), .C(n_467), .Y(n_460) );
AOI222xp33_ASAP7_75t_L g532 ( .A1(n_241), .A2(n_349), .B1(n_363), .B2(n_484), .C1(n_533), .C2(n_534), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_243), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_244), .A2(n_379), .B1(n_461), .B2(n_616), .Y(n_891) );
AND2x2_ASAP7_75t_L g389 ( .A(n_246), .B(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_248), .A2(n_281), .B1(n_490), .B2(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g1125 ( .A(n_251), .Y(n_1125) );
XNOR2xp5_ASAP7_75t_L g879 ( .A(n_253), .B(n_880), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_256), .A2(n_683), .B1(n_684), .B2(n_708), .Y(n_682) );
CKINVDCx14_ASAP7_75t_R g708 ( .A(n_256), .Y(n_708) );
INVx1_ASAP7_75t_L g1134 ( .A(n_257), .Y(n_1134) );
CKINVDCx20_ASAP7_75t_R g1091 ( .A(n_260), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_268), .A2(n_294), .B1(n_624), .B2(n_706), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_269), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_271), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_273), .A2(n_377), .B1(n_600), .B2(n_601), .Y(n_599) );
XOR2x2_ASAP7_75t_L g1026 ( .A(n_274), .B(n_1027), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_277), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_278), .A2(n_383), .B(n_391), .C(n_1082), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_280), .Y(n_468) );
OA22x2_ASAP7_75t_L g768 ( .A1(n_282), .A2(n_769), .B1(n_770), .B2(n_796), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_282), .Y(n_769) );
INVx1_ASAP7_75t_L g407 ( .A(n_286), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_286), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_291), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_292), .B(n_462), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_293), .Y(n_958) );
INVx1_ASAP7_75t_L g717 ( .A(n_295), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_296), .B(n_746), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_300), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_304), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_306), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_308), .B(n_489), .Y(n_1131) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_309), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_310), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_311), .A2(n_331), .B1(n_795), .B2(n_1019), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_312), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_313), .B(n_551), .Y(n_1055) );
OA22x2_ASAP7_75t_L g603 ( .A1(n_314), .A2(n_604), .B1(n_605), .B2(n_629), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_314), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_316), .A2(n_376), .B1(n_462), .B2(n_466), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_317), .A2(n_351), .B1(n_457), .B2(n_674), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g667 ( .A(n_319), .Y(n_667) );
INVx1_ASAP7_75t_L g390 ( .A(n_320), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_322), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_323), .B(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g386 ( .A(n_324), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_327), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_328), .A2(n_332), .B1(n_755), .B2(n_758), .Y(n_810) );
INVx1_ASAP7_75t_L g564 ( .A(n_329), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_330), .Y(n_440) );
AO22x2_ASAP7_75t_L g397 ( .A1(n_335), .A2(n_398), .B1(n_493), .B2(n_494), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_335), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_336), .Y(n_775) );
INVx1_ASAP7_75t_L g716 ( .A(n_338), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_340), .A2(n_361), .B1(n_542), .B2(n_900), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_344), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_346), .Y(n_1096) );
CKINVDCx20_ASAP7_75t_R g974 ( .A(n_350), .Y(n_974) );
INVx1_ASAP7_75t_L g545 ( .A(n_352), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_354), .B(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_355), .A2(n_374), .B1(n_524), .B2(n_1060), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_356), .B(n_513), .Y(n_584) );
XOR2x2_ASAP7_75t_L g497 ( .A(n_357), .B(n_498), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_359), .A2(n_639), .B1(n_676), .B2(n_677), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_359), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_364), .B(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_365), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_367), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_368), .Y(n_445) );
INVx1_ASAP7_75t_L g1133 ( .A(n_371), .Y(n_1133) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_372), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_378), .A2(n_852), .B1(n_877), .B2(n_878), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_378), .Y(n_877) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_386), .Y(n_1073) );
OAI21xp5_ASAP7_75t_L g1115 ( .A1(n_387), .A2(n_1072), .B(n_1116), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_815), .B1(n_1067), .B2(n_1068), .C(n_1069), .Y(n_391) );
INVx1_ASAP7_75t_L g1068 ( .A(n_392), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_633), .B1(n_634), .B2(n_814), .Y(n_392) );
INVx1_ASAP7_75t_SL g814 ( .A(n_393), .Y(n_814) );
OAI22xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_571), .B1(n_631), .B2(n_632), .Y(n_393) );
INVx1_ASAP7_75t_L g631 ( .A(n_394), .Y(n_631) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_495), .B2(n_496), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g494 ( .A(n_398), .Y(n_494) );
AND4x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_438), .C(n_460), .D(n_480), .Y(n_398) );
NOR2xp33_ASAP7_75t_SL g399 ( .A(n_400), .B(n_424), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_418), .B2(n_419), .Y(n_400) );
INVx3_ASAP7_75t_L g628 ( .A(n_402), .Y(n_628) );
INVx3_ASAP7_75t_L g1065 ( .A(n_402), .Y(n_1065) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx2_ASAP7_75t_SL g501 ( .A(n_403), .Y(n_501) );
BUFx2_ASAP7_75t_SL g590 ( .A(n_403), .Y(n_590) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_403), .Y(n_714) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_413), .Y(n_403) );
AND2x6_ASAP7_75t_L g442 ( .A(n_404), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g448 ( .A(n_404), .B(n_428), .Y(n_448) );
AND2x6_ASAP7_75t_L g484 ( .A(n_404), .B(n_477), .Y(n_484) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_410), .Y(n_404) );
AND2x2_ASAP7_75t_L g423 ( .A(n_405), .B(n_411), .Y(n_423) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g429 ( .A(n_406), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_406), .B(n_411), .Y(n_437) );
AND2x2_ASAP7_75t_L g471 ( .A(n_406), .B(n_415), .Y(n_471) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_409), .Y(n_412) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g430 ( .A(n_411), .Y(n_430) );
INVx1_ASAP7_75t_L g488 ( .A(n_411), .Y(n_488) );
AND2x4_ASAP7_75t_L g422 ( .A(n_413), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_413), .B(n_429), .Y(n_453) );
AND2x4_ASAP7_75t_L g458 ( .A(n_413), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g525 ( .A(n_413), .B(n_429), .Y(n_525) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .Y(n_413) );
AND2x2_ASAP7_75t_L g428 ( .A(n_414), .B(n_417), .Y(n_428) );
OR2x2_ASAP7_75t_L g444 ( .A(n_414), .B(n_417), .Y(n_444) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g477 ( .A(n_415), .B(n_417), .Y(n_477) );
INVx1_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
AND2x2_ASAP7_75t_L g487 ( .A(n_416), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g436 ( .A(n_417), .Y(n_436) );
OAI221xp5_ASAP7_75t_SL g854 ( .A1(n_419), .A2(n_855), .B1(n_856), .B2(n_857), .C(n_858), .Y(n_854) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g831 ( .A(n_421), .Y(n_831) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_422), .Y(n_504) );
INVx2_ASAP7_75t_L g592 ( .A(n_422), .Y(n_592) );
BUFx3_ASAP7_75t_L g795 ( .A(n_422), .Y(n_795) );
BUFx3_ASAP7_75t_L g931 ( .A(n_422), .Y(n_931) );
AND2x4_ASAP7_75t_L g464 ( .A(n_423), .B(n_443), .Y(n_464) );
AND2x6_ASAP7_75t_L g466 ( .A(n_423), .B(n_428), .Y(n_466) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_423), .B(n_428), .Y(n_548) );
INVx1_ASAP7_75t_L g645 ( .A(n_423), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_431), .B2(n_432), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_426), .A2(n_435), .B1(n_716), .B2(n_717), .Y(n_715) );
BUFx2_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AND2x2_ASAP7_75t_L g509 ( .A(n_428), .B(n_429), .Y(n_509) );
INVx1_ASAP7_75t_L g479 ( .A(n_430), .Y(n_479) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g510 ( .A(n_434), .Y(n_510) );
BUFx2_ASAP7_75t_L g594 ( .A(n_434), .Y(n_594) );
BUFx2_ASAP7_75t_L g702 ( .A(n_434), .Y(n_702) );
BUFx4f_ASAP7_75t_SL g1146 ( .A(n_434), .Y(n_1146) );
INVx6_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g669 ( .A(n_435), .Y(n_669) );
INVx1_ASAP7_75t_SL g900 ( .A(n_435), .Y(n_900) );
INVx1_ASAP7_75t_L g955 ( .A(n_435), .Y(n_955) );
OR2x6_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g519 ( .A(n_436), .Y(n_519) );
INVx1_ASAP7_75t_L g459 ( .A(n_437), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g438 ( .A(n_439), .B(n_449), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_445), .B2(n_446), .Y(n_439) );
INVx3_ASAP7_75t_L g563 ( .A(n_441), .Y(n_563) );
INVx2_ASAP7_75t_SL g600 ( .A(n_441), .Y(n_600) );
INVx4_ASAP7_75t_L g624 ( .A(n_441), .Y(n_624) );
INVx4_ASAP7_75t_L g672 ( .A(n_441), .Y(n_672) );
INVx11_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx11_ASAP7_75t_L g529 ( .A(n_442), .Y(n_529) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g644 ( .A(n_444), .B(n_645), .Y(n_644) );
OAI221xp5_ASAP7_75t_SL g859 ( .A1(n_446), .A2(n_557), .B1(n_860), .B2(n_861), .C(n_862), .Y(n_859) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx6_ASAP7_75t_L g531 ( .A(n_448), .Y(n_531) );
BUFx3_ASAP7_75t_L g601 ( .A(n_448), .Y(n_601) );
BUFx3_ASAP7_75t_L g757 ( .A(n_448), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_454), .B2(n_455), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_451), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g557 ( .A(n_452), .Y(n_557) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
BUFx2_ASAP7_75t_SL g598 ( .A(n_458), .Y(n_598) );
BUFx2_ASAP7_75t_SL g706 ( .A(n_458), .Y(n_706) );
BUFx3_ASAP7_75t_L g758 ( .A(n_458), .Y(n_758) );
BUFx3_ASAP7_75t_L g837 ( .A(n_458), .Y(n_837) );
INVx1_ASAP7_75t_L g985 ( .A(n_458), .Y(n_985) );
BUFx2_ASAP7_75t_L g1060 ( .A(n_458), .Y(n_1060) );
AND2x2_ASAP7_75t_L g752 ( .A(n_459), .B(n_472), .Y(n_752) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_462), .Y(n_919) );
INVx5_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g551 ( .A(n_463), .Y(n_551) );
INVx2_ASAP7_75t_L g744 ( .A(n_463), .Y(n_744) );
INVx2_ASAP7_75t_L g1037 ( .A(n_463), .Y(n_1037) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g514 ( .A(n_466), .Y(n_514) );
BUFx4f_ASAP7_75t_L g746 ( .A(n_466), .Y(n_746) );
BUFx2_ASAP7_75t_L g921 ( .A(n_466), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_473), .B2(n_474), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_469), .A2(n_475), .B1(n_728), .B2(n_729), .Y(n_727) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx4_ASAP7_75t_L g659 ( .A(n_470), .Y(n_659) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_470), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_470), .A2(n_474), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x4_ASAP7_75t_L g486 ( .A(n_471), .B(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g491 ( .A(n_471), .B(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g518 ( .A(n_471), .B(n_519), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_474), .A2(n_965), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g662 ( .A(n_475), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_475), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_475), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g521 ( .A(n_477), .B(n_479), .Y(n_521) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI21xp5_ASAP7_75t_SL g691 ( .A1(n_482), .A2(n_692), .B(n_693), .Y(n_691) );
BUFx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g774 ( .A(n_483), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_483), .A2(n_654), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_967) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_484), .Y(n_577) );
BUFx3_ASAP7_75t_L g609 ( .A(n_484), .Y(n_609) );
INVx2_ASAP7_75t_L g739 ( .A(n_484), .Y(n_739) );
INVx2_ASAP7_75t_SL g870 ( .A(n_484), .Y(n_870) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx4f_ASAP7_75t_SL g533 ( .A(n_486), .Y(n_533) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_486), .Y(n_568) );
BUFx2_ASAP7_75t_L g845 ( .A(n_486), .Y(n_845) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_486), .Y(n_885) );
INVx1_ASAP7_75t_L g492 ( .A(n_488), .Y(n_492) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g612 ( .A(n_490), .Y(n_612) );
INVx2_ASAP7_75t_L g654 ( .A(n_490), .Y(n_654) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx12f_ASAP7_75t_L g535 ( .A(n_491), .Y(n_535) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_491), .Y(n_569) );
INVx1_ASAP7_75t_L g887 ( .A(n_491), .Y(n_887) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
XOR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_536), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_497), .A2(n_638), .B1(n_678), .B2(n_679), .Y(n_637) );
INVx1_ASAP7_75t_L g678 ( .A(n_497), .Y(n_678) );
NAND4xp75_ASAP7_75t_L g498 ( .A(n_499), .B(n_511), .C(n_522), .D(n_532), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .Y(n_499) );
INVx1_ASAP7_75t_L g665 ( .A(n_501), .Y(n_665) );
INVx4_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g540 ( .A(n_503), .Y(n_540) );
OAI221xp5_ASAP7_75t_SL g664 ( .A1(n_503), .A2(n_665), .B1(n_666), .B2(n_667), .C(n_668), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_503), .A2(n_725), .B1(n_960), .B2(n_961), .Y(n_959) );
INVx4_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g1021 ( .A(n_507), .Y(n_1021) );
INVx5_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx3_ASAP7_75t_L g543 ( .A(n_508), .Y(n_543) );
INVx2_ASAP7_75t_L g621 ( .A(n_508), .Y(n_621) );
INVx1_ASAP7_75t_L g788 ( .A(n_508), .Y(n_788) );
INVx3_ASAP7_75t_L g938 ( .A(n_508), .Y(n_938) );
INVx8_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_SL g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_SL g616 ( .A(n_514), .Y(n_616) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g782 ( .A(n_518), .Y(n_782) );
BUFx3_ASAP7_75t_L g808 ( .A(n_518), .Y(n_808) );
BUFx2_ASAP7_75t_L g923 ( .A(n_518), .Y(n_923) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
BUFx3_ASAP7_75t_L g553 ( .A(n_521), .Y(n_553) );
BUFx2_ASAP7_75t_SL g587 ( .A(n_521), .Y(n_587) );
BUFx6f_ASAP7_75t_L g916 ( .A(n_521), .Y(n_916) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
BUFx2_ASAP7_75t_L g903 ( .A(n_524), .Y(n_903) );
INVx1_ASAP7_75t_L g1102 ( .A(n_524), .Y(n_1102) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx3_ASAP7_75t_L g597 ( .A(n_525), .Y(n_597) );
BUFx3_ASAP7_75t_L g626 ( .A(n_525), .Y(n_626) );
BUFx3_ASAP7_75t_L g755 ( .A(n_525), .Y(n_755) );
INVxp67_ASAP7_75t_L g558 ( .A(n_526), .Y(n_558) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g719 ( .A(n_529), .Y(n_719) );
INVx5_ASAP7_75t_SL g836 ( .A(n_529), .Y(n_836) );
INVx2_ASAP7_75t_SL g898 ( .A(n_529), .Y(n_898) );
INVx2_ASAP7_75t_L g1141 ( .A(n_529), .Y(n_1141) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx3_ASAP7_75t_L g566 ( .A(n_531), .Y(n_566) );
INVx2_ASAP7_75t_L g825 ( .A(n_531), .Y(n_825) );
INVx1_ASAP7_75t_L g650 ( .A(n_533), .Y(n_650) );
INVx1_ASAP7_75t_L g776 ( .A(n_533), .Y(n_776) );
BUFx4f_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g582 ( .A(n_535), .Y(n_582) );
XOR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_570), .Y(n_536) );
NAND4xp75_ASAP7_75t_L g537 ( .A(n_538), .B(n_544), .C(n_554), .D(n_567), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OA211x2_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B(n_549), .C(n_552), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_546), .A2(n_687), .B1(n_688), .B2(n_690), .Y(n_686) );
OA211x2_ASAP7_75t_L g939 ( .A1(n_546), .A2(n_940), .B(n_941), .C(n_942), .Y(n_939) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g648 ( .A(n_547), .Y(n_648) );
BUFx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g868 ( .A(n_548), .Y(n_868) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_557), .A2(n_823), .B1(n_824), .B2(n_826), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_557), .A2(n_565), .B1(n_957), .B2(n_958), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B1(n_564), .B2(n_565), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_568), .Y(n_580) );
INVx1_ASAP7_75t_L g778 ( .A(n_569), .Y(n_778) );
BUFx4f_ASAP7_75t_L g1094 ( .A(n_569), .Y(n_1094) );
INVx1_ASAP7_75t_L g632 ( .A(n_571), .Y(n_632) );
OAI22xp5_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_602), .B1(n_603), .B2(n_630), .Y(n_571) );
INVx1_ASAP7_75t_L g630 ( .A(n_572), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_588), .C(n_595), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_583), .Y(n_574) );
OAI21xp5_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_578), .B(n_579), .Y(n_575) );
OAI222xp33_ASAP7_75t_L g882 ( .A1(n_576), .A2(n_883), .B1(n_884), .B2(n_886), .C1(n_887), .C2(n_888), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g1005 ( .A1(n_576), .A2(n_1006), .B1(n_1007), .B2(n_1008), .C(n_1009), .Y(n_1005) );
OAI221xp5_ASAP7_75t_L g1090 ( .A1(n_576), .A2(n_776), .B1(n_1091), .B2(n_1092), .C(n_1093), .Y(n_1090) );
OAI221xp5_ASAP7_75t_L g1127 ( .A1(n_576), .A2(n_1128), .B1(n_1129), .B2(n_1130), .C(n_1131), .Y(n_1127) );
INVx2_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g652 ( .A(n_577), .Y(n_652) );
INVx2_ASAP7_75t_SL g1007 ( .A(n_580), .Y(n_1007) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .C(n_586), .Y(n_583) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .Y(n_588) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
INVx1_ASAP7_75t_L g675 ( .A(n_597), .Y(n_675) );
BUFx4f_ASAP7_75t_SL g705 ( .A(n_597), .Y(n_705) );
INVx1_ASAP7_75t_SL g725 ( .A(n_598), .Y(n_725) );
INVx3_ASAP7_75t_L g721 ( .A(n_601), .Y(n_721) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g629 ( .A(n_605), .Y(n_629) );
NAND3x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_617), .C(n_622), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_613), .Y(n_606) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_610), .B(n_611), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g1050 ( .A1(n_608), .A2(n_1051), .B(n_1052), .Y(n_1050) );
INVx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .Y(n_622) );
BUFx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
XNOR2xp5_ASAP7_75t_SL g634 ( .A(n_635), .B(n_765), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_680), .B2(n_764), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g679 ( .A(n_638), .Y(n_679) );
INVx1_ASAP7_75t_L g677 ( .A(n_639), .Y(n_677) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_663), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_641), .B(n_649), .C(n_656), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_646), .B2(n_647), .Y(n_641) );
OAI221xp5_ASAP7_75t_SL g840 ( .A1(n_643), .A2(n_647), .B1(n_841), .B2(n_842), .C(n_843), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_643), .A2(n_1002), .B1(n_1003), .B2(n_1004), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_643), .A2(n_1004), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g689 ( .A(n_644), .Y(n_689) );
BUFx3_ASAP7_75t_L g973 ( .A(n_644), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_647), .A2(n_1087), .B1(n_1088), .B2(n_1089), .Y(n_1086) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI222xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_652), .B2(n_653), .C1(n_654), .C2(n_655), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_658), .A2(n_661), .B1(n_875), .B2(n_876), .Y(n_874) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx3_ASAP7_75t_SL g965 ( .A(n_659), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_661), .A2(n_696), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_670), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g764 ( .A(n_680), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_709), .B1(n_762), .B2(n_763), .Y(n_680) );
INVx1_ASAP7_75t_L g762 ( .A(n_681), .Y(n_762) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_698), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_691), .C(n_694), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_688), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g1088 ( .A(n_689), .Y(n_1088) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_703), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_707), .Y(n_703) );
INVx1_ASAP7_75t_L g763 ( .A(n_709), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_733), .B1(n_760), .B2(n_761), .Y(n_709) );
INVx1_ASAP7_75t_L g761 ( .A(n_710), .Y(n_761) );
INVx1_ASAP7_75t_L g732 ( .A(n_711), .Y(n_732) );
AND4x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_718), .C(n_726), .D(n_730), .Y(n_711) );
INVx1_ASAP7_75t_SL g829 ( .A(n_713), .Y(n_829) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
BUFx3_ASAP7_75t_L g792 ( .A(n_714), .Y(n_792) );
INVx3_ASAP7_75t_L g855 ( .A(n_714), .Y(n_855) );
BUFx3_ASAP7_75t_L g1019 ( .A(n_714), .Y(n_1019) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g760 ( .A(n_735), .Y(n_760) );
AO22x2_ASAP7_75t_L g798 ( .A1(n_735), .A2(n_760), .B1(n_799), .B2(n_800), .Y(n_798) );
XOR2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_759), .Y(n_735) );
NAND2x1_ASAP7_75t_L g736 ( .A(n_737), .B(n_748), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .Y(n_737) );
OAI21xp5_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_740), .B(n_741), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .C(n_747), .Y(n_742) );
NOR2x1_ASAP7_75t_L g748 ( .A(n_749), .B(n_753), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g1045 ( .A(n_755), .Y(n_1045) );
INVx2_ASAP7_75t_L g1139 ( .A(n_758), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_797), .B2(n_798), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g796 ( .A(n_770), .Y(n_796) );
NAND3x1_ASAP7_75t_L g770 ( .A(n_771), .B(n_784), .C(n_789), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_780), .Y(n_771) );
OAI222xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_775), .B1(n_776), .B2(n_777), .C1(n_778), .C2(n_779), .Y(n_772) );
OAI21xp5_ASAP7_75t_SL g1029 ( .A1(n_773), .A2(n_1030), .B(n_1031), .Y(n_1029) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OAI221xp5_ASAP7_75t_L g869 ( .A1(n_776), .A2(n_870), .B1(n_871), .B2(n_872), .C(n_873), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_795), .Y(n_1144) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_813), .Y(n_800) );
NAND4xp75_ASAP7_75t_L g801 ( .A(n_802), .B(n_805), .C(n_809), .D(n_812), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AND2x2_ASAP7_75t_SL g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g1067 ( .A(n_815), .Y(n_1067) );
XOR2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_995), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B1(n_848), .B2(n_994), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_SL g847 ( .A(n_820), .Y(n_847) );
AND4x1_ASAP7_75t_L g820 ( .A(n_821), .B(n_832), .C(n_839), .D(n_844), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_827), .Y(n_821) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_827) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_838), .Y(n_832) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g994 ( .A(n_848), .Y(n_994) );
XOR2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_907), .Y(n_848) );
OAI22xp5_ASAP7_75t_SL g849 ( .A1(n_850), .A2(n_879), .B1(n_905), .B2(n_906), .Y(n_849) );
INVx2_ASAP7_75t_L g905 ( .A(n_850), .Y(n_905) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx2_ASAP7_75t_L g878 ( .A(n_852), .Y(n_878) );
AND2x2_ASAP7_75t_SL g852 ( .A(n_853), .B(n_863), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_859), .Y(n_853) );
INVx2_ASAP7_75t_L g895 ( .A(n_855), .Y(n_895) );
NOR3xp33_ASAP7_75t_L g863 ( .A(n_864), .B(n_869), .C(n_874), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_867), .A2(n_972), .B1(n_973), .B2(n_974), .Y(n_971) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_SL g1004 ( .A(n_868), .Y(n_1004) );
OAI21xp5_ASAP7_75t_SL g911 ( .A1(n_870), .A2(n_912), .B(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g906 ( .A(n_879), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_892), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_889), .Y(n_881) );
INVx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx4_ASAP7_75t_L g1033 ( .A(n_885), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_901), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_894), .B(n_899), .Y(n_893) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g907 ( .A1(n_908), .A2(n_932), .B1(n_992), .B2(n_993), .Y(n_907) );
INVx2_ASAP7_75t_L g992 ( .A(n_908), .Y(n_992) );
NAND2xp5_ASAP7_75t_SL g909 ( .A(n_910), .B(n_924), .Y(n_909) );
NOR2xp33_ASAP7_75t_SL g910 ( .A(n_911), .B(n_917), .Y(n_910) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_SL g915 ( .A(n_916), .Y(n_915) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_920), .C(n_922), .Y(n_917) );
NOR2x1_ASAP7_75t_L g924 ( .A(n_925), .B(n_928), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .Y(n_928) );
INVx1_ASAP7_75t_L g993 ( .A(n_932), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_948), .B1(n_990), .B2(n_991), .Y(n_932) );
INVx3_ASAP7_75t_SL g991 ( .A(n_933), .Y(n_991) );
XOR2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_947), .Y(n_933) );
NAND4xp75_ASAP7_75t_L g934 ( .A(n_935), .B(n_939), .C(n_943), .D(n_946), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
AND2x2_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g990 ( .A(n_948), .Y(n_990) );
XOR2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_976), .Y(n_948) );
XOR2xp5_ASAP7_75t_SL g949 ( .A(n_950), .B(n_975), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_951), .B(n_962), .Y(n_950) );
NOR3xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_956), .C(n_959), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_954), .Y(n_952) );
NOR3xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_967), .C(n_971), .Y(n_962) );
NAND4xp75_ASAP7_75t_L g977 ( .A(n_978), .B(n_981), .C(n_986), .D(n_989), .Y(n_977) );
AND2x2_ASAP7_75t_SL g978 ( .A(n_979), .B(n_980), .Y(n_978) );
AND2x2_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
AND2x2_ASAP7_75t_L g986 ( .A(n_987), .B(n_988), .Y(n_986) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B1(n_1024), .B2(n_1025), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1023 ( .A(n_999), .Y(n_1023) );
AND2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1013), .Y(n_999) );
NOR3xp33_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1005), .C(n_1010), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1017), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1016), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1020), .Y(n_1017) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
XNOR2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1047), .Y(n_1025) );
NAND3x2_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1039), .C(n_1042), .Y(n_1027) );
NOR2x1_ASAP7_75t_SL g1028 ( .A(n_1029), .B(n_1034), .Y(n_1028) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1032), .Y(n_1129) );
INVx3_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
NAND3xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .C(n_1038), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1041), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1046), .Y(n_1042) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
XOR2x2_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1066), .Y(n_1047) );
NAND2xp5_ASAP7_75t_SL g1048 ( .A(n_1049), .B(n_1057), .Y(n_1048) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1053), .Y(n_1049) );
NAND3xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .C(n_1056), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1062), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1061), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
INVx1_ASAP7_75t_SL g1069 ( .A(n_1070), .Y(n_1069) );
NOR2x1_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1075), .Y(n_1070) );
OR2x2_ASAP7_75t_SL g1150 ( .A(n_1071), .B(n_1076), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1074), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_1073), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1073), .B(n_1113), .Y(n_1116) );
CKINVDCx16_ASAP7_75t_R g1113 ( .A(n_1074), .Y(n_1113) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_1076), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1081), .Y(n_1079) );
OAI322xp33_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1109), .A3(n_1110), .B1(n_1114), .B2(n_1117), .C1(n_1118), .C2(n_1148), .Y(n_1082) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1084), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1098), .Y(n_1084) );
NOR3xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1090), .C(n_1095), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1104), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1103), .Y(n_1099) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1105), .B(n_1106), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx2_ASAP7_75t_SL g1147 ( .A(n_1122), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1135), .Y(n_1122) );
NOR3xp33_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1127), .C(n_1132), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1142), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1140), .Y(n_1136) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1145), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_1149), .Y(n_1148) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_1150), .Y(n_1149) );
endmodule