module fake_jpeg_1571_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.Y(n_60)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_43),
.B1(n_49),
.B2(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_57),
.B1(n_56),
.B2(n_55),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_37),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_51),
.B1(n_50),
.B2(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_69),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_42),
.C(n_45),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_82),
.B(n_0),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_55),
.B1(n_70),
.B2(n_41),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_96),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_65),
.B(n_60),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_24),
.B(n_32),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_41),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_79),
.B1(n_74),
.B2(n_76),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_51),
.B1(n_50),
.B2(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_93),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_1),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_97),
.C(n_90),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_108),
.B1(n_95),
.B2(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_2),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_82),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_114),
.B1(n_9),
.B2(n_11),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_125),
.B1(n_126),
.B2(n_114),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_104),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_97),
.B(n_33),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_124),
.C(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_6),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_7),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_12),
.B(n_14),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_99),
.C(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_133),
.C(n_123),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_117),
.C(n_122),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_123),
.A3(n_128),
.B1(n_120),
.B2(n_119),
.C1(n_107),
.C2(n_12),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_18),
.B(n_19),
.Y(n_138)
);

AOI31xp67_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_128),
.A3(n_107),
.B(n_20),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_138),
.C(n_25),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_26),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_14),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_136),
.C(n_15),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_16),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_16),
.Y(n_144)
);


endmodule