module fake_jpeg_29252_n_469 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_48),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_49),
.B(n_53),
.Y(n_118)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_10),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_10),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_56),
.B(n_59),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g130 ( 
.A(n_63),
.Y(n_130)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_66),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_30),
.B(n_11),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_76),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_30),
.B(n_11),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_96),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_82),
.B(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_11),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_89),
.Y(n_122)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_91),
.Y(n_105)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_97),
.B1(n_31),
.B2(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_29),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_98),
.B(n_92),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_40),
.B1(n_35),
.B2(n_33),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_102),
.A2(n_1),
.B(n_114),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_29),
.B1(n_47),
.B2(n_41),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_75),
.B1(n_68),
.B2(n_58),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_48),
.A2(n_40),
.B1(n_35),
.B2(n_43),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_108),
.A2(n_133),
.B1(n_137),
.B2(n_142),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_73),
.B(n_0),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_127),
.C(n_1),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_31),
.B1(n_41),
.B2(n_24),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_114),
.A2(n_117),
.B1(n_61),
.B2(n_55),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_116),
.A2(n_75),
.B(n_58),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_57),
.A2(n_43),
.B1(n_19),
.B2(n_28),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_54),
.A2(n_43),
.B1(n_28),
.B2(n_24),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_125),
.A2(n_128),
.B1(n_132),
.B2(n_153),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_28),
.C(n_23),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_66),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_60),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_67),
.A2(n_71),
.B1(n_78),
.B2(n_83),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_51),
.A2(n_21),
.B1(n_22),
.B2(n_4),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_65),
.A2(n_22),
.B1(n_12),
.B2(n_4),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_69),
.A2(n_22),
.B1(n_12),
.B2(n_4),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_90),
.A2(n_12),
.B1(n_16),
.B2(n_5),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_96),
.A2(n_87),
.B1(n_77),
.B2(n_70),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_88),
.A2(n_95),
.B1(n_94),
.B2(n_93),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_68),
.B(n_12),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_16),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_64),
.A2(n_91),
.B1(n_74),
.B2(n_62),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_98),
.B(n_97),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_155),
.B(n_162),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_156),
.A2(n_191),
.B1(n_130),
.B2(n_101),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_157),
.B(n_152),
.Y(n_211)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_100),
.B(n_32),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_58),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_178),
.Y(n_222)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_32),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_166),
.B(n_169),
.Y(n_236)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_168),
.A2(n_192),
.B1(n_139),
.B2(n_111),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_32),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_32),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_170),
.B(n_171),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_102),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_81),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_184),
.Y(n_234)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_174),
.A2(n_176),
.B(n_197),
.Y(n_246)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_99),
.A2(n_63),
.B(n_32),
.C(n_5),
.D(n_8),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_141),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_180),
.Y(n_237)
);

OR2x4_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_9),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_135),
.Y(n_221)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_105),
.A2(n_9),
.B(n_13),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_145),
.B(n_123),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_98),
.B(n_0),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_13),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_13),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_144),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_199),
.Y(n_242)
);

AO22x1_ASAP7_75t_SL g189 ( 
.A1(n_104),
.A2(n_0),
.B1(n_1),
.B2(n_15),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_130),
.B1(n_115),
.B2(n_119),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_126),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_112),
.A2(n_14),
.B1(n_15),
.B2(n_0),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_112),
.B(n_0),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_203),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_107),
.B(n_1),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_201),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_107),
.B(n_104),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_202),
.A2(n_109),
.B1(n_121),
.B2(n_182),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_105),
.B(n_127),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_136),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_124),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_126),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_205),
.B(n_130),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_117),
.B1(n_144),
.B2(n_123),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_209),
.A2(n_183),
.B(n_181),
.C(n_192),
.D(n_176),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_210),
.A2(n_218),
.B1(n_227),
.B2(n_155),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_211),
.B(n_225),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_168),
.A2(n_198),
.B1(n_177),
.B2(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_217),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_220),
.B(n_200),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_221),
.B(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_204),
.B(n_120),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_139),
.B1(n_119),
.B2(n_115),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_198),
.A2(n_111),
.B1(n_131),
.B2(n_120),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_124),
.B1(n_138),
.B2(n_121),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_178),
.B(n_138),
.C(n_135),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_167),
.C(n_202),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_248),
.Y(n_267)
);

AO21x2_ASAP7_75t_L g249 ( 
.A1(n_206),
.A2(n_174),
.B(n_186),
.Y(n_249)
);

AO22x1_ASAP7_75t_SL g301 ( 
.A1(n_249),
.A2(n_229),
.B1(n_219),
.B2(n_226),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_161),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_256),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_189),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_252),
.A2(n_214),
.B(n_244),
.Y(n_318)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_156),
.B1(n_177),
.B2(n_201),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_262),
.B1(n_242),
.B2(n_216),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_209),
.A2(n_205),
.B1(n_154),
.B2(n_158),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_255),
.A2(n_258),
.B1(n_281),
.B2(n_237),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_188),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_184),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_264),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_218),
.B1(n_160),
.B2(n_163),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_173),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_272),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_172),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_268),
.C(n_271),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_261),
.A2(n_277),
.B(n_237),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_221),
.A2(n_201),
.B1(n_199),
.B2(n_155),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_184),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_266),
.A2(n_270),
.B1(n_276),
.B2(n_286),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_172),
.C(n_162),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_162),
.B1(n_200),
.B2(n_189),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_212),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_196),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_275),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_286),
.C(n_220),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_240),
.B(n_165),
.Y(n_275)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_109),
.A3(n_180),
.B1(n_179),
.B2(n_175),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_232),
.B(n_193),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_278),
.B(n_280),
.Y(n_298)
);

BUFx4f_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_279),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_224),
.B(n_195),
.Y(n_280)
);

OAI22x1_ASAP7_75t_SL g281 ( 
.A1(n_246),
.A2(n_179),
.B1(n_190),
.B2(n_194),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_179),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_283),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_109),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_208),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_207),
.B(n_226),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_285),
.B(n_214),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_247),
.C(n_216),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_288),
.A2(n_292),
.B1(n_294),
.B2(n_302),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_289),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_250),
.A2(n_246),
.B1(n_243),
.B2(n_216),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_282),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_295),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_243),
.B1(n_242),
.B2(n_234),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_279),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_279),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_296),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_301),
.A2(n_277),
.B(n_283),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_234),
.B1(n_219),
.B2(n_229),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_269),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_304),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_284),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_315),
.Y(n_330)
);

NOR2x1p5_ASAP7_75t_SL g309 ( 
.A(n_281),
.B(n_244),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_230),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_314),
.B1(n_319),
.B2(n_252),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_272),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_312),
.A2(n_308),
.B1(n_294),
.B2(n_298),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_266),
.A2(n_276),
.B1(n_249),
.B2(n_270),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_317),
.A2(n_223),
.B(n_318),
.Y(n_347)
);

A2O1A1O1Ixp25_ASAP7_75t_L g339 ( 
.A1(n_318),
.A2(n_263),
.B(n_275),
.C(n_257),
.D(n_264),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_249),
.A2(n_230),
.B1(n_245),
.B2(n_233),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_228),
.C(n_215),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_274),
.C(n_262),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_321),
.A2(n_329),
.B1(n_332),
.B2(n_346),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_325),
.C(n_333),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_319),
.A2(n_252),
.B1(n_267),
.B2(n_249),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_314),
.B1(n_310),
.B2(n_293),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_290),
.B(n_268),
.C(n_271),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_309),
.A2(n_249),
.B1(n_267),
.B2(n_263),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_350),
.B1(n_301),
.B2(n_313),
.Y(n_356)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_301),
.Y(n_352)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_337),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_339),
.A2(n_347),
.B(n_348),
.Y(n_363)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_300),
.Y(n_340)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_273),
.C(n_228),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_345),
.C(n_316),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_342),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_304),
.B(n_261),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_343),
.Y(n_351)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_288),
.B(n_213),
.C(n_215),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_312),
.A2(n_245),
.B1(n_213),
.B2(n_223),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_292),
.B(n_302),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_303),
.Y(n_349)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_320),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_333),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_327),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_354),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_356),
.A2(n_359),
.B1(n_361),
.B2(n_377),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_329),
.A2(n_301),
.B1(n_308),
.B2(n_306),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_364),
.B1(n_367),
.B2(n_371),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_334),
.A2(n_313),
.B1(n_307),
.B2(n_311),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_350),
.A2(n_307),
.B1(n_298),
.B2(n_315),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_369),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_321),
.A2(n_306),
.B1(n_287),
.B2(n_305),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_332),
.A2(n_287),
.B1(n_291),
.B2(n_295),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_331),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_328),
.B(n_297),
.Y(n_370)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_342),
.A2(n_328),
.B1(n_347),
.B2(n_348),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_297),
.Y(n_372)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_323),
.C(n_337),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_336),
.A2(n_291),
.B1(n_296),
.B2(n_346),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_374),
.A2(n_322),
.B1(n_338),
.B2(n_349),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_343),
.A2(n_336),
.B1(n_331),
.B2(n_345),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_371),
.A2(n_336),
.B(n_338),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_380),
.B(n_386),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_381),
.B(n_387),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_382),
.A2(n_360),
.B1(n_366),
.B2(n_368),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_341),
.Y(n_385)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_335),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_325),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_364),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_391),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_363),
.A2(n_322),
.B(n_323),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_372),
.B(n_374),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_339),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_399),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_370),
.Y(n_392)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_392),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_398),
.C(n_354),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_356),
.A2(n_359),
.B1(n_376),
.B2(n_352),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_395),
.A2(n_358),
.B1(n_367),
.B2(n_355),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_326),
.C(n_340),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_344),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_402),
.C(n_393),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_362),
.C(n_377),
.Y(n_402)
);

XOR2x1_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_363),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_404),
.B(n_414),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_406),
.A2(n_384),
.B(n_397),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_361),
.B1(n_355),
.B2(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_408),
.A2(n_394),
.B1(n_383),
.B2(n_396),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_379),
.A2(n_358),
.B1(n_360),
.B2(n_366),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_380),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_397),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_396),
.Y(n_412)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_412),
.Y(n_423)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_384),
.Y(n_413)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_413),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_390),
.B(n_375),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_378),
.A2(n_326),
.B1(n_375),
.B2(n_382),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_416),
.B(n_395),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_426),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_419),
.B(n_411),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_420),
.A2(n_383),
.B(n_400),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_427),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_410),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_403),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_415),
.B(n_379),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_394),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_399),
.C(n_387),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_411),
.C(n_402),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_431),
.B(n_406),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_435),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_437),
.B(n_440),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_405),
.Y(n_438)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_420),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_405),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_441),
.A2(n_381),
.B(n_417),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_409),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_442),
.B(n_443),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_408),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_427),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_448),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_434),
.A2(n_428),
.B1(n_404),
.B2(n_412),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_449),
.B(n_439),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_423),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_452),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_437),
.C(n_436),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_444),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_454),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_442),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_458),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_400),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_459),
.A2(n_455),
.B(n_457),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_453),
.A2(n_449),
.B(n_429),
.Y(n_461)
);

AOI31xp33_ASAP7_75t_L g464 ( 
.A1(n_461),
.A2(n_452),
.A3(n_424),
.B(n_414),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_463),
.A2(n_464),
.B(n_462),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_463),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_466),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_467),
.B(n_460),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_SL g469 ( 
.A(n_468),
.B(n_424),
.Y(n_469)
);


endmodule