module fake_jpeg_15874_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_19),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_29),
.B(n_37),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_6),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_1),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_69),
.Y(n_77)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_54),
.B1(n_46),
.B2(n_49),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_72),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_46),
.B1(n_49),
.B2(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_62),
.B1(n_61),
.B2(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_47),
.Y(n_84)
);

OA22x2_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_53),
.B1(n_45),
.B2(n_56),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_90),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_102),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_4),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_60),
.C(n_44),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_4),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_100),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_82),
.B1(n_60),
.B2(n_44),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_101),
.B1(n_9),
.B2(n_13),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_5),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_86),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_110),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_112),
.B1(n_95),
.B2(n_91),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_25),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_98),
.B(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_109),
.B1(n_93),
.B2(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_122),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_109),
.B1(n_104),
.B2(n_89),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_123),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_30),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_122),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_129),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_125),
.Y(n_130)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_131),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_132),
.B1(n_125),
.B2(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_28),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_31),
.B(n_14),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_32),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_27),
.B(n_15),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_33),
.B(n_16),
.C(n_18),
.D(n_21),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_42),
.B1(n_23),
.B2(n_35),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_140),
.Y(n_141)
);


endmodule