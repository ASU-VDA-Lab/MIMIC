module fake_jpeg_9437_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

CKINVDCx9p33_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_1),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_3),
.B(n_4),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_3),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_22),
.Y(n_68)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_15),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_16),
.B1(n_13),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_21),
.B1(n_23),
.B2(n_15),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_49),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_28),
.B1(n_37),
.B2(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_63),
.B1(n_66),
.B2(n_45),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_47),
.B(n_50),
.C(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_60),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_16),
.B1(n_36),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_36),
.B1(n_27),
.B2(n_31),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_31),
.B1(n_36),
.B2(n_27),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_24),
.B(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_44),
.B1(n_39),
.B2(n_42),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_22),
.B1(n_25),
.B2(n_14),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_24),
.Y(n_81)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_24),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_46),
.B1(n_42),
.B2(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_58),
.B1(n_52),
.B2(n_68),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_25),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_35),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_69),
.B1(n_67),
.B2(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_90),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_93),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_76),
.C(n_74),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_67),
.B1(n_14),
.B2(n_19),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_4),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_82),
.B(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_73),
.B(n_75),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_92),
.B(n_90),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_104),
.C(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_91),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_76),
.C(n_72),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_107),
.B(n_92),
.Y(n_113)
);

FAx1_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_83),
.CI(n_70),
.CON(n_107),
.SN(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_19),
.C(n_14),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_116),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_107),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_97),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_105),
.C(n_19),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_97),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_6),
.C(n_7),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_112),
.B1(n_115),
.B2(n_8),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_125),
.B(n_9),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_11),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_118),
.C(n_117),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_9),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_124),
.B(n_10),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_10),
.B(n_131),
.Y(n_133)
);

BUFx24_ASAP7_75t_SL g134 ( 
.A(n_133),
.Y(n_134)
);


endmodule