module fake_jpeg_13768_n_199 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_SL g74 ( 
.A(n_38),
.B(n_8),
.C(n_0),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_2),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_89),
.Y(n_103)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_75),
.B1(n_50),
.B2(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_102),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_75),
.B1(n_50),
.B2(n_66),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_51),
.B1(n_76),
.B2(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_81),
.B1(n_62),
.B2(n_57),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_61),
.B1(n_70),
.B2(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_104),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_70),
.B1(n_52),
.B2(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_59),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_62),
.B1(n_73),
.B2(n_71),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_123),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_116),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_60),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_12),
.B(n_14),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_142),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_65),
.B1(n_79),
.B2(n_6),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_143),
.B1(n_10),
.B2(n_11),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_79),
.C(n_25),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_145),
.B(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_130),
.C(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_9),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_158),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_163),
.B1(n_168),
.B2(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_10),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_164),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_151),
.B1(n_147),
.B2(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_12),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_152),
.B1(n_154),
.B2(n_140),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_175),
.A2(n_178),
.B1(n_172),
.B2(n_156),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_140),
.A3(n_133),
.B1(n_131),
.B2(n_142),
.C1(n_23),
.C2(n_24),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_21),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_162),
.C(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_187),
.C(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_181),
.C(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_191),
.A2(n_180),
.B1(n_173),
.B2(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_192),
.B(n_167),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_167),
.B(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_26),
.B(n_32),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_34),
.B(n_39),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_42),
.Y(n_199)
);


endmodule