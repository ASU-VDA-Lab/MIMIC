module fake_jpeg_978_n_229 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_12),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_53),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_0),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_71),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_61),
.B1(n_78),
.B2(n_76),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_93),
.B1(n_74),
.B2(n_59),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_94),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_78),
.B1(n_71),
.B2(n_76),
.Y(n_93)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_59),
.B1(n_77),
.B2(n_68),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_55),
.B1(n_70),
.B2(n_62),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_95),
.A2(n_87),
.B1(n_62),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_118),
.B1(n_85),
.B2(n_91),
.Y(n_126)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_81),
.C(n_87),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_115),
.C(n_74),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_72),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_114),
.Y(n_127)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_81),
.B1(n_85),
.B2(n_63),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_109),
.B1(n_75),
.B2(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_117),
.Y(n_142)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_64),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_60),
.C(n_64),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_67),
.CI(n_63),
.CON(n_117),
.SN(n_117)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_56),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_5),
.Y(n_152)
);

OR2x4_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_67),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_75),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_134),
.B1(n_141),
.B2(n_1),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_7),
.Y(n_155)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_60),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_7),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_79),
.C(n_69),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.C(n_8),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_65),
.C(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_75),
.B(n_4),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_139),
.Y(n_157)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_140),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_75),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_145),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_147),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_116),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_148),
.Y(n_178)
);

XOR2x2_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_25),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_29),
.B1(n_49),
.B2(n_48),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_151),
.A2(n_121),
.B1(n_15),
.B2(n_16),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_163),
.Y(n_172)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_11),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_13),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_161),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_170),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_154),
.A2(n_137),
.B(n_132),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_174),
.B(n_177),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_140),
.B1(n_133),
.B2(n_17),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_151),
.B1(n_158),
.B2(n_162),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_14),
.B(n_15),
.C(n_18),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_36),
.Y(n_184)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_157),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_144),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_148),
.C(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_179),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_191),
.B1(n_193),
.B2(n_177),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_180),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_196),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_173),
.A2(n_164),
.B1(n_162),
.B2(n_20),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_14),
.B1(n_19),
.B2(n_20),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_37),
.B1(n_46),
.B2(n_22),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_175),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_170),
.B(n_186),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_202),
.A2(n_194),
.B(n_172),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_167),
.C(n_178),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_205),
.C(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_178),
.C(n_184),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_209),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_189),
.C(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_183),
.C(n_172),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_211),
.B(n_201),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_208),
.A2(n_191),
.B(n_193),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_174),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_200),
.A2(n_19),
.B1(n_21),
.B2(n_23),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

AOI321xp33_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_220),
.A3(n_212),
.B1(n_32),
.B2(n_33),
.C(n_38),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_205),
.C(n_31),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_222),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_218),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_42),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_221),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_203),
.B(n_45),
.C(n_50),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_43),
.Y(n_229)
);


endmodule