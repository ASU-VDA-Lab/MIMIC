module fake_jpeg_20153_n_267 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_267);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_27),
.B(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_44),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_12),
.B1(n_21),
.B2(n_19),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_42),
.B1(n_34),
.B2(n_30),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_12),
.B1(n_19),
.B2(n_15),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_29),
.C(n_33),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_60),
.B1(n_63),
.B2(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_27),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_41),
.B(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_29),
.B1(n_39),
.B2(n_30),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_29),
.C(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_37),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_43),
.B1(n_32),
.B2(n_12),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_67),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_27),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_47),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_26),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_39),
.B1(n_40),
.B2(n_35),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_78),
.B1(n_61),
.B2(n_50),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_77),
.B1(n_79),
.B2(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_14),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_68),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_61),
.C(n_54),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_68),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_98),
.B1(n_68),
.B2(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_60),
.B1(n_63),
.B2(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_94),
.B1(n_97),
.B2(n_99),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_32),
.B(n_18),
.C(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_52),
.B1(n_49),
.B2(n_48),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_32),
.B1(n_40),
.B2(n_33),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_79),
.B1(n_77),
.B2(n_72),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_59),
.B1(n_31),
.B2(n_28),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_59),
.B1(n_31),
.B2(n_28),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_82),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_105),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_112),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_81),
.B1(n_36),
.B2(n_65),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_68),
.B1(n_74),
.B2(n_65),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_90),
.B1(n_100),
.B2(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_113),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_116),
.C(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_26),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_26),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_95),
.B1(n_36),
.B2(n_46),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_99),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_91),
.B(n_86),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_135),
.B(n_143),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_131),
.B1(n_142),
.B2(n_144),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_128),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_96),
.C(n_91),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.C(n_36),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_136),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_116),
.C(n_117),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_92),
.B1(n_36),
.B2(n_37),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_46),
.B1(n_18),
.B2(n_23),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_101),
.A2(n_7),
.B(n_1),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_70),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_139),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_85),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_7),
.B(n_2),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_70),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_139),
.A2(n_112),
.B1(n_114),
.B2(n_104),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_150),
.B1(n_159),
.B2(n_163),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_26),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_161),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_46),
.B1(n_31),
.B2(n_28),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_28),
.C(n_26),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_123),
.C(n_140),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_156),
.B1(n_162),
.B2(n_8),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_156)
);

XOR2x2_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_24),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_143),
.B(n_132),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_124),
.B1(n_130),
.B2(n_138),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_24),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_9),
.B(n_3),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_144),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_20),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_174),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_153),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_126),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_25),
.Y(n_185)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_8),
.Y(n_186)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_22),
.B1(n_0),
.B2(n_5),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_162),
.B1(n_154),
.B2(n_155),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_149),
.C(n_151),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_201),
.C(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_181),
.A2(n_184),
.B1(n_172),
.B2(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_205),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_187),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_146),
.B1(n_166),
.B2(n_163),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_213),
.C(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_172),
.B(n_179),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_216),
.B(n_218),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_187),
.C(n_178),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_147),
.C(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_176),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_220),
.B(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_192),
.C(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_230),
.C(n_217),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_167),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_198),
.B(n_180),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_205),
.C(n_202),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_212),
.B1(n_206),
.B2(n_219),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_242),
.C(n_221),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_185),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_238),
.B(n_232),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_177),
.B1(n_188),
.B2(n_189),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_177),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_225),
.B(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_20),
.C(n_0),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_247),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_221),
.B(n_5),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_233),
.B(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_4),
.C(n_5),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_250),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_253),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_246),
.B(n_240),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_240),
.B(n_242),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_4),
.B(n_6),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_251),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_257),
.B(n_254),
.Y(n_260)
);

NAND4xp25_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_261),
.C(n_6),
.D(n_7),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_9),
.B(n_10),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_9),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_264),
.A2(n_9),
.B(n_10),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_10),
.C(n_11),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);


endmodule