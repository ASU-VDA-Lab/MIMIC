module real_jpeg_11770_n_17 (n_5, n_4, n_8, n_0, n_12, n_326, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_326;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_37),
.B1(n_59),
.B2(n_64),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_5),
.A2(n_59),
.B1(n_64),
.B2(n_146),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_146),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_146),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_6),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_6),
.B(n_59),
.C(n_63),
.Y(n_170)
);

NAND2x1_ASAP7_75t_SL g174 ( 
.A(n_6),
.B(n_31),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_6),
.A2(n_137),
.B(n_182),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_27),
.B(n_30),
.C(n_209),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_6),
.B(n_52),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_41),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_7),
.A2(n_51),
.B1(n_59),
.B2(n_64),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_75),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_75),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_9),
.A2(n_59),
.B1(n_64),
.B2(n_75),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_10),
.A2(n_59),
.B1(n_64),
.B2(n_178),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_178),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_178),
.Y(n_280)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_12),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_83),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_12),
.A2(n_59),
.B1(n_64),
.B2(n_83),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_83),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_112),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_14),
.A2(n_59),
.B1(n_64),
.B2(n_112),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_112),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_43),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_15),
.A2(n_43),
.B1(n_59),
.B2(n_64),
.Y(n_270)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_90),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_76),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_24),
.A2(n_31),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_24),
.B(n_216),
.Y(n_230)
);

NOR2x1_ASAP7_75t_R g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_26),
.A2(n_32),
.B(n_166),
.Y(n_209)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_30),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_28),
.B(n_47),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g265 ( 
.A1(n_30),
.A2(n_42),
.A3(n_48),
.B1(n_253),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_31),
.B(n_216),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_32),
.A2(n_33),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_33),
.B(n_170),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_45),
.B1(n_46),
.B2(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_42),
.A2(n_45),
.B(n_166),
.C(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_44),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_46),
.B1(n_74),
.B2(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_45),
.A2(n_145),
.B(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_45),
.A2(n_46),
.B1(n_145),
.B2(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_46),
.A2(n_82),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_46),
.B(n_111),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_46),
.A2(n_109),
.B(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_69),
.C(n_73),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_69),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_81),
.C(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_80),
.B1(n_85),
.B2(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_65),
.B(n_67),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_65),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_57),
.A2(n_65),
.B1(n_105),
.B2(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_57),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_57),
.A2(n_65),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_57),
.A2(n_65),
.B1(n_141),
.B2(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_58),
.A2(n_68),
.B1(n_107),
.B2(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_58),
.A2(n_177),
.B(n_179),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_58),
.B(n_166),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_58),
.A2(n_179),
.B(n_258),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_64),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_64),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_65),
.B(n_168),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_72),
.B1(n_87),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_70),
.A2(n_72),
.B1(n_116),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_70),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_70),
.A2(n_72),
.B1(n_229),
.B2(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_70),
.A2(n_215),
.B(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_72),
.A2(n_229),
.B(n_230),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_72),
.A2(n_143),
.B(n_230),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.C(n_84),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_77),
.A2(n_81),
.B1(n_122),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_81),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_85),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_154),
.B(n_322),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_149),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_124),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_93),
.B(n_124),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_113),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_94),
.B(n_114),
.C(n_119),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B(n_108),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_96),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_98),
.B1(n_108),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_97),
.A2(n_98),
.B1(n_103),
.B2(n_104),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_99),
.A2(n_100),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_99),
.B(n_183),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_99),
.A2(n_100),
.B1(n_136),
.B2(n_270),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_100),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_115),
.B(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_118),
.A2(n_165),
.B(n_167),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_118),
.A2(n_167),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_131),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_130),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_131),
.B(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_142),
.C(n_144),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_132),
.A2(n_133),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_134),
.A2(n_139),
.B1(n_140),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_134),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_137),
.A2(n_138),
.B1(n_211),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_137),
.A2(n_138),
.B1(n_236),
.B2(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_138),
.A2(n_188),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_166),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_138),
.A2(n_196),
.B(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_142),
.B(n_144),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_148),
.B(n_251),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_149),
.A2(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_150),
.B(n_153),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_316),
.B(n_321),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_304),
.B(n_315),
.Y(n_155)
);

OAI321xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_272),
.A3(n_297),
.B1(n_302),
.B2(n_303),
.C(n_326),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_245),
.B(n_271),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_223),
.B(n_244),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_204),
.B(n_222),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_184),
.B(n_203),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_171),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_162),
.B(n_171),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_164),
.B1(n_169),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_176),
.C(n_180),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_192),
.B(n_202),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_190),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_197),
.B(n_201),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_206),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_217),
.C(n_221),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_210),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_224),
.B(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_237),
.B2(n_238),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_240),
.C(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_232),
.C(n_235),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_246),
.B(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_261),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_262),
.C(n_263),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_254),
.B2(n_260),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_255),
.C(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_287),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_287),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.C(n_286),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_274),
.A2(n_275),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_281),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_281),
.C(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_286),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_296),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_291),
.C(n_296),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_294),
.C(n_295),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_314),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_314),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_309),
.C(n_310),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);


endmodule