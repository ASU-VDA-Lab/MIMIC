module fake_jpeg_6070_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_48),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_31),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_50),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_17),
.B1(n_24),
.B2(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_21),
.B1(n_18),
.B2(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_16),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_24),
.B1(n_29),
.B2(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_16),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_24),
.B1(n_29),
.B2(n_33),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_75),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_23),
.C(n_27),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_82),
.B(n_32),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_79),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_39),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_23),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_45),
.B(n_61),
.C(n_43),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_86),
.B(n_37),
.Y(n_123)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_88),
.Y(n_110)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_27),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_27),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_54),
.B1(n_56),
.B2(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_77),
.B1(n_59),
.B2(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_43),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_102),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_99),
.B(n_50),
.Y(n_116)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_51),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_38),
.B1(n_51),
.B2(n_35),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_107),
.B1(n_70),
.B2(n_76),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_75),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_19),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_40),
.B1(n_37),
.B2(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_114),
.B1(n_122),
.B2(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_112),
.Y(n_135)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_121),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_89),
.B(n_92),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_37),
.B1(n_40),
.B2(n_49),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_128),
.B1(n_86),
.B2(n_87),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_129),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_77),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_73),
.Y(n_127)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_92),
.B1(n_90),
.B2(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_97),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_106),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_137),
.C(n_138),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_139),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_142),
.B(n_144),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_99),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_91),
.C(n_93),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_100),
.B(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_150),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_86),
.B(n_96),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_96),
.B(n_68),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_68),
.C(n_73),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_148),
.C(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_147),
.B(n_151),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_58),
.C(n_40),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_116),
.B1(n_129),
.B2(n_121),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_169),
.B1(n_146),
.B2(n_139),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_166),
.B(n_168),
.Y(n_179)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx6_ASAP7_75t_SL g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_108),
.B1(n_97),
.B2(n_38),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_136),
.C(n_141),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_172),
.C(n_133),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_58),
.C(n_101),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_25),
.B(n_22),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_180),
.C(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_134),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_58),
.C(n_38),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_25),
.B(n_22),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_186),
.B1(n_166),
.B2(n_169),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_25),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_22),
.B1(n_15),
.B2(n_2),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_15),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_197),
.B(n_198),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_15),
.B(n_1),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_203),
.Y(n_216)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_155),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_171),
.B1(n_156),
.B2(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_175),
.B1(n_162),
.B2(n_178),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_SL g208 ( 
.A(n_206),
.B(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_185),
.C(n_181),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_215),
.B(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_160),
.C(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_213),
.C(n_214),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_180),
.C(n_172),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_200),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_0),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_212),
.B(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_226),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_206),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_205),
.B1(n_201),
.B2(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_227),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_3),
.B(n_4),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_218),
.C(n_209),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_232),
.C(n_233),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_6),
.B(n_8),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_225),
.C(n_224),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_0),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_3),
.B(n_5),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_3),
.CI(n_5),
.CON(n_241),
.SN(n_241)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_234),
.C(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_240),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_6),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_6),
.B(n_7),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_44),
.C2(n_247),
.Y(n_248)
);

AO221x1_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_240),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_9),
.B(n_10),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.C(n_245),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_9),
.B(n_11),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_44),
.Y(n_252)
);


endmodule