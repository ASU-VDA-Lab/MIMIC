module fake_netlist_1_427_n_671 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_671);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_671;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g75 ( .A(n_69), .Y(n_75) );
INVxp33_ASAP7_75t_SL g76 ( .A(n_7), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_47), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_23), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_13), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_58), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_63), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_46), .B(n_62), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_50), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_42), .Y(n_85) );
INVx1_ASAP7_75t_SL g86 ( .A(n_26), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_72), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_10), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_45), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_34), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_30), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_20), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_29), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_28), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_9), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_48), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_18), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_37), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_14), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_9), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_53), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_18), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_61), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_15), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_54), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_60), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_52), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_36), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_33), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_6), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_21), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_6), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_51), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_19), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_68), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_2), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_112), .Y(n_124) );
NAND2xp33_ASAP7_75t_SL g125 ( .A(n_75), .B(n_0), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_119), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_93), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_114), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_77), .B(n_1), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_101), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_76), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_102), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_92), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_108), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_108), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_110), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_108), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_109), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_91), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_109), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_77), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_78), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_110), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_78), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_79), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_91), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_98), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_105), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_110), .B(n_1), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_80), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_86), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_79), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_83), .B(n_2), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_91), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_81), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_84), .Y(n_161) );
NAND2x1_ASAP7_75t_L g162 ( .A(n_83), .B(n_3), .Y(n_162) );
INVx4_ASAP7_75t_SL g163 ( .A(n_130), .Y(n_163) );
BUFx2_ASAP7_75t_L g164 ( .A(n_126), .Y(n_164) );
NAND2x1p5_ASAP7_75t_L g165 ( .A(n_158), .B(n_89), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_149), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_134), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_135), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_140), .B(n_89), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_156), .B(n_100), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_157), .B(n_103), .Y(n_172) );
AND3x1_ASAP7_75t_L g173 ( .A(n_158), .B(n_121), .C(n_94), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
OAI22xp33_ASAP7_75t_SL g176 ( .A1(n_162), .A2(n_121), .B1(n_94), .B2(n_97), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_144), .B(n_145), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_162), .B(n_97), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_144), .B(n_100), .Y(n_181) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_127), .B(n_86), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_134), .Y(n_185) );
OR2x2_ASAP7_75t_SL g186 ( .A(n_152), .B(n_115), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_151), .B(n_104), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_148), .B(n_104), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_128), .B(n_120), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_124), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_132), .B(n_120), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_122), .Y(n_195) );
AND2x6_ASAP7_75t_L g196 ( .A(n_161), .B(n_120), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_154), .Y(n_197) );
BUFx10_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_154), .B(n_117), .Y(n_199) );
INVxp33_ASAP7_75t_L g200 ( .A(n_155), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_134), .Y(n_201) );
NAND2xp33_ASAP7_75t_L g202 ( .A(n_155), .B(n_110), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_134), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_122), .Y(n_204) );
AO22x2_ASAP7_75t_L g205 ( .A1(n_161), .A2(n_99), .B1(n_117), .B2(n_107), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_123), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_123), .B(n_96), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_131), .Y(n_208) );
OR2x2_ASAP7_75t_SL g209 ( .A(n_125), .B(n_107), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_131), .B(n_96), .Y(n_210) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_136), .Y(n_211) );
AO22x2_ASAP7_75t_L g212 ( .A1(n_129), .A2(n_115), .B1(n_116), .B2(n_95), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_136), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_142), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_142), .Y(n_215) );
NAND2x1p5_ASAP7_75t_L g216 ( .A(n_153), .B(n_95), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_150), .Y(n_218) );
OR2x2_ASAP7_75t_SL g219 ( .A(n_137), .B(n_84), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_159), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_137), .B(n_106), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_175), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_165), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_175), .B(n_90), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_200), .A2(n_159), .B1(n_139), .B2(n_143), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_199), .B(n_143), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_196), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_170), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_211), .B(n_111), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_165), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_173), .B(n_141), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_183), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_196), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_199), .B(n_141), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_196), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_174), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_214), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_177), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_169), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_196), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_218), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_211), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_212), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_221), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_173), .B(n_139), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_169), .A2(n_87), .B1(n_85), .B2(n_106), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_213), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_212), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_206), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_208), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_187), .B(n_111), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_191), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_197), .B(n_85), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_219), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_192), .B(n_194), .Y(n_263) );
BUFx4f_ASAP7_75t_L g264 ( .A(n_180), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_167), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_188), .B(n_116), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_181), .B(n_88), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_172), .B(n_3), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_205), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_167), .Y(n_270) );
NOR3xp33_ASAP7_75t_SL g271 ( .A(n_171), .B(n_88), .C(n_82), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_181), .B(n_118), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_190), .Y(n_273) );
INVx5_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
BUFx10_ASAP7_75t_L g275 ( .A(n_168), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_215), .Y(n_276) );
AND3x1_ASAP7_75t_SL g277 ( .A(n_209), .B(n_4), .C(n_5), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_179), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_198), .Y(n_279) );
INVx3_ASAP7_75t_L g280 ( .A(n_184), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_184), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_215), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_176), .B(n_118), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_189), .Y(n_284) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_182), .B(n_118), .C(n_113), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_242), .B(n_176), .Y(n_286) );
AOI22xp33_ASAP7_75t_SL g287 ( .A1(n_249), .A2(n_205), .B1(n_180), .B2(n_190), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
AND2x6_ASAP7_75t_L g289 ( .A(n_239), .B(n_222), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_224), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_224), .Y(n_291) );
OAI21xp33_ASAP7_75t_L g292 ( .A1(n_243), .A2(n_210), .B(n_207), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_239), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_245), .B(n_189), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_245), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_229), .A2(n_207), .B(n_222), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_223), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_225), .B(n_113), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_273), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_273), .B(n_216), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_239), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
NOR2x1_ASAP7_75t_L g306 ( .A(n_268), .B(n_113), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_249), .A2(n_186), .B1(n_216), .B2(n_110), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_240), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_240), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_229), .A2(n_202), .B(n_138), .Y(n_311) );
INVx5_ASAP7_75t_L g312 ( .A(n_239), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_225), .B(n_163), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_260), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_238), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_243), .A2(n_198), .B1(n_163), .B2(n_146), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_275), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_264), .B(n_163), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_234), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_231), .A2(n_138), .B(n_146), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_228), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_239), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_231), .A2(n_138), .B(n_146), .Y(n_323) );
INVx5_ASAP7_75t_L g324 ( .A(n_244), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_244), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_254), .Y(n_326) );
CKINVDCx8_ASAP7_75t_R g327 ( .A(n_235), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_275), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_254), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_268), .B(n_4), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_235), .B(n_5), .Y(n_331) );
INVx2_ASAP7_75t_SL g332 ( .A(n_264), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_233), .B(n_7), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_288), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_317), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_295), .A2(n_256), .B1(n_269), .B2(n_246), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_304), .B(n_312), .Y(n_337) );
AOI22xp33_ASAP7_75t_SL g338 ( .A1(n_290), .A2(n_251), .B1(n_262), .B2(n_235), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_298), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_310), .B(n_262), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_287), .A2(n_250), .B1(n_246), .B2(n_258), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_321), .B(n_252), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_296), .A2(n_258), .B(n_236), .Y(n_343) );
NAND2xp33_ASAP7_75t_SL g344 ( .A(n_322), .B(n_230), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_287), .A2(n_252), .B1(n_226), .B2(n_264), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_305), .B(n_252), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_326), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_297), .A2(n_283), .B1(n_276), .B2(n_282), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_291), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_315), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_328), .B(n_230), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_302), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_297), .B(n_276), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_322), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_286), .B(n_282), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_286), .A2(n_266), .B1(n_285), .B2(n_236), .Y(n_362) );
INVx6_ASAP7_75t_L g363 ( .A(n_304), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_339), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_343), .A2(n_296), .B(n_320), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_358), .A2(n_359), .B(n_323), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_350), .A2(n_307), .B1(n_292), .B2(n_253), .C(n_227), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_341), .A2(n_307), .B1(n_330), .B2(n_271), .C(n_263), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_337), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_327), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_361), .B(n_300), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_337), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_346), .A2(n_267), .B1(n_333), .B2(n_331), .C(n_300), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_357), .B1(n_338), .B2(n_306), .Y(n_374) );
OAI22xp33_ASAP7_75t_R g375 ( .A1(n_354), .A2(n_277), .B1(n_332), .B2(n_11), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_339), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_352), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g378 ( .A1(n_349), .A2(n_301), .B1(n_331), .B2(n_326), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_336), .A2(n_301), .B1(n_259), .B2(n_261), .C(n_272), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_334), .B(n_250), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_354), .B(n_299), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_353), .A2(n_303), .B1(n_232), .B2(n_294), .C(n_329), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_347), .A2(n_329), .B1(n_289), .B2(n_299), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_360), .A2(n_303), .B1(n_230), .B2(n_244), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_347), .A2(n_289), .B1(n_244), .B2(n_312), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_353), .A2(n_289), .B1(n_294), .B2(n_281), .Y(n_387) );
BUFx2_ASAP7_75t_SL g388 ( .A(n_347), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_348), .A2(n_289), .B1(n_284), .B2(n_281), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g390 ( .A1(n_362), .A2(n_316), .B1(n_247), .B2(n_257), .C(n_234), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_377), .B(n_352), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_377), .Y(n_393) );
AOI21x1_ASAP7_75t_L g394 ( .A1(n_365), .A2(n_320), .B(n_323), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_368), .B(n_146), .C(n_138), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_364), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_380), .A2(n_355), .B1(n_335), .B2(n_356), .C(n_247), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_375), .A2(n_340), .B1(n_289), .B2(n_351), .Y(n_398) );
OAI321xp33_ASAP7_75t_L g399 ( .A1(n_374), .A2(n_355), .A3(n_138), .B1(n_146), .B2(n_318), .C(n_257), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_382), .B(n_340), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_376), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_335), .B(n_356), .C(n_311), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_367), .A2(n_340), .B1(n_351), .B2(n_241), .C(n_255), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_381), .B(n_358), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_388), .Y(n_407) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_366), .A2(n_359), .B(n_311), .Y(n_408) );
NAND3xp33_ASAP7_75t_L g409 ( .A(n_383), .B(n_138), .C(n_146), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_379), .B(n_363), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_382), .A2(n_378), .B1(n_370), .B2(n_384), .C(n_375), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_369), .B(n_351), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_372), .B(n_363), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_369), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_371), .A2(n_241), .B(n_255), .C(n_274), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_372), .B(n_363), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_372), .B(n_241), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_388), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_387), .B(n_344), .C(n_324), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_385), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g424 ( .A1(n_385), .A2(n_363), .B1(n_312), .B2(n_304), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_390), .Y(n_425) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_421), .B(n_390), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_416), .B(n_389), .Y(n_427) );
NOR3xp33_ASAP7_75t_L g428 ( .A(n_411), .B(n_386), .C(n_344), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_411), .A2(n_318), .A3(n_313), .B(n_237), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g430 ( .A1(n_397), .A2(n_313), .B(n_248), .C(n_244), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_421), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_396), .B(n_8), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_396), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_401), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_393), .B(n_8), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_398), .A2(n_324), .B1(n_312), .B2(n_237), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_421), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_397), .A2(n_280), .B1(n_278), .B2(n_284), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_393), .B(n_10), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_401), .B(n_11), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_402), .B(n_12), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_416), .B(n_65), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
OAI211xp5_ASAP7_75t_L g448 ( .A1(n_407), .A2(n_255), .B(n_274), .C(n_278), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_391), .B(n_15), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_405), .B(n_16), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_405), .A2(n_278), .B1(n_280), .B2(n_248), .C(n_167), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_415), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_392), .B(n_17), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_392), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
INVx4_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_408), .Y(n_457) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_403), .B(n_178), .C(n_217), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_391), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_425), .A2(n_17), .A3(n_19), .B1(n_22), .B2(n_24), .B3(n_25), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_406), .B(n_27), .Y(n_462) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_403), .A2(n_248), .B(n_280), .C(n_322), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
BUFx3_ASAP7_75t_L g465 ( .A(n_410), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_408), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_420), .A2(n_324), .B1(n_325), .B2(n_293), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_420), .B(n_248), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_423), .B(n_31), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_400), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_408), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_420), .B(n_325), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_406), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_394), .Y(n_475) );
NAND4xp25_ASAP7_75t_L g476 ( .A(n_429), .B(n_404), .C(n_395), .D(n_400), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_471), .B(n_418), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_454), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_434), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_454), .B(n_425), .Y(n_480) );
NOR4xp25_ASAP7_75t_SL g481 ( .A(n_455), .B(n_399), .C(n_404), .D(n_395), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_460), .B(n_418), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_449), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_433), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_433), .B(n_414), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_455), .Y(n_486) );
AND4x1_ASAP7_75t_L g487 ( .A(n_430), .B(n_409), .C(n_422), .D(n_414), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_474), .B(n_413), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g489 ( .A1(n_430), .A2(n_428), .B(n_452), .Y(n_489) );
INVxp67_ASAP7_75t_L g490 ( .A(n_452), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_459), .B(n_419), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_459), .B(n_419), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_449), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_453), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_465), .A2(n_424), .B1(n_409), .B2(n_422), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_435), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_435), .B(n_424), .Y(n_498) );
BUFx2_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_436), .B(n_394), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_457), .B(n_32), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_437), .B(n_35), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_463), .B(n_399), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_437), .B(n_38), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_444), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_444), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_447), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_447), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_474), .B(n_39), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_465), .B(n_417), .Y(n_511) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_431), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_443), .B(n_417), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_464), .B(n_40), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_464), .B(n_41), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_466), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_456), .B(n_43), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_457), .B(n_44), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_475), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_443), .B(n_49), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_431), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_457), .B(n_55), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_440), .B(n_56), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_440), .B(n_57), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_466), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_440), .B(n_59), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_438), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_475), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_467), .Y(n_529) );
BUFx3_ASAP7_75t_L g530 ( .A(n_456), .Y(n_530) );
NAND2xp33_ASAP7_75t_R g531 ( .A(n_470), .B(n_64), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_467), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_530), .Y(n_533) );
AOI211xp5_ASAP7_75t_SL g534 ( .A1(n_489), .A2(n_463), .B(n_453), .C(n_432), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_483), .B(n_445), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_486), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_489), .A2(n_456), .B1(n_461), .B2(n_470), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_490), .B(n_472), .C(n_450), .Y(n_538) );
XOR2x2_ASAP7_75t_L g539 ( .A(n_493), .B(n_432), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_491), .B(n_445), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_491), .B(n_472), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_478), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_494), .B(n_438), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_480), .B(n_442), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_478), .Y(n_546) );
NAND2xp33_ASAP7_75t_SL g547 ( .A(n_531), .B(n_470), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_480), .B(n_442), .Y(n_548) );
OAI222xp33_ASAP7_75t_L g549 ( .A1(n_517), .A2(n_470), .B1(n_426), .B2(n_462), .C1(n_446), .C2(n_473), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_482), .A2(n_427), .B1(n_441), .B2(n_462), .C(n_458), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_484), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_477), .B(n_469), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_485), .B(n_427), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_485), .B(n_427), .Y(n_554) );
AOI21xp33_ASAP7_75t_L g555 ( .A1(n_511), .A2(n_426), .B(n_448), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_484), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_492), .B(n_427), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_497), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_530), .A2(n_446), .B(n_468), .C(n_473), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_501), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_497), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_496), .A2(n_446), .B1(n_451), .B2(n_439), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_499), .Y(n_563) );
NOR4xp25_ASAP7_75t_L g564 ( .A(n_476), .B(n_446), .C(n_67), .D(n_70), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_488), .B(n_66), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_504), .A2(n_73), .B(n_74), .C(n_274), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_517), .A2(n_274), .B(n_324), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_492), .B(n_248), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_527), .B(n_274), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_514), .A2(n_325), .B1(n_293), .B2(n_274), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_512), .B(n_178), .Y(n_571) );
OA21x2_ASAP7_75t_L g572 ( .A1(n_519), .A2(n_178), .B(n_185), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_498), .B(n_293), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_499), .A2(n_185), .B1(n_201), .B2(n_203), .Y(n_574) );
AOI211xp5_ASAP7_75t_L g575 ( .A1(n_476), .A2(n_185), .B(n_201), .C(n_203), .Y(n_575) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_498), .A2(n_201), .B(n_203), .C(n_217), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_500), .B(n_217), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_506), .B(n_265), .Y(n_579) );
XOR2x2_ASAP7_75t_L g580 ( .A(n_487), .B(n_265), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_507), .B(n_265), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g582 ( .A(n_487), .B(n_265), .C(n_270), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_533), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_542), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_546), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_534), .B(n_500), .C(n_521), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_551), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_536), .B(n_543), .Y(n_588) );
INVxp33_ASAP7_75t_L g589 ( .A(n_564), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_556), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_558), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_561), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_559), .A2(n_513), .B1(n_509), .B2(n_508), .C(n_520), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_555), .B(n_508), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_552), .Y(n_595) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_582), .B(n_515), .Y(n_596) );
OAI21xp33_ASAP7_75t_L g597 ( .A1(n_564), .A2(n_518), .B(n_522), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_540), .B(n_507), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_545), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_578), .B(n_509), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_560), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_563), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_553), .B(n_495), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_554), .B(n_516), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_549), .B(n_515), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_538), .B(n_510), .C(n_518), .Y(n_606) );
XNOR2xp5_ASAP7_75t_L g607 ( .A(n_539), .B(n_510), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_541), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_562), .B(n_514), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_535), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_557), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_544), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_548), .B(n_532), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_563), .B(n_495), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_569), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_547), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_573), .B(n_532), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_609), .A2(n_537), .B1(n_567), .B2(n_562), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_609), .A2(n_550), .B1(n_580), .B2(n_567), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_594), .B(n_534), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_589), .B(n_575), .C(n_576), .Y(n_621) );
OAI21xp5_ASAP7_75t_L g622 ( .A1(n_589), .A2(n_566), .B(n_570), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g623 ( .A1(n_616), .A2(n_570), .B1(n_565), .B2(n_502), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g624 ( .A(n_593), .B(n_481), .C(n_574), .Y(n_624) );
INVxp67_ASAP7_75t_L g625 ( .A(n_583), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_604), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_594), .B(n_571), .C(n_568), .Y(n_627) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_596), .B(n_502), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_604), .B(n_525), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_583), .B(n_577), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_595), .A2(n_516), .B1(n_525), .B2(n_529), .C(n_577), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_584), .Y(n_632) );
OA22x2_ASAP7_75t_L g633 ( .A1(n_607), .A2(n_502), .B1(n_526), .B2(n_524), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g634 ( .A(n_606), .B(n_523), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_615), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_585), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_597), .A2(n_522), .B(n_529), .C(n_502), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_590), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_618), .A2(n_605), .B(n_586), .C(n_610), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_633), .A2(n_605), .B(n_613), .Y(n_641) );
NAND3xp33_ASAP7_75t_SL g642 ( .A(n_622), .B(n_481), .C(n_602), .Y(n_642) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_633), .A2(n_602), .B(n_588), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_625), .Y(n_644) );
INVx4_ASAP7_75t_L g645 ( .A(n_630), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_618), .A2(n_612), .B1(n_608), .B2(n_611), .C(n_592), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_620), .B(n_591), .C(n_601), .Y(n_647) );
BUFx4f_ASAP7_75t_SL g648 ( .A(n_635), .Y(n_648) );
AOI222xp33_ASAP7_75t_L g649 ( .A1(n_634), .A2(n_603), .B1(n_614), .B2(n_600), .C1(n_599), .C2(n_505), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_637), .A2(n_598), .B1(n_599), .B2(n_617), .C(n_503), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g651 ( .A1(n_619), .A2(n_572), .B1(n_479), .B2(n_579), .Y(n_651) );
NOR2xp33_ASAP7_75t_R g652 ( .A(n_624), .B(n_523), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_621), .B(n_526), .C(n_524), .D(n_503), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_628), .A2(n_505), .B(n_479), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_631), .A2(n_572), .B(n_581), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_623), .A2(n_519), .B1(n_528), .B2(n_265), .Y(n_656) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_639), .A2(n_528), .B(n_270), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_627), .A2(n_270), .B1(n_626), .B2(n_632), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_638), .B(n_636), .C(n_629), .D(n_270), .Y(n_659) );
CKINVDCx12_ASAP7_75t_R g660 ( .A(n_648), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_644), .Y(n_661) );
AND2x4_ASAP7_75t_L g662 ( .A(n_645), .B(n_647), .Y(n_662) );
NAND4xp25_ASAP7_75t_L g663 ( .A(n_642), .B(n_640), .C(n_646), .D(n_641), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_658), .B1(n_659), .B2(n_645), .Y(n_664) );
OR4x1_ASAP7_75t_L g665 ( .A(n_660), .B(n_652), .C(n_643), .D(n_649), .Y(n_665) );
NAND4xp25_ASAP7_75t_SL g666 ( .A(n_662), .B(n_650), .C(n_656), .D(n_654), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_664), .B(n_661), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_665), .B(n_651), .Y(n_668) );
XNOR2xp5_ASAP7_75t_L g669 ( .A(n_667), .B(n_653), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_669), .A2(n_668), .B1(n_666), .B2(n_655), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_657), .B(n_270), .Y(n_671) );
endmodule