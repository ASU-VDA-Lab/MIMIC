module fake_jpeg_29121_n_424 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_424);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_424;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_378;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_62),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_18),
.B(n_9),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_18),
.B(n_16),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_81),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_19),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_67),
.A2(n_34),
.B(n_12),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_94),
.A2(n_111),
.B(n_107),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_52),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_107),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

CKINVDCx12_ASAP7_75t_R g159 ( 
.A(n_106),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_110),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_53),
.A2(n_41),
.B1(n_26),
.B2(n_39),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_121),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_40),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_36),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_39),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_45),
.A2(n_36),
.B1(n_24),
.B2(n_26),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_82),
.B1(n_47),
.B2(n_66),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_60),
.B(n_32),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_17),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_90),
.B(n_31),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_142),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_88),
.B(n_79),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_152),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_144),
.A2(n_165),
.B1(n_166),
.B2(n_120),
.Y(n_192)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_150),
.Y(n_191)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_17),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_23),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

BUFx2_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_61),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_167),
.C(n_96),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_69),
.B1(n_54),
.B2(n_24),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_168),
.B1(n_164),
.B2(n_157),
.Y(n_188)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_31),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_172),
.Y(n_175)
);

CKINVDCx9p33_ASAP7_75t_R g164 ( 
.A(n_85),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_SL g166 ( 
.A1(n_111),
.A2(n_30),
.B(n_65),
.C(n_63),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_90),
.A2(n_32),
.B(n_23),
.C(n_10),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_114),
.A2(n_24),
.B1(n_68),
.B2(n_15),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_99),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_121),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_167),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_134),
.B1(n_112),
.B2(n_119),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_190),
.B1(n_137),
.B2(n_86),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_158),
.B1(n_140),
.B2(n_109),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_134),
.B1(n_128),
.B2(n_97),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_125),
.B1(n_158),
.B2(n_108),
.Y(n_208)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_204),
.B1(n_214),
.B2(n_186),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_199),
.B(n_201),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_149),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_202),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_176),
.Y(n_201)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_87),
.B1(n_108),
.B2(n_115),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_89),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_187),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_89),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_156),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_148),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_10),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_217),
.Y(n_226)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_161),
.B1(n_169),
.B2(n_100),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_192),
.B1(n_193),
.B2(n_180),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_230),
.B1(n_231),
.B2(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_199),
.C(n_202),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_201),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_175),
.B1(n_193),
.B2(n_180),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_207),
.A2(n_132),
.B1(n_123),
.B2(n_181),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_207),
.A2(n_175),
.B(n_181),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_182),
.B1(n_185),
.B2(n_195),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_245),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_209),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_250),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_200),
.C(n_213),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_198),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_230),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_203),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_248),
.A2(n_227),
.B(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_249),
.Y(n_273)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_255),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_204),
.B1(n_217),
.B2(n_208),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_252),
.A2(n_231),
.B1(n_208),
.B2(n_235),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_258),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_218),
.B(n_212),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_218),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_197),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_217),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_221),
.C(n_229),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_223),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_226),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_215),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_268),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_233),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_226),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_251),
.B(n_233),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_274),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_238),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_238),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_225),
.B1(n_231),
.B2(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_279),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_242),
.B1(n_252),
.B2(n_255),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_245),
.C(n_247),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_203),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_267),
.B1(n_261),
.B2(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_292),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_298),
.B1(n_300),
.B2(n_265),
.Y(n_303)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_260),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_247),
.C(n_248),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_299),
.C(n_173),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_243),
.B1(n_249),
.B2(n_246),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_296),
.A2(n_210),
.B1(n_211),
.B2(n_206),
.Y(n_313)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_302),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_278),
.A2(n_243),
.B1(n_246),
.B2(n_232),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_221),
.C(n_220),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_259),
.A2(n_241),
.B1(n_229),
.B2(n_220),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_272),
.A2(n_250),
.B(n_219),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_303),
.A2(n_308),
.B1(n_143),
.B2(n_172),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_297),
.A2(n_281),
.B1(n_290),
.B2(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_305),
.B(n_307),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_273),
.B1(n_265),
.B2(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_275),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_273),
.B1(n_234),
.B2(n_206),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_293),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_316),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_315),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_211),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_182),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_323),
.C(n_326),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_285),
.B(n_184),
.Y(n_319)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_319),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_324),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_290),
.A2(n_203),
.B1(n_216),
.B2(n_196),
.Y(n_322)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_184),
.C(n_216),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_159),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_282),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_178),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_216),
.C(n_145),
.Y(n_326)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_345),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_292),
.B1(n_286),
.B2(n_283),
.Y(n_328)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_312),
.A2(n_286),
.B1(n_284),
.B2(n_280),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_332),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g332 ( 
.A(n_304),
.B(n_302),
.CI(n_280),
.CON(n_332),
.SN(n_332)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_178),
.C(n_195),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_336),
.B(n_344),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_307),
.B(n_11),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_341),
.B(n_10),
.Y(n_362)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_320),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_342),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_138),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_347),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_178),
.C(n_196),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_151),
.C(n_171),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_348),
.C(n_326),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_171),
.C(n_151),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_324),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_349),
.B(n_362),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g350 ( 
.A(n_345),
.B(n_314),
.Y(n_350)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_309),
.B(n_311),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_352),
.A2(n_363),
.B(n_343),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_357),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_308),
.B1(n_141),
.B2(n_153),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_359),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_174),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_170),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_348),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_340),
.B(n_162),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_174),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_339),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_332),
.A2(n_162),
.B(n_126),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_366),
.A2(n_346),
.B(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_333),
.C(n_336),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_376),
.C(n_378),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_377),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_361),
.A2(n_338),
.B1(n_327),
.B2(n_341),
.Y(n_374)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_375),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_339),
.C(n_133),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_122),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_103),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_379),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_103),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_135),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_372),
.A2(n_358),
.B1(n_363),
.B2(n_354),
.Y(n_383)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_383),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_368),
.A2(n_366),
.B1(n_350),
.B2(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_373),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_11),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_388),
.B(n_391),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_367),
.Y(n_391)
);

AOI21x1_ASAP7_75t_L g392 ( 
.A1(n_369),
.A2(n_15),
.B(n_14),
.Y(n_392)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_381),
.A2(n_390),
.B(n_385),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_393),
.A2(n_1),
.B(n_2),
.Y(n_406)
);

AOI31xp67_ASAP7_75t_SL g395 ( 
.A1(n_382),
.A2(n_371),
.A3(n_378),
.B(n_379),
.Y(n_395)
);

O2A1O1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_395),
.A2(n_92),
.B(n_129),
.C(n_130),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_396),
.B(n_129),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_388),
.A2(n_104),
.B1(n_131),
.B2(n_113),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_110),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_384),
.A2(n_387),
.B(n_124),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_401),
.A2(n_403),
.B(n_110),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_384),
.A2(n_170),
.B(n_24),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_397),
.A2(n_0),
.B(n_1),
.Y(n_404)
);

AOI322xp5_ASAP7_75t_L g412 ( 
.A1(n_404),
.A2(n_411),
.A3(n_398),
.B1(n_92),
.B2(n_24),
.C1(n_4),
.C2(n_5),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_407),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_406),
.A2(n_410),
.B(n_1),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_398),
.C(n_402),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_408),
.B(n_106),
.C(n_2),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_413),
.C(n_414),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_409),
.A2(n_1),
.B(n_2),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_3),
.C(n_5),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_416),
.A2(n_404),
.B(n_4),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_417),
.B(n_419),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_3),
.C(n_6),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_3),
.Y(n_422)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g423 ( 
.A1(n_422),
.A2(n_3),
.B(n_6),
.C(n_421),
.D(n_342),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_6),
.Y(n_424)
);


endmodule