module fake_ariane_2444_n_2817 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2817);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2817;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_762;
wire n_1661;
wire n_1468;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_727;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_2785;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1476;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_701;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1865;
wire n_1710;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_400),
.Y(n_617)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_188),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_40),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_560),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_442),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_242),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_219),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_350),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_539),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_304),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_149),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_26),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_316),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_375),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_159),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_128),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_553),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_558),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_491),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_311),
.Y(n_636)
);

BUFx8_ASAP7_75t_SL g637 ( 
.A(n_291),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_347),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_361),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_164),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_99),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_242),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_303),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_496),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_111),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_568),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_15),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_425),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_550),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_328),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_245),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_587),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_446),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_600),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_80),
.Y(n_655)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_344),
.Y(n_656)
);

CKINVDCx14_ASAP7_75t_R g657 ( 
.A(n_179),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_559),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_446),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_535),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_442),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_80),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_237),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_326),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_250),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_473),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_564),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_480),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_490),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_456),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_501),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_531),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_472),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_103),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_586),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_202),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_78),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_320),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_54),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_226),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_434),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_305),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_487),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_489),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_154),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_488),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_437),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_497),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_265),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_494),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_343),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_72),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_470),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_26),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_578),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_179),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_451),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_503),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_150),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_523),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_201),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_493),
.Y(n_702)
);

CKINVDCx16_ASAP7_75t_R g703 ( 
.A(n_540),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_87),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_430),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_367),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_85),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_407),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_200),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_437),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_77),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_119),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_236),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_188),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_334),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_224),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_163),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_500),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_52),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_114),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_107),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_485),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_581),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_122),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_201),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_433),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_264),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_309),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_137),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_251),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_391),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_70),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_228),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_566),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_176),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_497),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_206),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_346),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_178),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_555),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_44),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_527),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_495),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_231),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_185),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_362),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_5),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_342),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_291),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_164),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_283),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_462),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_226),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_534),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_87),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_507),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_454),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_574),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_152),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_466),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_45),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_104),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_362),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_491),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_71),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_452),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_414),
.Y(n_767)
);

CKINVDCx14_ASAP7_75t_R g768 ( 
.A(n_577),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_563),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_305),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_394),
.Y(n_771)
);

CKINVDCx16_ASAP7_75t_R g772 ( 
.A(n_222),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_402),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_247),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_258),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_509),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_273),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_588),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_116),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_573),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_160),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_112),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_392),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_457),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_440),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_239),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_27),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_256),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_0),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_160),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_348),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_522),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_392),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_474),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_375),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_204),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_57),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_289),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_37),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_369),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_606),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_562),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_500),
.Y(n_803)
);

BUFx10_ASAP7_75t_L g804 ( 
.A(n_607),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_333),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_447),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_157),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_360),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_611),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_57),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_517),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_91),
.Y(n_812)
);

INVxp33_ASAP7_75t_SL g813 ( 
.A(n_450),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_486),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_300),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_469),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_413),
.Y(n_817)
);

BUFx8_ASAP7_75t_SL g818 ( 
.A(n_315),
.Y(n_818)
);

BUFx10_ASAP7_75t_L g819 ( 
.A(n_546),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_398),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_23),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_371),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_315),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_46),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_241),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_410),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_97),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_373),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_526),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_9),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_287),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_245),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_379),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_135),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_390),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_12),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_428),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_290),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_389),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_499),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_161),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_463),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_111),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_45),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_529),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_33),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_359),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_181),
.Y(n_848)
);

BUFx10_ASAP7_75t_L g849 ( 
.A(n_86),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_281),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_477),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_5),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_37),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_322),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_294),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_492),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_286),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_484),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_209),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_498),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_308),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_221),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_185),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_3),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_166),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_443),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_386),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_659),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_657),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_659),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_710),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_668),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_668),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_711),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_711),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_712),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_710),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_710),
.Y(n_878)
);

INVxp33_ASAP7_75t_SL g879 ( 
.A(n_844),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_707),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_637),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_818),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_710),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_703),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_712),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_731),
.Y(n_886)
);

INVxp67_ASAP7_75t_SL g887 ( 
.A(n_713),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_731),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_731),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_731),
.Y(n_890)
);

INVxp33_ASAP7_75t_SL g891 ( 
.A(n_631),
.Y(n_891)
);

CKINVDCx16_ASAP7_75t_R g892 ( 
.A(n_618),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_753),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_713),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_753),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_734),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_778),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_753),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_753),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_810),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_810),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_810),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_829),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_810),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_828),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_734),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_812),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_718),
.Y(n_908)
);

INVxp33_ASAP7_75t_SL g909 ( 
.A(n_631),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_829),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_812),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_619),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_624),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_828),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_630),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_628),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_632),
.Y(n_917)
);

INVxp67_ASAP7_75t_SL g918 ( 
.A(n_828),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_828),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_674),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_638),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_674),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_639),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_644),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_645),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_648),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_693),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_663),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_669),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_620),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_620),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_670),
.Y(n_932)
);

INVxp33_ASAP7_75t_L g933 ( 
.A(n_817),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_620),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_693),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_658),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_706),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_706),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_656),
.Y(n_939)
);

BUFx10_ASAP7_75t_L g940 ( 
.A(n_633),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_721),
.Y(n_941)
);

INVxp33_ASAP7_75t_L g942 ( 
.A(n_679),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_721),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_766),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_766),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_660),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_787),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_787),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_662),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_789),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_667),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_630),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_772),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_789),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_723),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_796),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_804),
.Y(n_957)
);

INVxp33_ASAP7_75t_SL g958 ( 
.A(n_635),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_635),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_634),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_682),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_686),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_687),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_690),
.Y(n_964)
);

CKINVDCx14_ASAP7_75t_R g965 ( 
.A(n_768),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_742),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_754),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_769),
.Y(n_968)
);

BUFx5_ASAP7_75t_L g969 ( 
.A(n_845),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_960),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_960),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_871),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_918),
.B(n_633),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_881),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_960),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_960),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_871),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_960),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_883),
.Y(n_979)
);

BUFx12f_ASAP7_75t_L g980 ( 
.A(n_881),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_883),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_949),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_886),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_896),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_886),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_896),
.B(n_664),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_898),
.Y(n_987)
);

BUFx8_ASAP7_75t_SL g988 ( 
.A(n_915),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_930),
.B(n_776),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_874),
.B(n_885),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_898),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_901),
.Y(n_992)
);

BUFx8_ASAP7_75t_L g993 ( 
.A(n_939),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_906),
.B(n_664),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_901),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_914),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_887),
.B(n_634),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_914),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_877),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_877),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_878),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_878),
.Y(n_1002)
);

CKINVDCx16_ASAP7_75t_R g1003 ( 
.A(n_892),
.Y(n_1003)
);

CKINVDCx8_ASAP7_75t_R g1004 ( 
.A(n_882),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_888),
.Y(n_1005)
);

OA21x2_ASAP7_75t_L g1006 ( 
.A1(n_888),
.A2(n_890),
.B(n_889),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_939),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_889),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_936),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_890),
.Y(n_1010)
);

BUFx12f_ASAP7_75t_L g1011 ( 
.A(n_882),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_930),
.B(n_792),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_894),
.B(n_802),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_920),
.B(n_636),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_893),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_893),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_940),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_895),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_895),
.A2(n_802),
.B(n_796),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_899),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_952),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_959),
.Y(n_1022)
);

BUFx12f_ASAP7_75t_L g1023 ( 
.A(n_940),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_899),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_906),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_900),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_969),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_900),
.Y(n_1028)
);

OA21x2_ASAP7_75t_L g1029 ( 
.A1(n_902),
.A2(n_905),
.B(n_904),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_931),
.B(n_646),
.Y(n_1030)
);

AND2x6_ASAP7_75t_L g1031 ( 
.A(n_936),
.B(n_803),
.Y(n_1031)
);

OAI22x1_ASAP7_75t_L g1032 ( 
.A1(n_903),
.A2(n_647),
.B1(n_681),
.B2(n_640),
.Y(n_1032)
);

INVx5_ASAP7_75t_L g1033 ( 
.A(n_946),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_902),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_946),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1006),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1035),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_988),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_1017),
.B(n_940),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1035),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1006),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1035),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_1006),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_971),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1035),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1006),
.Y(n_1046)
);

AND2x6_ASAP7_75t_L g1047 ( 
.A(n_1014),
.B(n_1027),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1005),
.Y(n_1048)
);

CKINVDCx20_ASAP7_75t_R g1049 ( 
.A(n_1021),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_1023),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1005),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1008),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_989),
.A2(n_909),
.B1(n_958),
.B2(n_891),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1022),
.B(n_933),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_1004),
.B(n_965),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1008),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_R g1057 ( 
.A(n_1004),
.B(n_884),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_974),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1029),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1010),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_971),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_1007),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_R g1063 ( 
.A(n_1003),
.B(n_974),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1023),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_1023),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1017),
.B(n_957),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1029),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1010),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_1007),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_974),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_982),
.B(n_959),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1014),
.B(n_953),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_980),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1029),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_980),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_971),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_1003),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1016),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1012),
.B(n_884),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_984),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1016),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_984),
.B(n_955),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1020),
.Y(n_1083)
);

CKINVDCx11_ASAP7_75t_R g1084 ( 
.A(n_980),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1029),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1020),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_1011),
.Y(n_1087)
);

CKINVDCx6p67_ASAP7_75t_R g1088 ( 
.A(n_1011),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_R g1089 ( 
.A(n_986),
.B(n_903),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1028),
.Y(n_1090)
);

BUFx10_ASAP7_75t_L g1091 ( 
.A(n_1030),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_1011),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1028),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_993),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_993),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_993),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_990),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_999),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_993),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_984),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1025),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1025),
.B(n_973),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_999),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_986),
.B(n_897),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1025),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_999),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_997),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_1013),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_970),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_986),
.B(n_967),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_1009),
.B(n_957),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_970),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_973),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_986),
.B(n_897),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_994),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1019),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1032),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_1019),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_994),
.B(n_934),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_978),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_978),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_994),
.Y(n_1122)
);

XNOR2xp5_ASAP7_75t_L g1123 ( 
.A(n_1032),
.B(n_910),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_994),
.B(n_931),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1019),
.Y(n_1125)
);

AND2x2_ASAP7_75t_SL g1126 ( 
.A(n_1094),
.B(n_1095),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1100),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1097),
.B(n_934),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1048),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_L g1130 ( 
.A(n_1062),
.B(n_910),
.C(n_749),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1101),
.B(n_1027),
.Y(n_1131)
);

NAND2xp33_ASAP7_75t_L g1132 ( 
.A(n_1047),
.B(n_969),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1044),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1047),
.B(n_891),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_1050),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1054),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1051),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1101),
.B(n_1027),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1098),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_1125),
.B(n_1036),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1047),
.A2(n_879),
.B1(n_958),
.B2(n_909),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1098),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1119),
.B(n_813),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1052),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1049),
.Y(n_1145)
);

AND2x6_ASAP7_75t_L g1146 ( 
.A(n_1036),
.B(n_803),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1103),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1091),
.B(n_969),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1103),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1056),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1102),
.B(n_813),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1060),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1106),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1106),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1047),
.B(n_955),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1041),
.Y(n_1156)
);

OAI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1053),
.A2(n_717),
.B1(n_764),
.B2(n_738),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1041),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1077),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1047),
.B(n_1110),
.Y(n_1160)
);

NOR3xp33_ASAP7_75t_L g1161 ( 
.A(n_1079),
.B(n_825),
.C(n_701),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1038),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1046),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1046),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1068),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1110),
.B(n_951),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1078),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1044),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1038),
.Y(n_1169)
);

AND2x6_ASAP7_75t_L g1170 ( 
.A(n_1059),
.B(n_814),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1071),
.B(n_880),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1081),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1083),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1072),
.B(n_908),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1091),
.B(n_969),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1047),
.B(n_967),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1069),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1086),
.Y(n_1178)
);

INVx5_ASAP7_75t_L g1179 ( 
.A(n_1044),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1084),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1090),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_SL g1182 ( 
.A(n_1057),
.B(n_764),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1049),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1110),
.B(n_969),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1070),
.B(n_869),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1091),
.B(n_969),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_1044),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1059),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1067),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1104),
.B(n_942),
.Y(n_1190)
);

INVxp33_ASAP7_75t_SL g1191 ( 
.A(n_1063),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1111),
.B(n_1113),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1067),
.Y(n_1193)
);

NOR2x1p5_ASAP7_75t_L g1194 ( 
.A(n_1088),
.B(n_641),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1080),
.B(n_879),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1074),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1061),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1100),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1113),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1074),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1055),
.B(n_922),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_1088),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1093),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1085),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1089),
.Y(n_1205)
);

INVxp33_ASAP7_75t_SL g1206 ( 
.A(n_1070),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1082),
.Y(n_1207)
);

INVxp33_ASAP7_75t_L g1208 ( 
.A(n_1114),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1085),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1037),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1082),
.B(n_969),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1061),
.B(n_969),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1124),
.B(n_689),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_1050),
.Y(n_1214)
);

CKINVDCx6p67_ASAP7_75t_R g1215 ( 
.A(n_1084),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1043),
.A2(n_1019),
.B(n_1031),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1073),
.Y(n_1217)
);

AND2x2_ASAP7_75t_SL g1218 ( 
.A(n_1082),
.B(n_814),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1040),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1107),
.B(n_937),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1042),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1115),
.B(n_951),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1043),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1116),
.A2(n_717),
.B1(n_765),
.B2(n_738),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1116),
.A2(n_765),
.B1(n_791),
.B2(n_771),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1043),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1061),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1045),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1109),
.Y(n_1229)
);

AND2x6_ASAP7_75t_L g1230 ( 
.A(n_1105),
.B(n_820),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1122),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1112),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1120),
.Y(n_1233)
);

BUFx4f_ASAP7_75t_L g1234 ( 
.A(n_1121),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1061),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1118),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1076),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1118),
.A2(n_1031),
.B1(n_791),
.B2(n_800),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1073),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1076),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1076),
.Y(n_1241)
);

AO22x2_ASAP7_75t_L g1242 ( 
.A1(n_1117),
.A2(n_683),
.B1(n_862),
.B2(n_807),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1076),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1075),
.B(n_1087),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1107),
.B(n_966),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1108),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1064),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1108),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1039),
.Y(n_1249)
);

AOI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1066),
.A2(n_996),
.B(n_1015),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1064),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1117),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1123),
.A2(n_968),
.B(n_966),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1096),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1096),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1099),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1065),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1065),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1099),
.Y(n_1259)
);

INVx5_ASAP7_75t_L g1260 ( 
.A(n_1058),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1075),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1087),
.B(n_646),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1092),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1092),
.B(n_968),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1208),
.B(n_649),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1208),
.B(n_649),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1151),
.B(n_941),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1129),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1171),
.B(n_944),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1133),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1151),
.B(n_683),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1127),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1195),
.B(n_800),
.C(n_771),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1128),
.B(n_808),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1218),
.B(n_652),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1218),
.B(n_652),
.Y(n_1276)
);

NAND2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1258),
.B(n_808),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1137),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1143),
.B(n_830),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1166),
.B(n_1009),
.Y(n_1280)
);

NAND3xp33_ASAP7_75t_SL g1281 ( 
.A(n_1161),
.B(n_830),
.C(n_642),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1195),
.B(n_642),
.C(n_641),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1139),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1166),
.B(n_1009),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1166),
.B(n_1009),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1144),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1190),
.B(n_1009),
.Y(n_1287)
);

NAND2x1_ASAP7_75t_L g1288 ( 
.A(n_1187),
.B(n_971),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1143),
.B(n_643),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1234),
.A2(n_696),
.B(n_697),
.C(n_691),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_1260),
.B(n_868),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1187),
.Y(n_1292)
);

AOI221xp5_ASAP7_75t_L g1293 ( 
.A1(n_1157),
.A2(n_916),
.B1(n_917),
.B2(n_913),
.C(n_912),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1142),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1142),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1174),
.B(n_870),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1205),
.B(n_643),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1220),
.B(n_872),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1264),
.B(n_1009),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1160),
.B(n_654),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_L g1301 ( 
.A(n_1264),
.B(n_709),
.C(n_699),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1134),
.B(n_654),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1234),
.B(n_971),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_L g1304 ( 
.A(n_1148),
.B(n_650),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1147),
.Y(n_1305)
);

BUFx5_ASAP7_75t_L g1306 ( 
.A(n_1140),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1201),
.B(n_1033),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1177),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1150),
.B(n_1033),
.Y(n_1309)
);

NOR2xp67_ASAP7_75t_L g1310 ( 
.A(n_1260),
.B(n_873),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1207),
.B(n_650),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1147),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1152),
.B(n_1033),
.Y(n_1313)
);

NAND2xp33_ASAP7_75t_L g1314 ( 
.A(n_1148),
.B(n_651),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1165),
.B(n_1033),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1149),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1167),
.B(n_1033),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1207),
.B(n_651),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1207),
.B(n_653),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1172),
.B(n_1033),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1173),
.B(n_1031),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1178),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1260),
.B(n_653),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1181),
.B(n_1031),
.Y(n_1324)
);

NAND2xp33_ASAP7_75t_L g1325 ( 
.A(n_1175),
.B(n_842),
.Y(n_1325)
);

AO221x1_ASAP7_75t_L g1326 ( 
.A1(n_1242),
.A2(n_714),
.B1(n_726),
.B2(n_722),
.C(n_716),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1149),
.Y(n_1327)
);

BUFx8_ASAP7_75t_L g1328 ( 
.A(n_1217),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1203),
.B(n_1031),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1141),
.A2(n_1031),
.B1(n_621),
.B2(n_622),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1184),
.B(n_971),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1153),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1222),
.B(n_1031),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1245),
.B(n_1031),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1231),
.B(n_842),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1136),
.B(n_875),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1153),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1229),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1213),
.B(n_846),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1213),
.B(n_846),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1260),
.B(n_1261),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1154),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1154),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1229),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1156),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1232),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1156),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1261),
.B(n_847),
.Y(n_1348)
);

BUFx2_ASAP7_75t_R g1349 ( 
.A(n_1180),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1233),
.B(n_847),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1159),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1158),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1210),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1162),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1249),
.B(n_1155),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1249),
.B(n_850),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1199),
.Y(n_1357)
);

NOR3xp33_ASAP7_75t_L g1358 ( 
.A(n_1130),
.B(n_741),
.C(n_733),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1158),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1261),
.B(n_850),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1219),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1127),
.Y(n_1362)
);

NOR3xp33_ASAP7_75t_L g1363 ( 
.A(n_1262),
.B(n_750),
.C(n_744),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1126),
.B(n_876),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1145),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1192),
.B(n_853),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1126),
.B(n_907),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1132),
.A2(n_755),
.B(n_757),
.C(n_751),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1224),
.B(n_855),
.C(n_853),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1163),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1221),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1176),
.B(n_855),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1223),
.B(n_856),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1258),
.B(n_856),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1163),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1132),
.A2(n_763),
.B(n_770),
.C(n_760),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1192),
.B(n_858),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1223),
.B(n_858),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1246),
.B(n_911),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1183),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1226),
.B(n_1164),
.Y(n_1381)
);

NAND2xp33_ASAP7_75t_L g1382 ( 
.A(n_1175),
.B(n_860),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1164),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1258),
.B(n_1247),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1238),
.B(n_1262),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1259),
.B(n_860),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1228),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1188),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1259),
.B(n_863),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1188),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1244),
.B(n_921),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1247),
.B(n_863),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1189),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1248),
.B(n_1225),
.Y(n_1394)
);

NOR2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1215),
.B(n_864),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1189),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1211),
.A2(n_779),
.B(n_782),
.C(n_774),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_SL g1398 ( 
.A(n_1135),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1198),
.B(n_923),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1193),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1193),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1236),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1226),
.B(n_975),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1196),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1162),
.B(n_865),
.C(n_864),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1196),
.B(n_865),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1200),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1239),
.B(n_924),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_SL g1409 ( 
.A(n_1135),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1200),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1169),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1204),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1204),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1209),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1209),
.Y(n_1415)
);

NAND2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1247),
.B(n_866),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1250),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1133),
.B(n_975),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1257),
.B(n_925),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1202),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1140),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1140),
.Y(n_1422)
);

NAND3xp33_ASAP7_75t_L g1423 ( 
.A(n_1169),
.B(n_866),
.C(n_671),
.Y(n_1423)
);

NOR3xp33_ASAP7_75t_L g1424 ( 
.A(n_1251),
.B(n_797),
.C(n_794),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1251),
.B(n_617),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1253),
.B(n_820),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1237),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1140),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1253),
.B(n_836),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1251),
.B(n_623),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1237),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1240),
.Y(n_1432)
);

CKINVDCx16_ASAP7_75t_R g1433 ( 
.A(n_1185),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1140),
.Y(n_1434)
);

INVxp33_ASAP7_75t_L g1435 ( 
.A(n_1185),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1206),
.B(n_626),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1254),
.B(n_627),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1133),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1187),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1255),
.B(n_629),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1230),
.B(n_836),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1133),
.B(n_1186),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1257),
.B(n_661),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1240),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1241),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1146),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1179),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1191),
.B(n_665),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1230),
.B(n_843),
.Y(n_1449)
);

NOR3xp33_ASAP7_75t_L g1450 ( 
.A(n_1263),
.B(n_824),
.C(n_805),
.Y(n_1450)
);

NOR3xp33_ASAP7_75t_L g1451 ( 
.A(n_1182),
.B(n_837),
.C(n_832),
.Y(n_1451)
);

BUFx5_ASAP7_75t_L g1452 ( 
.A(n_1146),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1186),
.B(n_975),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1256),
.B(n_666),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1241),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1191),
.B(n_1135),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1182),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1252),
.B(n_673),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1252),
.B(n_676),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1214),
.B(n_677),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1230),
.B(n_1170),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1279),
.B(n_1214),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1268),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1278),
.Y(n_1464)
);

AO22x2_ASAP7_75t_L g1465 ( 
.A1(n_1273),
.A2(n_1242),
.B1(n_1138),
.B2(n_1131),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1354),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1393),
.Y(n_1467)
);

AO22x2_ASAP7_75t_L g1468 ( 
.A1(n_1301),
.A2(n_1242),
.B1(n_1138),
.B2(n_1131),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1362),
.B(n_1194),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1420),
.B(n_1179),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1279),
.A2(n_1214),
.B1(n_1202),
.B2(n_1180),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1400),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1433),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1269),
.B(n_1215),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1404),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1283),
.Y(n_1476)
);

AO22x2_ASAP7_75t_L g1477 ( 
.A1(n_1301),
.A2(n_1216),
.B1(n_935),
.B2(n_938),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1286),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1322),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1420),
.B(n_1179),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1274),
.B(n_1243),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1346),
.Y(n_1482)
);

BUFx8_ASAP7_75t_L g1483 ( 
.A(n_1398),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1328),
.Y(n_1484)
);

NAND2xp33_ASAP7_75t_L g1485 ( 
.A(n_1447),
.B(n_1230),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1294),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1289),
.A2(n_1170),
.B1(n_1227),
.B2(n_680),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1353),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1411),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1295),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1289),
.A2(n_1170),
.B1(n_1227),
.B2(n_684),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1361),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1305),
.Y(n_1493)
);

NAND2x1p5_ASAP7_75t_L g1494 ( 
.A(n_1365),
.B(n_1227),
.Y(n_1494)
);

AO22x2_ASAP7_75t_L g1495 ( 
.A1(n_1369),
.A2(n_935),
.B1(n_938),
.B2(n_927),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1312),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1308),
.B(n_1168),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1385),
.A2(n_1274),
.B1(n_1277),
.B2(n_1436),
.Y(n_1498)
);

NAND2x1p5_ASAP7_75t_L g1499 ( 
.A(n_1272),
.B(n_1168),
.Y(n_1499)
);

OAI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1358),
.A2(n_929),
.B1(n_932),
.B2(n_928),
.C(n_926),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1380),
.B(n_1168),
.Y(n_1501)
);

NAND2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1357),
.B(n_1197),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1267),
.B(n_1170),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1371),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1316),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1451),
.A2(n_943),
.B1(n_945),
.B2(n_927),
.Y(n_1506)
);

AO22x2_ASAP7_75t_L g1507 ( 
.A1(n_1451),
.A2(n_945),
.B1(n_947),
.B2(n_943),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1387),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1457),
.B(n_1456),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1338),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1447),
.B(n_1197),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1385),
.A2(n_1170),
.B1(n_685),
.B2(n_688),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1328),
.Y(n_1513)
);

AO22x2_ASAP7_75t_L g1514 ( 
.A1(n_1394),
.A2(n_948),
.B1(n_950),
.B2(n_947),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1395),
.B(n_961),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1327),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1344),
.Y(n_1517)
);

OAI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1358),
.A2(n_964),
.B1(n_963),
.B2(n_962),
.C(n_851),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1424),
.A2(n_1235),
.B(n_1197),
.C(n_1212),
.Y(n_1519)
);

AO22x2_ASAP7_75t_L g1520 ( 
.A1(n_1281),
.A2(n_950),
.B1(n_954),
.B2(n_948),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1402),
.B(n_1235),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1447),
.B(n_1235),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1271),
.A2(n_1212),
.B1(n_692),
.B2(n_694),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1332),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1399),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1419),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1436),
.A2(n_852),
.B1(n_854),
.B2(n_848),
.C(n_840),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1337),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1342),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1402),
.B(n_954),
.Y(n_1530)
);

BUFx8_ASAP7_75t_L g1531 ( 
.A(n_1398),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1343),
.Y(n_1532)
);

AO22x2_ASAP7_75t_L g1533 ( 
.A1(n_1281),
.A2(n_956),
.B1(n_859),
.B2(n_861),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1364),
.B(n_636),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1336),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1415),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1345),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1347),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1308),
.Y(n_1539)
);

AO22x2_ASAP7_75t_L g1540 ( 
.A1(n_1363),
.A2(n_956),
.B1(n_857),
.B2(n_996),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1447),
.B(n_985),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1352),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1367),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1292),
.Y(n_1544)
);

AO22x2_ASAP7_75t_L g1545 ( 
.A1(n_1363),
.A2(n_1018),
.B1(n_1024),
.B2(n_1015),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1359),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1391),
.B(n_985),
.Y(n_1547)
);

AND2x6_ASAP7_75t_L g1548 ( 
.A(n_1421),
.B(n_1015),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1370),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1375),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1296),
.B(n_636),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1383),
.Y(n_1552)
);

AO22x2_ASAP7_75t_L g1553 ( 
.A1(n_1426),
.A2(n_1024),
.B1(n_1026),
.B2(n_1018),
.Y(n_1553)
);

AO22x2_ASAP7_75t_L g1554 ( 
.A1(n_1429),
.A2(n_1024),
.B1(n_1026),
.B2(n_1018),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1388),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1390),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1396),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1298),
.B(n_678),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1401),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1292),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1339),
.B(n_702),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1340),
.B(n_704),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1407),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1410),
.Y(n_1564)
);

OAI221xp5_ASAP7_75t_L g1565 ( 
.A1(n_1450),
.A2(n_708),
.B1(n_719),
.B2(n_715),
.C(n_705),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1351),
.B(n_985),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1326),
.A2(n_655),
.B1(n_745),
.B2(n_724),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1412),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1413),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1351),
.B(n_720),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1414),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1408),
.B(n_1379),
.Y(n_1572)
);

NOR2xp67_ASAP7_75t_L g1573 ( 
.A(n_1380),
.B(n_985),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1435),
.B(n_725),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1349),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1297),
.B(n_727),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1297),
.B(n_728),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1458),
.A2(n_655),
.B1(n_745),
.B2(n_724),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1427),
.Y(n_1579)
);

AO22x2_ASAP7_75t_L g1580 ( 
.A1(n_1450),
.A2(n_1026),
.B1(n_724),
.B2(n_745),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1431),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1432),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1444),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1424),
.A2(n_730),
.B1(n_735),
.B2(n_732),
.C(n_729),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1445),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1270),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1430),
.B(n_736),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1455),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1381),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1458),
.A2(n_739),
.B1(n_747),
.B2(n_743),
.C(n_737),
.Y(n_1590)
);

AND2x2_ASAP7_75t_SL g1591 ( 
.A(n_1366),
.B(n_804),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1406),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1373),
.Y(n_1593)
);

AO22x2_ASAP7_75t_L g1594 ( 
.A1(n_1275),
.A2(n_849),
.B1(n_655),
.B2(n_972),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1417),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1311),
.B(n_849),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1439),
.B(n_979),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1291),
.B(n_1310),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1311),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1459),
.A2(n_752),
.B1(n_759),
.B2(n_748),
.C(n_746),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1318),
.B(n_849),
.Y(n_1601)
);

NAND2x1p5_ASAP7_75t_L g1602 ( 
.A(n_1439),
.B(n_979),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1409),
.Y(n_1603)
);

OAI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1459),
.A2(n_773),
.B1(n_775),
.B2(n_762),
.C(n_761),
.Y(n_1604)
);

AO22x2_ASAP7_75t_L g1605 ( 
.A1(n_1276),
.A2(n_977),
.B1(n_983),
.B2(n_972),
.Y(n_1605)
);

OAI221xp5_ASAP7_75t_L g1606 ( 
.A1(n_1386),
.A2(n_781),
.B1(n_783),
.B2(n_777),
.C(n_767),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1430),
.B(n_784),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1378),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1350),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1403),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1441),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1443),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1449),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1446),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1321),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1282),
.B(n_1318),
.Y(n_1616)
);

NAND2x1p5_ASAP7_75t_L g1617 ( 
.A(n_1270),
.B(n_979),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1416),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1324),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1319),
.A2(n_786),
.B1(n_788),
.B2(n_785),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1386),
.B(n_790),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1389),
.B(n_793),
.Y(n_1622)
);

NAND2x1p5_ASAP7_75t_L g1623 ( 
.A(n_1270),
.B(n_979),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1329),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1389),
.B(n_795),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1319),
.B(n_798),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1355),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1422),
.Y(n_1628)
);

AO22x2_ASAP7_75t_L g1629 ( 
.A1(n_1428),
.A2(n_977),
.B1(n_983),
.B2(n_972),
.Y(n_1629)
);

AO22x2_ASAP7_75t_L g1630 ( 
.A1(n_1434),
.A2(n_983),
.B1(n_987),
.B2(n_977),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1384),
.B(n_987),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1356),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1437),
.A2(n_815),
.B1(n_816),
.B2(n_806),
.C(n_799),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1397),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1437),
.B(n_821),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1334),
.Y(n_1636)
);

NAND2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1270),
.B(n_979),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1440),
.A2(n_823),
.B1(n_826),
.B2(n_822),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1335),
.Y(n_1639)
);

NAND2x1p5_ASAP7_75t_L g1640 ( 
.A(n_1438),
.B(n_979),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1290),
.Y(n_1641)
);

AND2x6_ASAP7_75t_L g1642 ( 
.A(n_1438),
.B(n_987),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_SL g1643 ( 
.A(n_1409),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1438),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1366),
.B(n_827),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1440),
.A2(n_833),
.B1(n_834),
.B2(n_831),
.Y(n_1646)
);

AO22x2_ASAP7_75t_L g1647 ( 
.A1(n_1302),
.A2(n_998),
.B1(n_991),
.B2(n_904),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1377),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1372),
.A2(n_838),
.B1(n_839),
.B2(n_835),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1287),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1309),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1438),
.B(n_981),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1377),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1280),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1313),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1448),
.Y(n_1656)
);

NOR2xp67_ASAP7_75t_L g1657 ( 
.A(n_1423),
.B(n_1405),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1341),
.B(n_991),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1315),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1306),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1317),
.Y(n_1661)
);

OAI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1454),
.A2(n_867),
.B1(n_841),
.B2(n_919),
.C(n_905),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1454),
.B(n_819),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1284),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1660),
.A2(n_1299),
.B(n_1442),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1663),
.A2(n_1376),
.B(n_1368),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1498),
.A2(n_1330),
.B1(n_1266),
.B2(n_1265),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1485),
.A2(n_1442),
.B(n_1453),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1572),
.B(n_1293),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1526),
.B(n_1374),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1576),
.A2(n_1302),
.B(n_1453),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1519),
.A2(n_1331),
.B(n_1303),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1651),
.A2(n_1331),
.B(n_1303),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1577),
.A2(n_1300),
.B(n_1304),
.Y(n_1674)
);

O2A1O1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1616),
.A2(n_1348),
.B(n_1392),
.C(n_1360),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1481),
.A2(n_1325),
.B(n_1382),
.C(n_1314),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1655),
.A2(n_1418),
.B(n_1461),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1599),
.B(n_1460),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1659),
.A2(n_1418),
.B(n_1288),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1661),
.A2(n_1300),
.B(n_1425),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1636),
.A2(n_1320),
.B(n_1333),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1653),
.B(n_1323),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1525),
.B(n_1307),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1587),
.A2(n_1285),
.B1(n_1306),
.B2(n_672),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1648),
.B(n_1591),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1534),
.B(n_1543),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1535),
.B(n_1306),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1503),
.A2(n_1306),
.B(n_1452),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1551),
.B(n_819),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_R g1690 ( 
.A(n_1466),
.B(n_1306),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1607),
.A2(n_1306),
.B(n_1452),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1462),
.B(n_1452),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1539),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1621),
.A2(n_998),
.B(n_2),
.C(n_0),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1615),
.A2(n_1619),
.B(n_1624),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1474),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1615),
.A2(n_1452),
.B(n_976),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1622),
.A2(n_675),
.B1(n_695),
.B2(n_625),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1521),
.B(n_1509),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1619),
.A2(n_1452),
.B(n_976),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1626),
.B(n_819),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1468),
.A2(n_1465),
.B1(n_1514),
.B2(n_1533),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1650),
.A2(n_976),
.B(n_975),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1586),
.A2(n_1635),
.B(n_1610),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1544),
.A2(n_976),
.B(n_700),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1463),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1521),
.B(n_981),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1544),
.A2(n_976),
.B(n_740),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1645),
.B(n_1001),
.C(n_1000),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1560),
.A2(n_756),
.B(n_698),
.Y(n_1710)
);

O2A1O1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1625),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1641),
.A2(n_1001),
.B(n_1002),
.C(n_1000),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1561),
.A2(n_780),
.B(n_758),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1464),
.Y(n_1714)
);

O2A1O1Ixp33_ASAP7_75t_L g1715 ( 
.A1(n_1527),
.A2(n_6),
.B(n_1),
.C(n_4),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1476),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1468),
.A2(n_1001),
.B1(n_1002),
.B2(n_1000),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1562),
.A2(n_809),
.B(n_801),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1596),
.B(n_1601),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1609),
.A2(n_811),
.B(n_4),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1489),
.B(n_6),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1471),
.A2(n_1001),
.B1(n_1002),
.B2(n_1000),
.Y(n_1722)
);

AO32x1_ASAP7_75t_L g1723 ( 
.A1(n_1595),
.A2(n_995),
.A3(n_992),
.B1(n_981),
.B2(n_9),
.Y(n_1723)
);

AO32x2_ASAP7_75t_L g1724 ( 
.A1(n_1523),
.A2(n_995),
.A3(n_992),
.B1(n_981),
.B2(n_1000),
.Y(n_1724)
);

BUFx4f_ASAP7_75t_L g1725 ( 
.A(n_1515),
.Y(n_1725)
);

BUFx4f_ASAP7_75t_L g1726 ( 
.A(n_1515),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1639),
.B(n_1530),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1483),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1560),
.A2(n_1001),
.B(n_1000),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1530),
.B(n_1001),
.Y(n_1730)
);

AOI21xp33_ASAP7_75t_L g1731 ( 
.A1(n_1662),
.A2(n_992),
.B(n_981),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1597),
.A2(n_1034),
.B(n_1002),
.Y(n_1732)
);

A2O1A1Ixp33_ASAP7_75t_L g1733 ( 
.A1(n_1512),
.A2(n_1034),
.B(n_1002),
.C(n_992),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1602),
.A2(n_1034),
.B(n_1002),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1477),
.A2(n_1034),
.B(n_992),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1509),
.B(n_1501),
.Y(n_1736)
);

BUFx4f_ASAP7_75t_L g1737 ( 
.A(n_1469),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1486),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1490),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1533),
.B(n_7),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1632),
.A2(n_1608),
.B(n_1593),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1477),
.A2(n_1034),
.B(n_992),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1627),
.A2(n_1491),
.B(n_1487),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_SL g1744 ( 
.A(n_1575),
.B(n_981),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1618),
.B(n_7),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1638),
.A2(n_1034),
.B1(n_995),
.B2(n_11),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1627),
.A2(n_995),
.B(n_504),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1473),
.A2(n_995),
.B1(n_11),
.B2(n_8),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1612),
.B(n_995),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1497),
.A2(n_505),
.B(n_502),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1592),
.A2(n_508),
.B(n_506),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1558),
.B(n_8),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1649),
.A2(n_10),
.B(n_12),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1617),
.A2(n_1637),
.B(n_1623),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1478),
.B(n_10),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_L g1756 ( 
.A(n_1484),
.B(n_510),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1470),
.Y(n_1757)
);

AOI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1553),
.A2(n_512),
.B(n_511),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1479),
.B(n_13),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1640),
.A2(n_1652),
.B(n_1628),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1482),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1488),
.B(n_13),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1492),
.B(n_14),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1566),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1480),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1628),
.A2(n_514),
.B(n_513),
.Y(n_1766)
);

AO22x1_ASAP7_75t_L g1767 ( 
.A1(n_1483),
.A2(n_1531),
.B1(n_1513),
.B2(n_1603),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_SL g1768 ( 
.A(n_1643),
.B(n_515),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1634),
.A2(n_16),
.B(n_17),
.C(n_15),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1598),
.B(n_516),
.Y(n_1770)
);

NAND2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1598),
.B(n_518),
.Y(n_1771)
);

O2A1O1Ixp33_ASAP7_75t_SL g1772 ( 
.A1(n_1570),
.A2(n_17),
.B(n_14),
.C(n_16),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1631),
.A2(n_1554),
.B(n_1589),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1631),
.A2(n_520),
.B(n_519),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1646),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1578),
.B(n_18),
.C(n_19),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1554),
.A2(n_524),
.B(n_521),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1642),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1493),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1504),
.B(n_20),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1584),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1511),
.A2(n_528),
.B(n_525),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1574),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1522),
.A2(n_1605),
.B(n_1644),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1508),
.B(n_21),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1496),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1520),
.B(n_22),
.Y(n_1787)
);

AOI21x1_ASAP7_75t_L g1788 ( 
.A1(n_1605),
.A2(n_532),
.B(n_530),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1510),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1620),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1514),
.B(n_24),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1502),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1465),
.B(n_25),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1467),
.A2(n_536),
.B(n_533),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1565),
.B(n_28),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1467),
.A2(n_538),
.B(n_537),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1517),
.Y(n_1797)
);

BUFx2_ASAP7_75t_L g1798 ( 
.A(n_1566),
.Y(n_1798)
);

OAI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1590),
.A2(n_1600),
.B1(n_1604),
.B2(n_1606),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1472),
.A2(n_542),
.B(n_541),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1494),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1642),
.Y(n_1802)
);

O2A1O1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1633),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1642),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1642),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1531),
.Y(n_1806)
);

O2A1O1Ixp5_ASAP7_75t_L g1807 ( 
.A1(n_1658),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1520),
.B(n_31),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1499),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1505),
.Y(n_1810)
);

A2O1A1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1657),
.A2(n_34),
.B(n_35),
.C(n_33),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1472),
.A2(n_544),
.B(n_543),
.Y(n_1812)
);

O2A1O1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1656),
.A2(n_35),
.B(n_32),
.C(n_34),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1475),
.A2(n_547),
.B(n_545),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1573),
.B(n_32),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1547),
.Y(n_1816)
);

OA22x2_ASAP7_75t_L g1817 ( 
.A1(n_1654),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1547),
.A2(n_1664),
.B(n_1611),
.C(n_1613),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1541),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1580),
.B(n_36),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1475),
.A2(n_549),
.B(n_548),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1540),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1536),
.B(n_41),
.Y(n_1823)
);

O2A1O1Ixp33_ASAP7_75t_L g1824 ( 
.A1(n_1518),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1516),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1658),
.Y(n_1826)
);

AOI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1594),
.A2(n_42),
.B(n_43),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1567),
.A2(n_47),
.B(n_44),
.C(n_46),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1647),
.A2(n_552),
.B(n_551),
.Y(n_1829)
);

INVx1_ASAP7_75t_SL g1830 ( 
.A(n_1579),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1647),
.A2(n_556),
.B(n_554),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1580),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1614),
.A2(n_561),
.B(n_557),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1643),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1540),
.B(n_48),
.Y(n_1835)
);

NAND2x1p5_ASAP7_75t_L g1836 ( 
.A(n_1581),
.B(n_565),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1500),
.B(n_49),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1594),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1838)
);

INVx11_ASAP7_75t_L g1839 ( 
.A(n_1548),
.Y(n_1839)
);

BUFx6f_ASAP7_75t_L g1840 ( 
.A(n_1548),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1506),
.B(n_50),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1506),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_L g1843 ( 
.A(n_1582),
.B(n_53),
.C(n_55),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1507),
.B(n_55),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1507),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1524),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1528),
.B(n_56),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1529),
.B(n_58),
.Y(n_1848)
);

A2O1A1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1583),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_1849)
);

AOI33xp33_ASAP7_75t_L g1850 ( 
.A1(n_1585),
.A2(n_62),
.A3(n_64),
.B1(n_60),
.B2(n_61),
.B3(n_63),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1588),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1548),
.Y(n_1852)
);

NAND3xp33_ASAP7_75t_SL g1853 ( 
.A(n_1532),
.B(n_65),
.C(n_66),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1545),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_R g1855 ( 
.A(n_1728),
.B(n_1548),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1669),
.B(n_1537),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1693),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1727),
.B(n_1538),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1706),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1719),
.B(n_1495),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1799),
.A2(n_1666),
.B(n_1667),
.C(n_1837),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1737),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1798),
.Y(n_1863)
);

O2A1O1Ixp5_ASAP7_75t_SL g1864 ( 
.A1(n_1827),
.A2(n_1838),
.B(n_1793),
.C(n_1736),
.Y(n_1864)
);

A2O1A1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1674),
.A2(n_1795),
.B(n_1720),
.C(n_1803),
.Y(n_1865)
);

A2O1A1Ixp33_ASAP7_75t_L g1866 ( 
.A1(n_1675),
.A2(n_1542),
.B(n_1546),
.C(n_1549),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1741),
.B(n_1552),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1665),
.A2(n_1545),
.B(n_1629),
.Y(n_1868)
);

O2A1O1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1676),
.A2(n_1556),
.B(n_1557),
.C(n_1555),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1691),
.A2(n_1672),
.B(n_1712),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1690),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1686),
.B(n_1559),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1783),
.B(n_1696),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1764),
.B(n_1563),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1816),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1685),
.B(n_1568),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1714),
.B(n_1569),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1689),
.B(n_1495),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1721),
.B(n_67),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1671),
.B(n_1542),
.Y(n_1880)
);

O2A1O1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1811),
.A2(n_1571),
.B(n_1546),
.C(n_1564),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1761),
.B(n_1550),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1716),
.Y(n_1883)
);

A2O1A1Ixp33_ASAP7_75t_L g1884 ( 
.A1(n_1715),
.A2(n_1630),
.B(n_70),
.C(n_68),
.Y(n_1884)
);

A2O1A1Ixp33_ASAP7_75t_L g1885 ( 
.A1(n_1743),
.A2(n_71),
.B(n_68),
.C(n_69),
.Y(n_1885)
);

OAI21xp33_ASAP7_75t_SL g1886 ( 
.A1(n_1753),
.A2(n_69),
.B(n_72),
.Y(n_1886)
);

HB1xp67_ASAP7_75t_L g1887 ( 
.A(n_1789),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1802),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1832),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1702),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1682),
.B(n_76),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1668),
.A2(n_76),
.B(n_77),
.Y(n_1892)
);

OAI22x1_ASAP7_75t_L g1893 ( 
.A1(n_1820),
.A2(n_81),
.B1(n_78),
.B2(n_79),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1835),
.A2(n_82),
.B1(n_79),
.B2(n_81),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1697),
.A2(n_82),
.B(n_83),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1738),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1701),
.B(n_83),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1700),
.A2(n_84),
.B(n_85),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1681),
.A2(n_84),
.B(n_86),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1740),
.B(n_88),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1739),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1737),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1797),
.B(n_88),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1679),
.A2(n_89),
.B(n_90),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1673),
.A2(n_89),
.B(n_90),
.Y(n_1905)
);

OAI21x1_ASAP7_75t_L g1906 ( 
.A1(n_1688),
.A2(n_569),
.B(n_567),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1840),
.B(n_1852),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1792),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1683),
.B(n_91),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1725),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_1910)
);

BUFx4f_ASAP7_75t_SL g1911 ( 
.A(n_1806),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1733),
.A2(n_92),
.B(n_93),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1748),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_1913)
);

O2A1O1Ixp5_ASAP7_75t_L g1914 ( 
.A1(n_1777),
.A2(n_97),
.B(n_95),
.C(n_96),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1678),
.B(n_98),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1802),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1725),
.B(n_98),
.Y(n_1917)
);

OAI22xp5_ASAP7_75t_L g1918 ( 
.A1(n_1844),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1918)
);

NOR3xp33_ASAP7_75t_L g1919 ( 
.A(n_1776),
.B(n_100),
.C(n_101),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1745),
.B(n_102),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1752),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1816),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1699),
.Y(n_1923)
);

INVxp67_ASAP7_75t_L g1924 ( 
.A(n_1670),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1726),
.B(n_105),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1841),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1816),
.B(n_106),
.Y(n_1927)
);

BUFx4f_ASAP7_75t_L g1928 ( 
.A(n_1840),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1726),
.B(n_108),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1802),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1826),
.B(n_108),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1834),
.Y(n_1932)
);

AOI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1824),
.A2(n_112),
.B1(n_109),
.B2(n_110),
.C(n_113),
.Y(n_1933)
);

INVx1_ASAP7_75t_SL g1934 ( 
.A(n_1830),
.Y(n_1934)
);

NOR3xp33_ASAP7_75t_SL g1935 ( 
.A(n_1775),
.B(n_1790),
.C(n_1853),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_SL g1936 ( 
.A1(n_1822),
.A2(n_113),
.B1(n_109),
.B2(n_110),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1754),
.A2(n_114),
.B(n_115),
.Y(n_1937)
);

O2A1O1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1828),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1809),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1759),
.B(n_117),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1791),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1840),
.B(n_118),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1755),
.B(n_120),
.Y(n_1943)
);

BUFx4f_ASAP7_75t_SL g1944 ( 
.A(n_1809),
.Y(n_1944)
);

INVx4_ASAP7_75t_L g1945 ( 
.A(n_1839),
.Y(n_1945)
);

O2A1O1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1769),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_1946)
);

NAND3xp33_ASAP7_75t_SL g1947 ( 
.A(n_1850),
.B(n_1711),
.C(n_1713),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1788),
.A2(n_571),
.B(n_570),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1781),
.A2(n_124),
.B1(n_121),
.B2(n_123),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1746),
.A2(n_124),
.B(n_125),
.Y(n_1950)
);

A2O1A1Ixp33_ASAP7_75t_L g1951 ( 
.A1(n_1718),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1694),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1852),
.B(n_129),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1851),
.A2(n_1831),
.B(n_1829),
.C(n_1808),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_R g1955 ( 
.A(n_1768),
.B(n_572),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1804),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1787),
.B(n_129),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1817),
.A2(n_1717),
.B1(n_1786),
.B2(n_1779),
.Y(n_1958)
);

NOR3xp33_ASAP7_75t_SL g1959 ( 
.A(n_1823),
.B(n_130),
.C(n_131),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1810),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1767),
.B(n_130),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1852),
.B(n_131),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1804),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1809),
.Y(n_1964)
);

NOR2xp67_ASAP7_75t_SL g1965 ( 
.A(n_1804),
.B(n_132),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1825),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1846),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1847),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1848),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1762),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1763),
.B(n_132),
.Y(n_1971)
);

NAND3xp33_ASAP7_75t_L g1972 ( 
.A(n_1849),
.B(n_133),
.C(n_134),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1780),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1785),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1826),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1801),
.B(n_133),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1842),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1687),
.Y(n_1978)
);

A2O1A1Ixp33_ASAP7_75t_L g1979 ( 
.A1(n_1680),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1760),
.A2(n_138),
.B(n_139),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1818),
.B(n_139),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1826),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1698),
.B(n_140),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1707),
.Y(n_1984)
);

BUFx3_ASAP7_75t_L g1985 ( 
.A(n_1801),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1684),
.A2(n_140),
.B(n_141),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1801),
.B(n_141),
.Y(n_1987)
);

INVxp67_ASAP7_75t_L g1988 ( 
.A(n_1744),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1747),
.A2(n_142),
.B(n_143),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1695),
.B(n_142),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1677),
.A2(n_576),
.B(n_575),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1773),
.Y(n_1992)
);

A2O1A1Ixp33_ASAP7_75t_SL g1993 ( 
.A1(n_1813),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1815),
.B(n_144),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1703),
.A2(n_1692),
.B(n_1709),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1757),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1843),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1723),
.A2(n_146),
.B(n_147),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1730),
.Y(n_1999)
);

A2O1A1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1751),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1749),
.B(n_148),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1707),
.B(n_151),
.Y(n_2002)
);

O2A1O1Ixp5_ASAP7_75t_L g2003 ( 
.A1(n_1722),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1757),
.B(n_153),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1756),
.B(n_154),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1854),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1819),
.B(n_155),
.Y(n_2007)
);

INVx3_ASAP7_75t_L g2008 ( 
.A(n_1778),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1704),
.Y(n_2009)
);

OAI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1735),
.A2(n_155),
.B(n_156),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1757),
.B(n_156),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1723),
.A2(n_157),
.B(n_158),
.Y(n_2012)
);

OA22x2_ASAP7_75t_L g2013 ( 
.A1(n_1845),
.A2(n_161),
.B1(n_158),
.B2(n_159),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1836),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1770),
.A2(n_165),
.B1(n_162),
.B2(n_163),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1807),
.Y(n_2016)
);

O2A1O1Ixp33_ASAP7_75t_L g2017 ( 
.A1(n_1772),
.A2(n_166),
.B(n_162),
.C(n_165),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1771),
.Y(n_2018)
);

INVxp67_ASAP7_75t_SL g2019 ( 
.A(n_1784),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1765),
.B(n_1819),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_1819),
.B(n_167),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1778),
.A2(n_1805),
.B1(n_1774),
.B2(n_1796),
.Y(n_2022)
);

AND2x4_ASAP7_75t_L g2023 ( 
.A(n_1805),
.B(n_167),
.Y(n_2023)
);

CKINVDCx8_ASAP7_75t_R g2024 ( 
.A(n_1765),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1765),
.B(n_168),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_1758),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1731),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_2027)
);

OAI21x1_ASAP7_75t_L g2028 ( 
.A1(n_1870),
.A2(n_1995),
.B(n_1948),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1861),
.A2(n_1723),
.B(n_1742),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1924),
.B(n_169),
.Y(n_2030)
);

OAI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1865),
.A2(n_1800),
.B(n_1794),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_2008),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_2022),
.A2(n_1814),
.B(n_1812),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_1868),
.A2(n_1766),
.B(n_1821),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1887),
.Y(n_2035)
);

A2O1A1Ixp33_ASAP7_75t_L g2036 ( 
.A1(n_1983),
.A2(n_1833),
.B(n_1782),
.C(n_1750),
.Y(n_2036)
);

OAI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1885),
.A2(n_1729),
.B(n_1708),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1857),
.B(n_170),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1860),
.B(n_1724),
.Y(n_2039)
);

AND2x2_ASAP7_75t_SL g2040 ( 
.A(n_1871),
.B(n_1724),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1863),
.B(n_171),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_SL g2042 ( 
.A1(n_1954),
.A2(n_1705),
.B(n_1710),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1900),
.B(n_1724),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1913),
.A2(n_1734),
.B1(n_1732),
.B2(n_173),
.Y(n_2044)
);

OA21x2_ASAP7_75t_L g2045 ( 
.A1(n_2010),
.A2(n_171),
.B(n_172),
.Y(n_2045)
);

OAI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1972),
.A2(n_172),
.B(n_173),
.Y(n_2046)
);

O2A1O1Ixp5_ASAP7_75t_L g2047 ( 
.A1(n_1950),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1934),
.B(n_579),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_R g2049 ( 
.A(n_1955),
.B(n_174),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1872),
.B(n_175),
.Y(n_2050)
);

AO21x2_ASAP7_75t_L g2051 ( 
.A1(n_2010),
.A2(n_582),
.B(n_580),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1926),
.A2(n_180),
.B1(n_177),
.B2(n_178),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1876),
.B(n_177),
.Y(n_2053)
);

OAI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1991),
.A2(n_584),
.B(n_583),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1934),
.B(n_180),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1974),
.B(n_181),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_SL g2057 ( 
.A(n_1920),
.B(n_182),
.C(n_183),
.Y(n_2057)
);

AO21x2_ASAP7_75t_L g2058 ( 
.A1(n_2009),
.A2(n_2019),
.B(n_1992),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_2022),
.A2(n_182),
.B(n_183),
.Y(n_2059)
);

AOI21x1_ASAP7_75t_SL g2060 ( 
.A1(n_1994),
.A2(n_1897),
.B(n_1971),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1912),
.A2(n_184),
.B(n_186),
.Y(n_2061)
);

OA21x2_ASAP7_75t_L g2062 ( 
.A1(n_1914),
.A2(n_184),
.B(n_186),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1932),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_1908),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1859),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1891),
.A2(n_190),
.B1(n_187),
.B2(n_189),
.Y(n_2066)
);

BUFx10_ASAP7_75t_L g2067 ( 
.A(n_1862),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1856),
.B(n_187),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_2008),
.Y(n_2069)
);

OAI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1972),
.A2(n_189),
.B(n_190),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1970),
.B(n_191),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1878),
.B(n_191),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_2018),
.B(n_585),
.Y(n_2073)
);

OAI21x1_ASAP7_75t_L g2074 ( 
.A1(n_1906),
.A2(n_590),
.B(n_589),
.Y(n_2074)
);

OAI21x1_ASAP7_75t_L g2075 ( 
.A1(n_1905),
.A2(n_1904),
.B(n_1898),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1990),
.A2(n_192),
.B(n_193),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1999),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_1975),
.B(n_591),
.Y(n_2078)
);

AO31x2_ASAP7_75t_L g2079 ( 
.A1(n_1866),
.A2(n_593),
.A3(n_594),
.B(n_592),
.Y(n_2079)
);

INVxp67_ASAP7_75t_SL g2080 ( 
.A(n_1867),
.Y(n_2080)
);

AOI21xp33_ASAP7_75t_L g2081 ( 
.A1(n_1886),
.A2(n_1946),
.B(n_1993),
.Y(n_2081)
);

AO31x2_ASAP7_75t_L g2082 ( 
.A1(n_2016),
.A2(n_596),
.A3(n_597),
.B(n_595),
.Y(n_2082)
);

OA21x2_ASAP7_75t_L g2083 ( 
.A1(n_2006),
.A2(n_192),
.B(n_193),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1978),
.Y(n_2084)
);

BUFx2_ASAP7_75t_R g2085 ( 
.A(n_1902),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1973),
.B(n_194),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_1911),
.Y(n_2087)
);

OAI21x1_ASAP7_75t_L g2088 ( 
.A1(n_1895),
.A2(n_599),
.B(n_598),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1950),
.A2(n_194),
.B(n_195),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1968),
.B(n_195),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2002),
.B(n_196),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1969),
.B(n_196),
.Y(n_2092)
);

AO31x2_ASAP7_75t_L g2093 ( 
.A1(n_2014),
.A2(n_1883),
.A3(n_1901),
.B(n_1896),
.Y(n_2093)
);

OAI21x1_ASAP7_75t_L g2094 ( 
.A1(n_1989),
.A2(n_602),
.B(n_601),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1877),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1928),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_1930),
.Y(n_2097)
);

NAND4xp25_ASAP7_75t_SL g2098 ( 
.A(n_1910),
.B(n_199),
.C(n_197),
.D(n_198),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1882),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1967),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1930),
.B(n_603),
.Y(n_2101)
);

OAI21xp5_ASAP7_75t_SL g2102 ( 
.A1(n_1879),
.A2(n_197),
.B(n_198),
.Y(n_2102)
);

INVx5_ASAP7_75t_SL g2103 ( 
.A(n_1875),
.Y(n_2103)
);

BUFx10_ASAP7_75t_L g2104 ( 
.A(n_2005),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1858),
.B(n_199),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1960),
.Y(n_2106)
);

AOI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1899),
.A2(n_200),
.B(n_202),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1944),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1923),
.B(n_203),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1873),
.B(n_203),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_1880),
.A2(n_204),
.B(n_205),
.Y(n_2111)
);

OA21x2_ASAP7_75t_L g2112 ( 
.A1(n_2003),
.A2(n_205),
.B(n_206),
.Y(n_2112)
);

INVxp67_ASAP7_75t_L g2113 ( 
.A(n_1939),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_1981),
.A2(n_207),
.B(n_208),
.Y(n_2114)
);

NOR2xp67_ASAP7_75t_L g2115 ( 
.A(n_2026),
.B(n_604),
.Y(n_2115)
);

AOI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_1947),
.A2(n_207),
.B(n_208),
.Y(n_2116)
);

OAI21x1_ASAP7_75t_L g2117 ( 
.A1(n_1869),
.A2(n_608),
.B(n_605),
.Y(n_2117)
);

BUFx2_ASAP7_75t_R g2118 ( 
.A(n_2024),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1966),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1931),
.B(n_209),
.Y(n_2120)
);

OAI21x1_ASAP7_75t_L g2121 ( 
.A1(n_1892),
.A2(n_610),
.B(n_609),
.Y(n_2121)
);

OA21x2_ASAP7_75t_L g2122 ( 
.A1(n_1998),
.A2(n_210),
.B(n_211),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_1875),
.B(n_612),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1930),
.B(n_613),
.Y(n_2124)
);

NAND3xp33_ASAP7_75t_L g2125 ( 
.A(n_1935),
.B(n_210),
.C(n_211),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1915),
.B(n_212),
.Y(n_2126)
);

BUFx10_ASAP7_75t_L g2127 ( 
.A(n_2021),
.Y(n_2127)
);

AOI21x1_ASAP7_75t_SL g2128 ( 
.A1(n_1903),
.A2(n_212),
.B(n_213),
.Y(n_2128)
);

AOI221x1_ASAP7_75t_L g2129 ( 
.A1(n_1894),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.C(n_216),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1956),
.B(n_614),
.Y(n_2130)
);

AO31x2_ASAP7_75t_L g2131 ( 
.A1(n_1884),
.A2(n_616),
.A3(n_615),
.B(n_216),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_2000),
.A2(n_214),
.B(n_215),
.Y(n_2132)
);

A2O1A1Ixp33_ASAP7_75t_L g2133 ( 
.A1(n_1938),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_2020),
.Y(n_2134)
);

AOI21xp5_ASAP7_75t_L g2135 ( 
.A1(n_1986),
.A2(n_217),
.B(n_218),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_1881),
.A2(n_220),
.B(n_221),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1909),
.B(n_220),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1874),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1957),
.B(n_1940),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2001),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_R g2141 ( 
.A(n_1855),
.B(n_222),
.Y(n_2141)
);

AO21x2_ASAP7_75t_L g2142 ( 
.A1(n_1952),
.A2(n_223),
.B(n_224),
.Y(n_2142)
);

AOI21xp5_ASAP7_75t_L g2143 ( 
.A1(n_2026),
.A2(n_223),
.B(n_225),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1984),
.B(n_225),
.Y(n_2144)
);

CKINVDCx20_ASAP7_75t_R g2145 ( 
.A(n_2087),
.Y(n_2145)
);

BUFx12f_ASAP7_75t_L g2146 ( 
.A(n_2067),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2033),
.A2(n_2017),
.B(n_1936),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2077),
.B(n_2064),
.Y(n_2148)
);

AOI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_2031),
.A2(n_1936),
.B(n_1951),
.Y(n_2149)
);

BUFx12f_ASAP7_75t_L g2150 ( 
.A(n_2067),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2035),
.B(n_1943),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2065),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_2063),
.Y(n_2153)
);

AOI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2031),
.A2(n_1913),
.B(n_1928),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2093),
.Y(n_2155)
);

OAI221xp5_ASAP7_75t_L g2156 ( 
.A1(n_2102),
.A2(n_1889),
.B1(n_1961),
.B2(n_1921),
.C(n_1941),
.Y(n_2156)
);

NOR2xp67_ASAP7_75t_L g2157 ( 
.A(n_2030),
.B(n_1988),
.Y(n_2157)
);

OAI21xp5_ASAP7_75t_L g2158 ( 
.A1(n_2125),
.A2(n_1921),
.B(n_1979),
.Y(n_2158)
);

OAI21x1_ASAP7_75t_L g2159 ( 
.A1(n_2028),
.A2(n_1864),
.B(n_1980),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2064),
.B(n_2113),
.Y(n_2160)
);

A2O1A1Ixp33_ASAP7_75t_L g2161 ( 
.A1(n_2102),
.A2(n_1933),
.B(n_1959),
.C(n_1941),
.Y(n_2161)
);

OR2x4_ASAP7_75t_L g2162 ( 
.A(n_2057),
.B(n_1875),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2084),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2039),
.B(n_2023),
.Y(n_2164)
);

HB1xp67_ASAP7_75t_L g2165 ( 
.A(n_2058),
.Y(n_2165)
);

AO21x2_ASAP7_75t_L g2166 ( 
.A1(n_2029),
.A2(n_2012),
.B(n_1919),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2043),
.B(n_2023),
.Y(n_2167)
);

CKINVDCx11_ASAP7_75t_R g2168 ( 
.A(n_2104),
.Y(n_2168)
);

OAI21x1_ASAP7_75t_L g2169 ( 
.A1(n_2034),
.A2(n_1937),
.B(n_1907),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2100),
.Y(n_2170)
);

AOI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2052),
.A2(n_1893),
.B1(n_1894),
.B2(n_1918),
.C(n_1889),
.Y(n_2171)
);

INVx4_ASAP7_75t_L g2172 ( 
.A(n_2097),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2085),
.Y(n_2173)
);

BUFx8_ASAP7_75t_SL g2174 ( 
.A(n_2108),
.Y(n_2174)
);

OR2x6_ASAP7_75t_L g2175 ( 
.A(n_2042),
.B(n_1956),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_2104),
.B(n_1917),
.Y(n_2176)
);

INVx4_ASAP7_75t_L g2177 ( 
.A(n_2097),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_2096),
.Y(n_2178)
);

BUFx3_ASAP7_75t_L g2179 ( 
.A(n_2127),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2080),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2099),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2072),
.B(n_1927),
.Y(n_2182)
);

AO21x2_ASAP7_75t_L g2183 ( 
.A1(n_2058),
.A2(n_1997),
.B(n_1953),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_2125),
.B(n_1925),
.Y(n_2184)
);

OAI21x1_ASAP7_75t_L g2185 ( 
.A1(n_2059),
.A2(n_1916),
.B(n_1888),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_2117),
.A2(n_1963),
.B(n_1918),
.Y(n_2186)
);

CKINVDCx16_ASAP7_75t_R g2187 ( 
.A(n_2049),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_2118),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_2040),
.B(n_2026),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2095),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2106),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2126),
.B(n_1929),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2138),
.Y(n_2193)
);

OAI21x1_ASAP7_75t_L g2194 ( 
.A1(n_2075),
.A2(n_1963),
.B(n_1962),
.Y(n_2194)
);

O2A1O1Ixp33_ASAP7_75t_SL g2195 ( 
.A1(n_2046),
.A2(n_1942),
.B(n_1949),
.C(n_1976),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2140),
.Y(n_2196)
);

OAI21x1_ASAP7_75t_L g2197 ( 
.A1(n_2136),
.A2(n_2013),
.B(n_1958),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_2037),
.A2(n_1982),
.B(n_2027),
.Y(n_2198)
);

OAI21x1_ASAP7_75t_L g2199 ( 
.A1(n_2037),
.A2(n_2011),
.B(n_2004),
.Y(n_2199)
);

AOI22xp33_ASAP7_75t_L g2200 ( 
.A1(n_2046),
.A2(n_2070),
.B1(n_2098),
.B2(n_2052),
.Y(n_2200)
);

OAI21x1_ASAP7_75t_L g2201 ( 
.A1(n_2054),
.A2(n_2025),
.B(n_2007),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_2127),
.Y(n_2202)
);

O2A1O1Ixp33_ASAP7_75t_L g2203 ( 
.A1(n_2066),
.A2(n_1987),
.B(n_2015),
.C(n_1977),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2119),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2134),
.B(n_1931),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_2083),
.Y(n_2206)
);

AO21x1_ASAP7_75t_L g2207 ( 
.A1(n_2070),
.A2(n_1927),
.B(n_1945),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2139),
.B(n_1964),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_L g2209 ( 
.A1(n_2074),
.A2(n_1890),
.B(n_1965),
.Y(n_2209)
);

BUFx3_ASAP7_75t_L g2210 ( 
.A(n_2032),
.Y(n_2210)
);

OAI21x1_ASAP7_75t_L g2211 ( 
.A1(n_2128),
.A2(n_2094),
.B(n_2088),
.Y(n_2211)
);

OAI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2089),
.A2(n_1945),
.B(n_1985),
.Y(n_2212)
);

OAI21x1_ASAP7_75t_L g2213 ( 
.A1(n_2121),
.A2(n_1956),
.B(n_1996),
.Y(n_2213)
);

A2O1A1Ixp33_ASAP7_75t_L g2214 ( 
.A1(n_2044),
.A2(n_1922),
.B(n_1996),
.C(n_229),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2083),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2056),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2180),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2164),
.B(n_2032),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2152),
.Y(n_2219)
);

BUFx2_ASAP7_75t_L g2220 ( 
.A(n_2210),
.Y(n_2220)
);

BUFx2_ASAP7_75t_SL g2221 ( 
.A(n_2207),
.Y(n_2221)
);

NAND2x1p5_ASAP7_75t_L g2222 ( 
.A(n_2194),
.B(n_2045),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2155),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2200),
.A2(n_2044),
.B1(n_2133),
.B2(n_2045),
.Y(n_2224)
);

NAND2x1p5_ASAP7_75t_L g2225 ( 
.A(n_2186),
.B(n_2115),
.Y(n_2225)
);

NOR2x1_ASAP7_75t_SL g2226 ( 
.A(n_2175),
.B(n_2051),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_2156),
.A2(n_2142),
.B1(n_2081),
.B2(n_2051),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2171),
.A2(n_2200),
.B1(n_2161),
.B2(n_2184),
.Y(n_2228)
);

NOR2xp67_ASAP7_75t_SL g2229 ( 
.A(n_2149),
.B(n_2096),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2164),
.B(n_2069),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2161),
.A2(n_2141),
.B1(n_2142),
.B2(n_2116),
.Y(n_2231)
);

CKINVDCx20_ASAP7_75t_R g2232 ( 
.A(n_2174),
.Y(n_2232)
);

NAND2x1p5_ASAP7_75t_L g2233 ( 
.A(n_2185),
.B(n_2115),
.Y(n_2233)
);

OAI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_2154),
.A2(n_2129),
.B1(n_2132),
.B2(n_2135),
.Y(n_2234)
);

CKINVDCx5p33_ASAP7_75t_R g2235 ( 
.A(n_2174),
.Y(n_2235)
);

OA21x2_ASAP7_75t_L g2236 ( 
.A1(n_2165),
.A2(n_2143),
.B(n_2047),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2170),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_2175),
.Y(n_2238)
);

INVx6_ASAP7_75t_L g2239 ( 
.A(n_2146),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_2210),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_L g2241 ( 
.A1(n_2158),
.A2(n_2061),
.B1(n_2114),
.B2(n_2107),
.Y(n_2241)
);

BUFx3_ASAP7_75t_L g2242 ( 
.A(n_2146),
.Y(n_2242)
);

OAI21xp5_ASAP7_75t_SL g2243 ( 
.A1(n_2147),
.A2(n_2076),
.B(n_2111),
.Y(n_2243)
);

AOI22xp33_ASAP7_75t_L g2244 ( 
.A1(n_2184),
.A2(n_2122),
.B1(n_2048),
.B2(n_2112),
.Y(n_2244)
);

AO21x1_ASAP7_75t_L g2245 ( 
.A1(n_2189),
.A2(n_2215),
.B(n_2206),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2164),
.B(n_2069),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2214),
.A2(n_2048),
.B1(n_2120),
.B2(n_2091),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2214),
.A2(n_2137),
.B(n_2110),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2163),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2190),
.Y(n_2250)
);

AOI22xp33_ASAP7_75t_L g2251 ( 
.A1(n_2187),
.A2(n_2166),
.B1(n_2197),
.B2(n_2216),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2181),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2148),
.B(n_2055),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2151),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2160),
.Y(n_2255)
);

HB1xp67_ASAP7_75t_L g2256 ( 
.A(n_2196),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2191),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2204),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2167),
.B(n_2053),
.Y(n_2259)
);

INVx1_ASAP7_75t_SL g2260 ( 
.A(n_2168),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2256),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_2224),
.A2(n_2166),
.B1(n_2183),
.B2(n_2206),
.Y(n_2262)
);

INVxp67_ASAP7_75t_L g2263 ( 
.A(n_2221),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_2232),
.Y(n_2264)
);

AOI22xp33_ASAP7_75t_L g2265 ( 
.A1(n_2231),
.A2(n_2183),
.B1(n_2157),
.B2(n_2189),
.Y(n_2265)
);

OAI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_2228),
.A2(n_2162),
.B1(n_2202),
.B2(n_2179),
.Y(n_2266)
);

AO22x1_ASAP7_75t_L g2267 ( 
.A1(n_2248),
.A2(n_2188),
.B1(n_2173),
.B2(n_2176),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2255),
.B(n_2179),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2227),
.A2(n_2192),
.B1(n_2122),
.B2(n_2176),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2218),
.B(n_2153),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2260),
.B(n_2202),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2218),
.B(n_2153),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2254),
.B(n_2192),
.Y(n_2273)
);

AOI22xp33_ASAP7_75t_SL g2274 ( 
.A1(n_2221),
.A2(n_2226),
.B1(n_2236),
.B2(n_2222),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_2234),
.A2(n_2182),
.B1(n_2112),
.B2(n_2062),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2217),
.B(n_2199),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_SL g2277 ( 
.A1(n_2226),
.A2(n_2188),
.B1(n_2165),
.B2(n_2175),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2251),
.A2(n_2062),
.B1(n_2205),
.B2(n_2193),
.Y(n_2278)
);

OAI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_2247),
.A2(n_2162),
.B1(n_2212),
.B2(n_2036),
.Y(n_2279)
);

AOI22xp33_ASAP7_75t_SL g2280 ( 
.A1(n_2236),
.A2(n_2159),
.B1(n_2105),
.B2(n_2050),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_2242),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2223),
.Y(n_2282)
);

BUFx6f_ASAP7_75t_L g2283 ( 
.A(n_2242),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2217),
.B(n_2208),
.Y(n_2284)
);

AOI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_2241),
.A2(n_2198),
.B1(n_2201),
.B2(n_2209),
.Y(n_2285)
);

OAI21xp33_ASAP7_75t_L g2286 ( 
.A1(n_2243),
.A2(n_2041),
.B(n_2038),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_2263),
.B(n_2230),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_R g2288 ( 
.A(n_2264),
.B(n_2232),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2264),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_2281),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2261),
.Y(n_2291)
);

NAND2xp33_ASAP7_75t_R g2292 ( 
.A(n_2268),
.B(n_2235),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_R g2293 ( 
.A(n_2281),
.B(n_2235),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2268),
.B(n_2220),
.Y(n_2294)
);

XNOR2xp5_ASAP7_75t_L g2295 ( 
.A(n_2267),
.B(n_2145),
.Y(n_2295)
);

BUFx10_ASAP7_75t_L g2296 ( 
.A(n_2281),
.Y(n_2296)
);

BUFx10_ASAP7_75t_L g2297 ( 
.A(n_2281),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2290),
.B(n_2274),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2291),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_2290),
.B(n_2262),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2294),
.B(n_2287),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2296),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_2296),
.Y(n_2303)
);

BUFx6f_ASAP7_75t_L g2304 ( 
.A(n_2296),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2301),
.B(n_2287),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2301),
.B(n_2298),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2299),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2299),
.B(n_2280),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2299),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2301),
.B(n_2287),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2302),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2298),
.B(n_2294),
.Y(n_2312)
);

OAI22xp33_ASAP7_75t_L g2313 ( 
.A1(n_2300),
.A2(n_2279),
.B1(n_2266),
.B2(n_2292),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2302),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2309),
.Y(n_2315)
);

INVxp67_ASAP7_75t_L g2316 ( 
.A(n_2306),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2306),
.B(n_2298),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2312),
.B(n_2302),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2309),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2308),
.B(n_2273),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2307),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2314),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2305),
.B(n_2302),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2314),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2310),
.B(n_2303),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2311),
.B(n_2303),
.Y(n_2326)
);

INVxp67_ASAP7_75t_L g2327 ( 
.A(n_2317),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2315),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2317),
.B(n_2303),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2318),
.B(n_2303),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2316),
.B(n_2303),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2325),
.B(n_2304),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2319),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2322),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_2323),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2324),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2335),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_SL g2338 ( 
.A(n_2335),
.B(n_2313),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2335),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2332),
.Y(n_2340)
);

BUFx2_ASAP7_75t_L g2341 ( 
.A(n_2340),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2339),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2337),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_2338),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2341),
.Y(n_2345)
);

XNOR2x1_ASAP7_75t_L g2346 ( 
.A(n_2343),
.B(n_2320),
.Y(n_2346)
);

OAI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2344),
.A2(n_2338),
.B1(n_2327),
.B2(n_2313),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2341),
.B(n_2329),
.Y(n_2348)
);

OAI21xp33_ASAP7_75t_SL g2349 ( 
.A1(n_2342),
.A2(n_2329),
.B(n_2330),
.Y(n_2349)
);

AOI22xp33_ASAP7_75t_L g2350 ( 
.A1(n_2344),
.A2(n_2308),
.B1(n_2300),
.B2(n_2334),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2349),
.B(n_2331),
.Y(n_2351)
);

BUFx2_ASAP7_75t_SL g2352 ( 
.A(n_2345),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_L g2353 ( 
.A(n_2348),
.B(n_2331),
.C(n_2336),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2346),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2347),
.Y(n_2355)
);

AOI22xp5_ASAP7_75t_L g2356 ( 
.A1(n_2350),
.A2(n_2318),
.B1(n_2333),
.B2(n_2328),
.Y(n_2356)
);

OAI322xp33_ASAP7_75t_L g2357 ( 
.A1(n_2347),
.A2(n_2321),
.A3(n_2326),
.B1(n_2330),
.B2(n_2331),
.C1(n_2325),
.C2(n_2295),
.Y(n_2357)
);

NAND3xp33_ASAP7_75t_L g2358 ( 
.A(n_2345),
.B(n_2332),
.C(n_2326),
.Y(n_2358)
);

AOI32xp33_ASAP7_75t_L g2359 ( 
.A1(n_2347),
.A2(n_2332),
.A3(n_2300),
.B1(n_2323),
.B2(n_2286),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2348),
.B(n_2323),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2352),
.Y(n_2361)
);

OAI21xp5_ASAP7_75t_SL g2362 ( 
.A1(n_2351),
.A2(n_2300),
.B(n_2304),
.Y(n_2362)
);

A2O1A1Ixp33_ASAP7_75t_L g2363 ( 
.A1(n_2359),
.A2(n_2300),
.B(n_2289),
.C(n_2269),
.Y(n_2363)
);

OAI22xp33_ASAP7_75t_L g2364 ( 
.A1(n_2354),
.A2(n_2300),
.B1(n_2304),
.B2(n_2283),
.Y(n_2364)
);

INVx2_ASAP7_75t_SL g2365 ( 
.A(n_2360),
.Y(n_2365)
);

OAI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2358),
.A2(n_2086),
.B(n_2071),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2353),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2356),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2357),
.A2(n_2355),
.B(n_2289),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2352),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2352),
.B(n_2288),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2352),
.Y(n_2372)
);

INVx1_ASAP7_75t_SL g2373 ( 
.A(n_2360),
.Y(n_2373)
);

NOR3xp33_ASAP7_75t_L g2374 ( 
.A(n_2373),
.B(n_2267),
.C(n_2168),
.Y(n_2374)
);

INVx2_ASAP7_75t_SL g2375 ( 
.A(n_2371),
.Y(n_2375)
);

INVx2_ASAP7_75t_SL g2376 ( 
.A(n_2365),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2361),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2362),
.B(n_2367),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2370),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2372),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2368),
.Y(n_2381)
);

NOR3x1_ASAP7_75t_L g2382 ( 
.A(n_2362),
.B(n_2271),
.C(n_2092),
.Y(n_2382)
);

AOI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2369),
.A2(n_2145),
.B(n_2304),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2366),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2364),
.B(n_2239),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2363),
.B(n_2304),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2373),
.B(n_2304),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2362),
.A2(n_2304),
.B(n_2283),
.Y(n_2388)
);

OAI211xp5_ASAP7_75t_L g2389 ( 
.A1(n_2378),
.A2(n_2293),
.B(n_2304),
.C(n_2283),
.Y(n_2389)
);

OAI221xp5_ASAP7_75t_L g2390 ( 
.A1(n_2374),
.A2(n_2239),
.B1(n_2304),
.B2(n_2281),
.C(n_2283),
.Y(n_2390)
);

AOI21xp33_ASAP7_75t_L g2391 ( 
.A1(n_2381),
.A2(n_2090),
.B(n_2068),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2376),
.B(n_2283),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2387),
.Y(n_2393)
);

HAxp5_ASAP7_75t_SL g2394 ( 
.A(n_2379),
.B(n_2239),
.CON(n_2394),
.SN(n_2394)
);

AOI221xp5_ASAP7_75t_L g2395 ( 
.A1(n_2384),
.A2(n_2265),
.B1(n_2245),
.B2(n_2285),
.C(n_2195),
.Y(n_2395)
);

OAI21xp5_ASAP7_75t_SL g2396 ( 
.A1(n_2383),
.A2(n_2277),
.B(n_2109),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2386),
.A2(n_2276),
.B(n_2195),
.Y(n_2397)
);

OAI211xp5_ASAP7_75t_SL g2398 ( 
.A1(n_2377),
.A2(n_2275),
.B(n_229),
.C(n_227),
.Y(n_2398)
);

OAI22xp5_ASAP7_75t_L g2399 ( 
.A1(n_2380),
.A2(n_2375),
.B1(n_2385),
.B2(n_2388),
.Y(n_2399)
);

AOI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2382),
.A2(n_2245),
.B1(n_2278),
.B2(n_2244),
.C(n_2203),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2382),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2376),
.Y(n_2402)
);

AOI321xp33_ASAP7_75t_L g2403 ( 
.A1(n_2399),
.A2(n_2144),
.A3(n_2078),
.B1(n_2073),
.B2(n_2101),
.C(n_2130),
.Y(n_2403)
);

OAI211xp5_ASAP7_75t_L g2404 ( 
.A1(n_2402),
.A2(n_230),
.B(n_227),
.C(n_228),
.Y(n_2404)
);

AOI321xp33_ASAP7_75t_L g2405 ( 
.A1(n_2401),
.A2(n_2078),
.A3(n_2124),
.B1(n_2123),
.B2(n_2253),
.C(n_2060),
.Y(n_2405)
);

OAI221xp5_ASAP7_75t_L g2406 ( 
.A1(n_2393),
.A2(n_2239),
.B1(n_2253),
.B2(n_2229),
.C(n_2222),
.Y(n_2406)
);

O2A1O1Ixp33_ASAP7_75t_SL g2407 ( 
.A1(n_2389),
.A2(n_2390),
.B(n_2397),
.C(n_2391),
.Y(n_2407)
);

O2A1O1Ixp33_ASAP7_75t_L g2408 ( 
.A1(n_2392),
.A2(n_2259),
.B(n_232),
.C(n_230),
.Y(n_2408)
);

AOI211xp5_ASAP7_75t_L g2409 ( 
.A1(n_2398),
.A2(n_2229),
.B(n_2211),
.C(n_2123),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2396),
.B(n_2297),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_2394),
.B(n_2150),
.Y(n_2411)
);

AOI222xp33_ASAP7_75t_L g2412 ( 
.A1(n_2395),
.A2(n_2150),
.B1(n_2297),
.B2(n_2284),
.C1(n_2252),
.C2(n_2250),
.Y(n_2412)
);

O2A1O1Ixp33_ASAP7_75t_L g2413 ( 
.A1(n_2400),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2413)
);

NAND3xp33_ASAP7_75t_L g2414 ( 
.A(n_2394),
.B(n_2096),
.C(n_2236),
.Y(n_2414)
);

O2A1O1Ixp33_ASAP7_75t_L g2415 ( 
.A1(n_2399),
.A2(n_235),
.B(n_233),
.C(n_234),
.Y(n_2415)
);

O2A1O1Ixp33_ASAP7_75t_L g2416 ( 
.A1(n_2399),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_2416)
);

OAI21x1_ASAP7_75t_L g2417 ( 
.A1(n_2399),
.A2(n_2272),
.B(n_2270),
.Y(n_2417)
);

AOI211xp5_ASAP7_75t_L g2418 ( 
.A1(n_2401),
.A2(n_239),
.B(n_237),
.C(n_238),
.Y(n_2418)
);

NAND4xp75_ASAP7_75t_L g2419 ( 
.A(n_2402),
.B(n_241),
.C(n_238),
.D(n_240),
.Y(n_2419)
);

OAI321xp33_ASAP7_75t_L g2420 ( 
.A1(n_2401),
.A2(n_2233),
.A3(n_2225),
.B1(n_2222),
.B2(n_2257),
.C(n_2238),
.Y(n_2420)
);

AOI21xp5_ASAP7_75t_L g2421 ( 
.A1(n_2399),
.A2(n_2272),
.B(n_2270),
.Y(n_2421)
);

AOI211x1_ASAP7_75t_SL g2422 ( 
.A1(n_2399),
.A2(n_2297),
.B(n_244),
.C(n_240),
.Y(n_2422)
);

OAI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2393),
.A2(n_2219),
.B1(n_2249),
.B2(n_2237),
.Y(n_2423)
);

AOI22xp5_ASAP7_75t_L g2424 ( 
.A1(n_2401),
.A2(n_2178),
.B1(n_2225),
.B2(n_2220),
.Y(n_2424)
);

AOI322xp5_ASAP7_75t_L g2425 ( 
.A1(n_2411),
.A2(n_2131),
.A3(n_2258),
.B1(n_2282),
.B2(n_2082),
.C1(n_2178),
.C2(n_2079),
.Y(n_2425)
);

AOI211x1_ASAP7_75t_SL g2426 ( 
.A1(n_2410),
.A2(n_246),
.B(n_243),
.C(n_244),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2404),
.B(n_243),
.Y(n_2427)
);

OAI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2424),
.A2(n_2178),
.B1(n_2225),
.B2(n_2233),
.Y(n_2428)
);

AOI221xp5_ASAP7_75t_L g2429 ( 
.A1(n_2413),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.C(n_249),
.Y(n_2429)
);

AOI221xp5_ASAP7_75t_L g2430 ( 
.A1(n_2407),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_2430)
);

AOI222xp33_ASAP7_75t_L g2431 ( 
.A1(n_2414),
.A2(n_2420),
.B1(n_2406),
.B2(n_2417),
.C1(n_2422),
.C2(n_2412),
.Y(n_2431)
);

AOI221xp5_ASAP7_75t_L g2432 ( 
.A1(n_2408),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.C(n_255),
.Y(n_2432)
);

AOI221xp5_ASAP7_75t_L g2433 ( 
.A1(n_2415),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.C(n_255),
.Y(n_2433)
);

INVxp67_ASAP7_75t_L g2434 ( 
.A(n_2419),
.Y(n_2434)
);

OAI211xp5_ASAP7_75t_L g2435 ( 
.A1(n_2416),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_2435)
);

OAI211xp5_ASAP7_75t_L g2436 ( 
.A1(n_2418),
.A2(n_260),
.B(n_257),
.C(n_259),
.Y(n_2436)
);

XOR2x2_ASAP7_75t_L g2437 ( 
.A(n_2409),
.B(n_259),
.Y(n_2437)
);

OAI21xp33_ASAP7_75t_L g2438 ( 
.A1(n_2421),
.A2(n_2240),
.B(n_2230),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_R g2439 ( 
.A(n_2403),
.B(n_260),
.Y(n_2439)
);

OAI222xp33_ASAP7_75t_L g2440 ( 
.A1(n_2423),
.A2(n_2233),
.B1(n_2172),
.B2(n_2177),
.C1(n_2240),
.C2(n_2246),
.Y(n_2440)
);

AOI21xp5_ASAP7_75t_L g2441 ( 
.A1(n_2405),
.A2(n_261),
.B(n_262),
.Y(n_2441)
);

NOR3xp33_ASAP7_75t_L g2442 ( 
.A(n_2404),
.B(n_261),
.C(n_262),
.Y(n_2442)
);

AOI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2411),
.A2(n_2178),
.B1(n_2246),
.B2(n_2240),
.Y(n_2443)
);

NAND2xp33_ASAP7_75t_SL g2444 ( 
.A(n_2410),
.B(n_263),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2422),
.Y(n_2445)
);

OAI211xp5_ASAP7_75t_L g2446 ( 
.A1(n_2415),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_2446)
);

NOR3xp33_ASAP7_75t_L g2447 ( 
.A(n_2404),
.B(n_266),
.C(n_267),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2411),
.B(n_2238),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2422),
.B(n_2131),
.Y(n_2449)
);

A2O1A1Ixp33_ASAP7_75t_L g2450 ( 
.A1(n_2411),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_2450)
);

NAND3xp33_ASAP7_75t_L g2451 ( 
.A(n_2418),
.B(n_1996),
.C(n_268),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2422),
.B(n_2131),
.Y(n_2452)
);

AOI221xp5_ASAP7_75t_L g2453 ( 
.A1(n_2413),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.C(n_272),
.Y(n_2453)
);

OAI221xp5_ASAP7_75t_L g2454 ( 
.A1(n_2411),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.C(n_272),
.Y(n_2454)
);

OAI221xp5_ASAP7_75t_L g2455 ( 
.A1(n_2411),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.C(n_276),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2411),
.B(n_2238),
.Y(n_2456)
);

OAI211xp5_ASAP7_75t_L g2457 ( 
.A1(n_2415),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2457)
);

NOR4xp25_ASAP7_75t_L g2458 ( 
.A(n_2407),
.B(n_279),
.C(n_277),
.D(n_278),
.Y(n_2458)
);

OAI211xp5_ASAP7_75t_SL g2459 ( 
.A1(n_2422),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_2459)
);

AOI222xp33_ASAP7_75t_L g2460 ( 
.A1(n_2414),
.A2(n_2282),
.B1(n_2082),
.B2(n_282),
.C1(n_283),
.C2(n_284),
.Y(n_2460)
);

NOR2x1_ASAP7_75t_L g2461 ( 
.A(n_2419),
.B(n_280),
.Y(n_2461)
);

OAI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2449),
.A2(n_2238),
.B1(n_2172),
.B2(n_2177),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2426),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2461),
.Y(n_2464)
);

NAND4xp75_ASAP7_75t_L g2465 ( 
.A(n_2430),
.B(n_282),
.C(n_280),
.D(n_281),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2445),
.Y(n_2466)
);

NOR2x1_ASAP7_75t_L g2467 ( 
.A(n_2454),
.B(n_2455),
.Y(n_2467)
);

NOR2xp67_ASAP7_75t_SL g2468 ( 
.A(n_2436),
.B(n_284),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2434),
.Y(n_2469)
);

NAND4xp25_ASAP7_75t_L g2470 ( 
.A(n_2459),
.B(n_287),
.C(n_285),
.D(n_286),
.Y(n_2470)
);

NOR3xp33_ASAP7_75t_L g2471 ( 
.A(n_2444),
.B(n_285),
.C(n_288),
.Y(n_2471)
);

NAND3xp33_ASAP7_75t_L g2472 ( 
.A(n_2450),
.B(n_288),
.C(n_289),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2452),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_2458),
.B(n_290),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_L g2475 ( 
.A(n_2435),
.B(n_292),
.C(n_293),
.Y(n_2475)
);

AOI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2442),
.A2(n_2447),
.B1(n_2427),
.B2(n_2431),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2446),
.Y(n_2477)
);

AO22x1_ASAP7_75t_L g2478 ( 
.A1(n_2457),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2451),
.Y(n_2479)
);

NAND3xp33_ASAP7_75t_L g2480 ( 
.A(n_2433),
.B(n_295),
.C(n_296),
.Y(n_2480)
);

AOI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2432),
.A2(n_2103),
.B1(n_2238),
.B2(n_2213),
.Y(n_2481)
);

OAI221xp5_ASAP7_75t_L g2482 ( 
.A1(n_2441),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.C(n_298),
.Y(n_2482)
);

NOR3xp33_ASAP7_75t_L g2483 ( 
.A(n_2429),
.B(n_297),
.C(n_298),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2437),
.Y(n_2484)
);

NAND3xp33_ASAP7_75t_L g2485 ( 
.A(n_2453),
.B(n_299),
.C(n_300),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2439),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2448),
.Y(n_2487)
);

NOR2x1_ASAP7_75t_L g2488 ( 
.A(n_2456),
.B(n_299),
.Y(n_2488)
);

OAI21xp33_ASAP7_75t_L g2489 ( 
.A1(n_2443),
.A2(n_301),
.B(n_302),
.Y(n_2489)
);

OAI21xp5_ASAP7_75t_SL g2490 ( 
.A1(n_2460),
.A2(n_301),
.B(n_302),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2438),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2428),
.Y(n_2492)
);

NAND3xp33_ASAP7_75t_L g2493 ( 
.A(n_2425),
.B(n_303),
.C(n_304),
.Y(n_2493)
);

NOR2x1_ASAP7_75t_L g2494 ( 
.A(n_2440),
.B(n_306),
.Y(n_2494)
);

NAND4xp75_ASAP7_75t_L g2495 ( 
.A(n_2461),
.B(n_308),
.C(n_306),
.D(n_307),
.Y(n_2495)
);

NOR2x1_ASAP7_75t_L g2496 ( 
.A(n_2445),
.B(n_307),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2426),
.Y(n_2497)
);

NOR3xp33_ASAP7_75t_L g2498 ( 
.A(n_2444),
.B(n_309),
.C(n_310),
.Y(n_2498)
);

INVx2_ASAP7_75t_SL g2499 ( 
.A(n_2461),
.Y(n_2499)
);

NOR2x1_ASAP7_75t_L g2500 ( 
.A(n_2495),
.B(n_310),
.Y(n_2500)
);

NAND4xp75_ASAP7_75t_L g2501 ( 
.A(n_2496),
.B(n_313),
.C(n_311),
.D(n_312),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2463),
.Y(n_2502)
);

NAND4xp75_ASAP7_75t_L g2503 ( 
.A(n_2499),
.B(n_314),
.C(n_312),
.D(n_313),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2474),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2470),
.B(n_314),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2497),
.B(n_2082),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2478),
.B(n_316),
.Y(n_2507)
);

NOR2x1_ASAP7_75t_L g2508 ( 
.A(n_2464),
.B(n_317),
.Y(n_2508)
);

NAND3x2_ASAP7_75t_L g2509 ( 
.A(n_2466),
.B(n_317),
.C(n_318),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2465),
.Y(n_2510)
);

OA21x2_ASAP7_75t_L g2511 ( 
.A1(n_2469),
.A2(n_318),
.B(n_319),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2477),
.B(n_2487),
.Y(n_2512)
);

NAND3xp33_ASAP7_75t_L g2513 ( 
.A(n_2486),
.B(n_2476),
.C(n_2471),
.Y(n_2513)
);

OAI211xp5_ASAP7_75t_L g2514 ( 
.A1(n_2489),
.A2(n_321),
.B(n_319),
.C(n_320),
.Y(n_2514)
);

NAND4xp25_ASAP7_75t_L g2515 ( 
.A(n_2498),
.B(n_323),
.C(n_321),
.D(n_322),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2468),
.Y(n_2516)
);

NOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2473),
.B(n_323),
.Y(n_2517)
);

NAND3xp33_ASAP7_75t_L g2518 ( 
.A(n_2484),
.B(n_324),
.C(n_325),
.Y(n_2518)
);

NOR2xp67_ASAP7_75t_L g2519 ( 
.A(n_2472),
.B(n_324),
.Y(n_2519)
);

NAND3x1_ASAP7_75t_L g2520 ( 
.A(n_2494),
.B(n_325),
.C(n_326),
.Y(n_2520)
);

NAND2xp33_ASAP7_75t_SL g2521 ( 
.A(n_2491),
.B(n_327),
.Y(n_2521)
);

NOR3xp33_ASAP7_75t_L g2522 ( 
.A(n_2479),
.B(n_327),
.C(n_328),
.Y(n_2522)
);

NOR2x1_ASAP7_75t_L g2523 ( 
.A(n_2485),
.B(n_329),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_L g2524 ( 
.A(n_2488),
.B(n_329),
.C(n_330),
.Y(n_2524)
);

NOR2x1_ASAP7_75t_L g2525 ( 
.A(n_2480),
.B(n_2482),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2475),
.B(n_330),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2490),
.B(n_331),
.Y(n_2527)
);

NOR3xp33_ASAP7_75t_L g2528 ( 
.A(n_2467),
.B(n_331),
.C(n_332),
.Y(n_2528)
);

NOR3x2_ASAP7_75t_L g2529 ( 
.A(n_2483),
.B(n_332),
.C(n_333),
.Y(n_2529)
);

AOI21xp5_ASAP7_75t_L g2530 ( 
.A1(n_2492),
.A2(n_334),
.B(n_335),
.Y(n_2530)
);

NOR2x1_ASAP7_75t_L g2531 ( 
.A(n_2493),
.B(n_335),
.Y(n_2531)
);

NOR2x1_ASAP7_75t_L g2532 ( 
.A(n_2462),
.B(n_336),
.Y(n_2532)
);

INVxp67_ASAP7_75t_L g2533 ( 
.A(n_2481),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2481),
.Y(n_2534)
);

NOR3x1_ASAP7_75t_L g2535 ( 
.A(n_2495),
.B(n_336),
.C(n_337),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2499),
.B(n_337),
.Y(n_2536)
);

CKINVDCx20_ASAP7_75t_R g2537 ( 
.A(n_2469),
.Y(n_2537)
);

NOR3xp33_ASAP7_75t_L g2538 ( 
.A(n_2469),
.B(n_338),
.C(n_339),
.Y(n_2538)
);

NAND2xp33_ASAP7_75t_L g2539 ( 
.A(n_2469),
.B(n_338),
.Y(n_2539)
);

NOR3xp33_ASAP7_75t_L g2540 ( 
.A(n_2469),
.B(n_339),
.C(n_340),
.Y(n_2540)
);

INVxp67_ASAP7_75t_SL g2541 ( 
.A(n_2496),
.Y(n_2541)
);

INVxp67_ASAP7_75t_L g2542 ( 
.A(n_2496),
.Y(n_2542)
);

INVx1_ASAP7_75t_SL g2543 ( 
.A(n_2495),
.Y(n_2543)
);

NAND3xp33_ASAP7_75t_L g2544 ( 
.A(n_2469),
.B(n_340),
.C(n_341),
.Y(n_2544)
);

NOR3xp33_ASAP7_75t_L g2545 ( 
.A(n_2469),
.B(n_341),
.C(n_342),
.Y(n_2545)
);

NOR3x1_ASAP7_75t_L g2546 ( 
.A(n_2495),
.B(n_343),
.C(n_344),
.Y(n_2546)
);

INVx3_ASAP7_75t_L g2547 ( 
.A(n_2495),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2463),
.B(n_345),
.Y(n_2548)
);

INVxp33_ASAP7_75t_SL g2549 ( 
.A(n_2469),
.Y(n_2549)
);

NOR3xp33_ASAP7_75t_L g2550 ( 
.A(n_2469),
.B(n_345),
.C(n_346),
.Y(n_2550)
);

NOR2x1_ASAP7_75t_L g2551 ( 
.A(n_2495),
.B(n_347),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2496),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2496),
.Y(n_2553)
);

NAND3xp33_ASAP7_75t_SL g2554 ( 
.A(n_2469),
.B(n_348),
.C(n_349),
.Y(n_2554)
);

NAND4xp75_ASAP7_75t_L g2555 ( 
.A(n_2496),
.B(n_349),
.C(n_350),
.D(n_351),
.Y(n_2555)
);

NOR3xp33_ASAP7_75t_L g2556 ( 
.A(n_2469),
.B(n_351),
.C(n_352),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2470),
.B(n_352),
.Y(n_2557)
);

NOR2x1_ASAP7_75t_L g2558 ( 
.A(n_2495),
.B(n_353),
.Y(n_2558)
);

NOR3xp33_ASAP7_75t_L g2559 ( 
.A(n_2469),
.B(n_353),
.C(n_354),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2499),
.B(n_354),
.Y(n_2560)
);

XNOR2x1_ASAP7_75t_L g2561 ( 
.A(n_2469),
.B(n_355),
.Y(n_2561)
);

NAND4xp75_ASAP7_75t_L g2562 ( 
.A(n_2517),
.B(n_355),
.C(n_356),
.D(n_357),
.Y(n_2562)
);

NAND4xp75_ASAP7_75t_L g2563 ( 
.A(n_2508),
.B(n_2512),
.C(n_2553),
.D(n_2552),
.Y(n_2563)
);

AOI22xp33_ASAP7_75t_L g2564 ( 
.A1(n_2537),
.A2(n_2103),
.B1(n_2213),
.B2(n_1922),
.Y(n_2564)
);

INVx1_ASAP7_75t_SL g2565 ( 
.A(n_2529),
.Y(n_2565)
);

OAI221xp5_ASAP7_75t_L g2566 ( 
.A1(n_2502),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.C(n_359),
.Y(n_2566)
);

XNOR2x1_ASAP7_75t_L g2567 ( 
.A(n_2561),
.B(n_358),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2511),
.Y(n_2568)
);

OA22x2_ASAP7_75t_L g2569 ( 
.A1(n_2504),
.A2(n_360),
.B1(n_361),
.B2(n_363),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2549),
.B(n_363),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2513),
.B(n_364),
.Y(n_2571)
);

NAND4xp75_ASAP7_75t_L g2572 ( 
.A(n_2535),
.B(n_364),
.C(n_365),
.D(n_366),
.Y(n_2572)
);

INVx2_ASAP7_75t_SL g2573 ( 
.A(n_2500),
.Y(n_2573)
);

OAI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2520),
.A2(n_2169),
.B(n_365),
.Y(n_2574)
);

AOI211xp5_ASAP7_75t_L g2575 ( 
.A1(n_2554),
.A2(n_366),
.B(n_367),
.C(n_368),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2541),
.B(n_368),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2511),
.Y(n_2577)
);

XNOR2xp5_ASAP7_75t_L g2578 ( 
.A(n_2509),
.B(n_369),
.Y(n_2578)
);

AND3x4_ASAP7_75t_L g2579 ( 
.A(n_2524),
.B(n_370),
.C(n_371),
.Y(n_2579)
);

AO21x1_ASAP7_75t_L g2580 ( 
.A1(n_2521),
.A2(n_370),
.B(n_372),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_R g2581 ( 
.A(n_2547),
.B(n_372),
.Y(n_2581)
);

OR2x6_ASAP7_75t_L g2582 ( 
.A(n_2542),
.B(n_373),
.Y(n_2582)
);

XNOR2x1_ASAP7_75t_L g2583 ( 
.A(n_2501),
.B(n_2555),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2551),
.Y(n_2584)
);

NOR5xp2_ASAP7_75t_SL g2585 ( 
.A(n_2548),
.B(n_374),
.C(n_376),
.D(n_377),
.E(n_378),
.Y(n_2585)
);

XNOR2x1_ASAP7_75t_L g2586 ( 
.A(n_2558),
.B(n_374),
.Y(n_2586)
);

NAND4xp75_ASAP7_75t_L g2587 ( 
.A(n_2546),
.B(n_376),
.C(n_377),
.D(n_378),
.Y(n_2587)
);

NAND3xp33_ASAP7_75t_SL g2588 ( 
.A(n_2543),
.B(n_379),
.C(n_380),
.Y(n_2588)
);

AOI21x1_ASAP7_75t_L g2589 ( 
.A1(n_2560),
.A2(n_380),
.B(n_381),
.Y(n_2589)
);

INVx1_ASAP7_75t_SL g2590 ( 
.A(n_2507),
.Y(n_2590)
);

OAI322xp33_ASAP7_75t_L g2591 ( 
.A1(n_2516),
.A2(n_381),
.A3(n_382),
.B1(n_383),
.B2(n_384),
.C1(n_385),
.C2(n_386),
.Y(n_2591)
);

AOI221xp5_ASAP7_75t_SL g2592 ( 
.A1(n_2539),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.C(n_385),
.Y(n_2592)
);

NAND4xp75_ASAP7_75t_L g2593 ( 
.A(n_2531),
.B(n_387),
.C(n_388),
.D(n_389),
.Y(n_2593)
);

OAI21xp33_ASAP7_75t_L g2594 ( 
.A1(n_2515),
.A2(n_387),
.B(n_388),
.Y(n_2594)
);

NAND3x1_ASAP7_75t_L g2595 ( 
.A(n_2536),
.B(n_390),
.C(n_391),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2547),
.B(n_393),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2503),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_SL g2598 ( 
.A(n_2510),
.B(n_393),
.Y(n_2598)
);

NAND4xp25_ASAP7_75t_SL g2599 ( 
.A(n_2528),
.B(n_394),
.C(n_395),
.D(n_396),
.Y(n_2599)
);

OR2x2_ASAP7_75t_L g2600 ( 
.A(n_2505),
.B(n_395),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_2519),
.Y(n_2601)
);

OAI211xp5_ASAP7_75t_L g2602 ( 
.A1(n_2527),
.A2(n_396),
.B(n_397),
.C(n_398),
.Y(n_2602)
);

AOI311xp33_ASAP7_75t_L g2603 ( 
.A1(n_2534),
.A2(n_397),
.A3(n_399),
.B(n_400),
.C(n_401),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2557),
.Y(n_2604)
);

NOR2x1_ASAP7_75t_SL g2605 ( 
.A(n_2514),
.B(n_2544),
.Y(n_2605)
);

OAI32xp33_ASAP7_75t_L g2606 ( 
.A1(n_2526),
.A2(n_399),
.A3(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_2606)
);

NOR2xp67_ASAP7_75t_SL g2607 ( 
.A(n_2518),
.B(n_403),
.Y(n_2607)
);

BUFx2_ASAP7_75t_L g2608 ( 
.A(n_2523),
.Y(n_2608)
);

NOR2x1_ASAP7_75t_L g2609 ( 
.A(n_2530),
.B(n_404),
.Y(n_2609)
);

NOR2x1_ASAP7_75t_L g2610 ( 
.A(n_2525),
.B(n_404),
.Y(n_2610)
);

NAND5xp2_ASAP7_75t_L g2611 ( 
.A(n_2533),
.B(n_405),
.C(n_406),
.D(n_407),
.E(n_408),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2538),
.Y(n_2612)
);

INVx1_ASAP7_75t_SL g2613 ( 
.A(n_2532),
.Y(n_2613)
);

NOR2xp67_ASAP7_75t_L g2614 ( 
.A(n_2506),
.B(n_405),
.Y(n_2614)
);

AND2x4_ASAP7_75t_L g2615 ( 
.A(n_2540),
.B(n_2545),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2550),
.Y(n_2616)
);

NAND4xp75_ASAP7_75t_L g2617 ( 
.A(n_2522),
.B(n_2556),
.C(n_2559),
.D(n_409),
.Y(n_2617)
);

AOI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2549),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.C(n_410),
.Y(n_2618)
);

NOR2x1_ASAP7_75t_L g2619 ( 
.A(n_2537),
.B(n_411),
.Y(n_2619)
);

NAND4xp25_ASAP7_75t_L g2620 ( 
.A(n_2549),
.B(n_411),
.C(n_412),
.D(n_413),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2549),
.B(n_412),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2512),
.B(n_414),
.Y(n_2622)
);

NAND3x1_ASAP7_75t_L g2623 ( 
.A(n_2508),
.B(n_415),
.C(n_416),
.Y(n_2623)
);

NOR3xp33_ASAP7_75t_L g2624 ( 
.A(n_2513),
.B(n_415),
.C(n_416),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2549),
.B(n_417),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2537),
.B(n_417),
.Y(n_2626)
);

NAND4xp75_ASAP7_75t_L g2627 ( 
.A(n_2517),
.B(n_418),
.C(n_419),
.D(n_420),
.Y(n_2627)
);

NOR3x2_ASAP7_75t_L g2628 ( 
.A(n_2501),
.B(n_418),
.C(n_419),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_R g2629 ( 
.A(n_2570),
.B(n_420),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2581),
.B(n_421),
.Y(n_2630)
);

NAND2xp33_ASAP7_75t_SL g2631 ( 
.A(n_2621),
.B(n_421),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_R g2632 ( 
.A(n_2625),
.B(n_422),
.Y(n_2632)
);

NOR2xp33_ASAP7_75t_R g2633 ( 
.A(n_2588),
.B(n_422),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2573),
.B(n_423),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_R g2635 ( 
.A(n_2599),
.B(n_423),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_R g2636 ( 
.A(n_2584),
.B(n_424),
.Y(n_2636)
);

NAND2xp33_ASAP7_75t_SL g2637 ( 
.A(n_2622),
.B(n_424),
.Y(n_2637)
);

NAND2xp33_ASAP7_75t_SL g2638 ( 
.A(n_2607),
.B(n_425),
.Y(n_2638)
);

NAND2xp33_ASAP7_75t_SL g2639 ( 
.A(n_2583),
.B(n_426),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_R g2640 ( 
.A(n_2589),
.B(n_426),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_R g2641 ( 
.A(n_2596),
.B(n_427),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2568),
.B(n_427),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_R g2643 ( 
.A(n_2578),
.B(n_428),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_R g2644 ( 
.A(n_2577),
.B(n_429),
.Y(n_2644)
);

NAND2xp33_ASAP7_75t_SL g2645 ( 
.A(n_2586),
.B(n_429),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_R g2646 ( 
.A(n_2598),
.B(n_430),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_2603),
.B(n_431),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_R g2648 ( 
.A(n_2600),
.B(n_431),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_SL g2649 ( 
.A(n_2613),
.B(n_432),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2601),
.B(n_432),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_R g2651 ( 
.A(n_2608),
.B(n_433),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_SL g2652 ( 
.A(n_2571),
.B(n_434),
.Y(n_2652)
);

NOR2xp33_ASAP7_75t_R g2653 ( 
.A(n_2597),
.B(n_2612),
.Y(n_2653)
);

NAND3xp33_ASAP7_75t_L g2654 ( 
.A(n_2610),
.B(n_435),
.C(n_436),
.Y(n_2654)
);

NAND3xp33_ASAP7_75t_L g2655 ( 
.A(n_2619),
.B(n_435),
.C(n_436),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_R g2656 ( 
.A(n_2616),
.B(n_438),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2592),
.B(n_438),
.Y(n_2657)
);

NAND2xp33_ASAP7_75t_SL g2658 ( 
.A(n_2579),
.B(n_439),
.Y(n_2658)
);

NAND2xp33_ASAP7_75t_SL g2659 ( 
.A(n_2567),
.B(n_439),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_R g2660 ( 
.A(n_2604),
.B(n_440),
.Y(n_2660)
);

NAND3xp33_ASAP7_75t_L g2661 ( 
.A(n_2624),
.B(n_441),
.C(n_443),
.Y(n_2661)
);

NOR3xp33_ASAP7_75t_SL g2662 ( 
.A(n_2563),
.B(n_441),
.C(n_444),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2580),
.B(n_444),
.Y(n_2663)
);

NOR3xp33_ASAP7_75t_SL g2664 ( 
.A(n_2572),
.B(n_445),
.C(n_447),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2614),
.B(n_445),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2590),
.B(n_448),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_2575),
.B(n_448),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2565),
.B(n_449),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2626),
.B(n_449),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_R g2670 ( 
.A(n_2576),
.B(n_450),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2576),
.B(n_451),
.Y(n_2671)
);

XNOR2xp5_ASAP7_75t_L g2672 ( 
.A(n_2623),
.B(n_452),
.Y(n_2672)
);

NAND3xp33_ASAP7_75t_L g2673 ( 
.A(n_2609),
.B(n_453),
.C(n_454),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2615),
.B(n_453),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_R g2675 ( 
.A(n_2585),
.B(n_455),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2582),
.B(n_455),
.Y(n_2676)
);

XNOR2xp5_ASAP7_75t_L g2677 ( 
.A(n_2628),
.B(n_456),
.Y(n_2677)
);

XNOR2xp5_ASAP7_75t_L g2678 ( 
.A(n_2595),
.B(n_457),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_R g2679 ( 
.A(n_2611),
.B(n_458),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_R g2680 ( 
.A(n_2587),
.B(n_458),
.Y(n_2680)
);

NAND3xp33_ASAP7_75t_L g2681 ( 
.A(n_2602),
.B(n_459),
.C(n_460),
.Y(n_2681)
);

NOR3xp33_ASAP7_75t_SL g2682 ( 
.A(n_2617),
.B(n_459),
.C(n_460),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_R g2683 ( 
.A(n_2569),
.B(n_461),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_R g2684 ( 
.A(n_2620),
.B(n_461),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2594),
.B(n_462),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2645),
.A2(n_2593),
.B1(n_2562),
.B2(n_2627),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2678),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2672),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2677),
.Y(n_2689)
);

INVxp33_ASAP7_75t_SL g2690 ( 
.A(n_2643),
.Y(n_2690)
);

BUFx2_ASAP7_75t_L g2691 ( 
.A(n_2675),
.Y(n_2691)
);

AOI22xp5_ASAP7_75t_L g2692 ( 
.A1(n_2647),
.A2(n_2566),
.B1(n_2574),
.B2(n_2618),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2665),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2663),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2671),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2676),
.Y(n_2696)
);

HB1xp67_ASAP7_75t_L g2697 ( 
.A(n_2679),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2642),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2670),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2654),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2655),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2662),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2669),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2630),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2673),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2666),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2653),
.B(n_2582),
.Y(n_2707)
);

CKINVDCx20_ASAP7_75t_R g2708 ( 
.A(n_2659),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2650),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2637),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2668),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2658),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2657),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2664),
.Y(n_2714)
);

BUFx6f_ASAP7_75t_L g2715 ( 
.A(n_2674),
.Y(n_2715)
);

OR3x2_ASAP7_75t_L g2716 ( 
.A(n_2648),
.B(n_2605),
.C(n_2606),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2682),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2652),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2640),
.Y(n_2719)
);

CKINVDCx20_ASAP7_75t_R g2720 ( 
.A(n_2631),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2639),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2644),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2651),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2634),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2649),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_2685),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2667),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2636),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2699),
.Y(n_2729)
);

AOI22xp5_ASAP7_75t_L g2730 ( 
.A1(n_2691),
.A2(n_2638),
.B1(n_2661),
.B2(n_2681),
.Y(n_2730)
);

XNOR2x1_ASAP7_75t_L g2731 ( 
.A(n_2697),
.B(n_2641),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_L g2732 ( 
.A(n_2690),
.B(n_2591),
.Y(n_2732)
);

XOR2xp5_ASAP7_75t_L g2733 ( 
.A(n_2719),
.B(n_2629),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2723),
.Y(n_2734)
);

XOR2xp5_ASAP7_75t_L g2735 ( 
.A(n_2716),
.B(n_2632),
.Y(n_2735)
);

XNOR2xp5_ASAP7_75t_SL g2736 ( 
.A(n_2686),
.B(n_2714),
.Y(n_2736)
);

OA22x2_ASAP7_75t_L g2737 ( 
.A1(n_2692),
.A2(n_2683),
.B1(n_2660),
.B2(n_2684),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2715),
.Y(n_2738)
);

AO22x2_ASAP7_75t_L g2739 ( 
.A1(n_2710),
.A2(n_2656),
.B1(n_2646),
.B2(n_2680),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2715),
.Y(n_2740)
);

AOI22xp5_ASAP7_75t_L g2741 ( 
.A1(n_2702),
.A2(n_2564),
.B1(n_2635),
.B2(n_2633),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2715),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2707),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2720),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2708),
.Y(n_2745)
);

AO22x2_ASAP7_75t_L g2746 ( 
.A1(n_2721),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.Y(n_2746)
);

XNOR2x1_ASAP7_75t_L g2747 ( 
.A(n_2687),
.B(n_464),
.Y(n_2747)
);

INVx2_ASAP7_75t_SL g2748 ( 
.A(n_2713),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2722),
.B(n_465),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2726),
.Y(n_2750)
);

AOI22x1_ASAP7_75t_L g2751 ( 
.A1(n_2688),
.A2(n_466),
.B1(n_467),
.B2(n_468),
.Y(n_2751)
);

XNOR2xp5_ASAP7_75t_L g2752 ( 
.A(n_2689),
.B(n_467),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2712),
.Y(n_2753)
);

OA22x2_ASAP7_75t_L g2754 ( 
.A1(n_2717),
.A2(n_468),
.B1(n_469),
.B2(n_470),
.Y(n_2754)
);

INVxp67_ASAP7_75t_SL g2755 ( 
.A(n_2694),
.Y(n_2755)
);

BUFx3_ASAP7_75t_L g2756 ( 
.A(n_2728),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2706),
.Y(n_2757)
);

AND2x4_ASAP7_75t_L g2758 ( 
.A(n_2755),
.B(n_2718),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2738),
.B(n_2693),
.Y(n_2759)
);

AO21x2_ASAP7_75t_L g2760 ( 
.A1(n_2740),
.A2(n_2696),
.B(n_2711),
.Y(n_2760)
);

OAI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2748),
.A2(n_2704),
.B(n_2724),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2739),
.Y(n_2762)
);

OA22x2_ASAP7_75t_L g2763 ( 
.A1(n_2735),
.A2(n_2733),
.B1(n_2730),
.B2(n_2744),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2739),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2742),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2750),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2737),
.Y(n_2767)
);

XNOR2xp5_ASAP7_75t_L g2768 ( 
.A(n_2731),
.B(n_2736),
.Y(n_2768)
);

XNOR2xp5_ASAP7_75t_L g2769 ( 
.A(n_2745),
.B(n_2709),
.Y(n_2769)
);

AOI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2729),
.A2(n_2695),
.B1(n_2701),
.B2(n_2700),
.Y(n_2770)
);

OAI21x1_ASAP7_75t_L g2771 ( 
.A1(n_2734),
.A2(n_2725),
.B(n_2705),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2757),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2752),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2747),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2756),
.B(n_2698),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2749),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2746),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2753),
.A2(n_2703),
.B1(n_2727),
.B2(n_2726),
.Y(n_2778)
);

CKINVDCx20_ASAP7_75t_R g2779 ( 
.A(n_2768),
.Y(n_2779)
);

OAI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2758),
.A2(n_2743),
.B(n_2732),
.Y(n_2780)
);

XOR2xp5_ASAP7_75t_L g2781 ( 
.A(n_2769),
.B(n_2741),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2766),
.B(n_2754),
.Y(n_2782)
);

BUFx2_ASAP7_75t_L g2783 ( 
.A(n_2761),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2760),
.Y(n_2784)
);

NOR3xp33_ASAP7_75t_L g2785 ( 
.A(n_2775),
.B(n_2726),
.C(n_2751),
.Y(n_2785)
);

OAI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2771),
.A2(n_2746),
.B(n_472),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2772),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2777),
.Y(n_2788)
);

OAI22x1_ASAP7_75t_L g2789 ( 
.A1(n_2770),
.A2(n_471),
.B1(n_473),
.B2(n_474),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2763),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2759),
.A2(n_471),
.B(n_475),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2779),
.Y(n_2792)
);

BUFx2_ASAP7_75t_L g2793 ( 
.A(n_2783),
.Y(n_2793)
);

INVxp67_ASAP7_75t_L g2794 ( 
.A(n_2790),
.Y(n_2794)
);

OAI22xp5_ASAP7_75t_SL g2795 ( 
.A1(n_2781),
.A2(n_2765),
.B1(n_2762),
.B2(n_2764),
.Y(n_2795)
);

AO22x2_ASAP7_75t_L g2796 ( 
.A1(n_2784),
.A2(n_2778),
.B1(n_2767),
.B2(n_2773),
.Y(n_2796)
);

INVx1_ASAP7_75t_SL g2797 ( 
.A(n_2787),
.Y(n_2797)
);

XOR2xp5_ASAP7_75t_L g2798 ( 
.A(n_2780),
.B(n_2774),
.Y(n_2798)
);

CKINVDCx20_ASAP7_75t_R g2799 ( 
.A(n_2788),
.Y(n_2799)
);

HB1xp67_ASAP7_75t_L g2800 ( 
.A(n_2782),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2793),
.B(n_2786),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2792),
.B(n_2776),
.Y(n_2802)
);

INVxp67_ASAP7_75t_L g2803 ( 
.A(n_2800),
.Y(n_2803)
);

XOR2xp5_ASAP7_75t_L g2804 ( 
.A(n_2798),
.B(n_2789),
.Y(n_2804)
);

OR2x6_ASAP7_75t_L g2805 ( 
.A(n_2795),
.B(n_2785),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2794),
.A2(n_2791),
.B(n_476),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2803),
.Y(n_2807)
);

OAI22xp5_ASAP7_75t_SL g2808 ( 
.A1(n_2805),
.A2(n_2799),
.B1(n_2797),
.B2(n_2796),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2801),
.Y(n_2809)
);

OAI22xp5_ASAP7_75t_L g2810 ( 
.A1(n_2802),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_2810)
);

NAND3xp33_ASAP7_75t_L g2811 ( 
.A(n_2807),
.B(n_2806),
.C(n_2804),
.Y(n_2811)
);

OAI21xp5_ASAP7_75t_L g2812 ( 
.A1(n_2809),
.A2(n_478),
.B(n_479),
.Y(n_2812)
);

AOI33xp33_ASAP7_75t_L g2813 ( 
.A1(n_2811),
.A2(n_2808),
.A3(n_2810),
.B1(n_480),
.B2(n_481),
.B3(n_482),
.Y(n_2813)
);

AOI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2813),
.A2(n_2812),
.B1(n_479),
.B2(n_481),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2814),
.B(n_478),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2815),
.A2(n_482),
.B(n_483),
.Y(n_2816)
);

AOI211xp5_ASAP7_75t_L g2817 ( 
.A1(n_2816),
.A2(n_483),
.B(n_484),
.C(n_485),
.Y(n_2817)
);


endmodule