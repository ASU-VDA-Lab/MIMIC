module fake_jpeg_167_n_183 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_183);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_66),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_51),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_52),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_58),
.B1(n_65),
.B2(n_57),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_61),
.B(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_50),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_65),
.B1(n_57),
.B2(n_52),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_91),
.B1(n_64),
.B2(n_61),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_63),
.B(n_60),
.C(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_107),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_80),
.B1(n_81),
.B2(n_59),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_103),
.A2(n_101),
.B1(n_88),
.B2(n_92),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_7),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_62),
.B1(n_22),
.B2(n_24),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_4),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g119 ( 
.A(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_1),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_21),
.B(n_45),
.C(n_44),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_33),
.B(n_41),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_0),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_121),
.B(n_2),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_123),
.B(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_1),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_128),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_3),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_5),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_6),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_138),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_139),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_9),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_137),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_12),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_12),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_13),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_113),
.B(n_13),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_141),
.B(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_14),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_131),
.B(n_133),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_108),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_31),
.C(n_40),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_138),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_113),
.B1(n_122),
.B2(n_135),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_156),
.B1(n_143),
.B2(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_153),
.C(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_29),
.C(n_39),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_27),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_169),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_171),
.B1(n_156),
.B2(n_165),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_154),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_171),
.B1(n_143),
.B2(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_157),
.B(n_152),
.C(n_168),
.Y(n_176)
);

AOI31xp67_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_176),
.A3(n_173),
.B(n_174),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_14),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_15),
.C(n_16),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_25),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_34),
.B(n_38),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_46),
.Y(n_183)
);


endmodule