module fake_jpeg_20975_n_31 (n_3, n_2, n_1, n_0, n_4, n_5, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_1),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_18),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_11),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_6),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_16),
.A2(n_17),
.B1(n_9),
.B2(n_10),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_8),
.A2(n_2),
.B1(n_5),
.B2(n_10),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_13),
.C(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_22),
.A2(n_9),
.B(n_16),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_25),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_20),
.B(n_21),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_19),
.C(n_20),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_29),
.C(n_13),
.Y(n_31)
);


endmodule