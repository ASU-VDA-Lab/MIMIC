module fake_jpeg_7991_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_47),
.B1(n_64),
.B2(n_68),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_19),
.B1(n_34),
.B2(n_20),
.Y(n_47)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_53),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_65),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_20),
.B1(n_19),
.B2(n_34),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_32),
.B(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_26),
.B1(n_29),
.B2(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_74),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_43),
.C(n_23),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_86),
.C(n_25),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_25),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_21),
.B(n_18),
.Y(n_99)
);

AO21x2_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_24),
.B(n_43),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_43),
.C(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_90),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_34),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_17),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_49),
.B1(n_58),
.B2(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_115),
.B1(n_93),
.B2(n_95),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_46),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_97),
.A2(n_121),
.B(n_28),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_103),
.B1(n_121),
.B2(n_21),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_48),
.B1(n_60),
.B2(n_69),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_17),
.B1(n_31),
.B2(n_22),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_105),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_33),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_113),
.C(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_111),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_70),
.C(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_49),
.B1(n_48),
.B2(n_69),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_29),
.B1(n_31),
.B2(n_21),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_27),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_17),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_96),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_78),
.B1(n_70),
.B2(n_79),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_131),
.B1(n_136),
.B2(n_143),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_144),
.B(n_9),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_78),
.B1(n_79),
.B2(n_26),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_130),
.A2(n_145),
.B1(n_123),
.B2(n_114),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_76),
.B1(n_73),
.B2(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_151),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_31),
.C(n_17),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_139),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_80),
.B1(n_28),
.B2(n_27),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_27),
.B1(n_29),
.B2(n_18),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_110),
.B1(n_98),
.B2(n_100),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_18),
.B1(n_30),
.B2(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_104),
.B(n_107),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_146),
.A2(n_98),
.B1(n_100),
.B2(n_105),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_158),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_104),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_102),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_162),
.C(n_166),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_136),
.B1(n_145),
.B2(n_127),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_101),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_164),
.B(n_170),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_109),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_112),
.A3(n_115),
.B1(n_33),
.B2(n_30),
.C1(n_31),
.C2(n_22),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_130),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_22),
.B(n_112),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_171),
.B(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_22),
.B(n_1),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_128),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_179),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_180),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_112),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_177),
.B1(n_169),
.B2(n_176),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_156),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_191),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_195),
.Y(n_212)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_137),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_195),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_132),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_197),
.C(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_134),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_134),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_136),
.B1(n_146),
.B2(n_140),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_204),
.B1(n_165),
.B2(n_172),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_171),
.B(n_136),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_160),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_146),
.B1(n_22),
.B2(n_2),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_0),
.C(n_1),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_212),
.B(n_215),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_170),
.C(n_158),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_225),
.C(n_228),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_177),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_218),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_168),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_222),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_174),
.B1(n_173),
.B2(n_153),
.Y(n_220)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_229),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_231),
.B1(n_234),
.B2(n_232),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_165),
.C(n_161),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_161),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_189),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_16),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_185),
.B(n_191),
.C(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_182),
.C(n_185),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_182),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_0),
.B(n_3),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_213),
.B(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_245),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_183),
.C(n_189),
.Y(n_244)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_250),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_203),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_184),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_202),
.C(n_181),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_205),
.C(n_204),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_217),
.C(n_211),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_207),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_10),
.B(n_15),
.C(n_14),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_257),
.A2(n_231),
.B1(n_221),
.B2(n_11),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_228),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_210),
.C(n_216),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_264),
.C(n_268),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_232),
.C(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_16),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_240),
.B1(n_238),
.B2(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_0),
.C(n_3),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_274),
.C(n_4),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_4),
.C(n_5),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_259),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_280),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_274),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_288),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_245),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_283),
.C(n_12),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_247),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_273),
.A2(n_243),
.B1(n_249),
.B2(n_255),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_284),
.A2(n_286),
.B1(n_290),
.B2(n_285),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_257),
.B1(n_12),
.B2(n_13),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_289),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_16),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_290),
.B(n_5),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_263),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_291),
.B(n_300),
.Y(n_312)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_262),
.B1(n_272),
.B2(n_261),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_5),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_268),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_299),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_270),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_12),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_277),
.A2(n_259),
.B(n_270),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_13),
.B(n_14),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_303),
.B(n_297),
.C(n_294),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_305),
.B(n_307),
.Y(n_320)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_7),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_6),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_6),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_302),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_300),
.B1(n_7),
.B2(n_8),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_7),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_7),
.B(n_8),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_320),
.B(n_308),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_326),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_305),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_327),
.B(n_323),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_325),
.C(n_311),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_316),
.B(n_307),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_316),
.Y(n_332)
);


endmodule