module fake_jpeg_4641_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_15),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_28),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_61),
.Y(n_81)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_63),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_71),
.Y(n_115)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_77),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_23),
.B1(n_46),
.B2(n_48),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_91),
.B1(n_93),
.B2(n_36),
.Y(n_111)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_85),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_80)
);

OAI22x1_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_87),
.B1(n_94),
.B2(n_99),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_60),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_17),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_46),
.B1(n_40),
.B2(n_45),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_58),
.B1(n_54),
.B2(n_38),
.Y(n_110)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_51),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_41),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_46),
.B1(n_37),
.B2(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g122 ( 
.A(n_92),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_48),
.B1(n_39),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_29),
.B1(n_19),
.B2(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_53),
.A2(n_19),
.B1(n_29),
.B2(n_37),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_104),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_55),
.B1(n_38),
.B2(n_45),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_110),
.B1(n_79),
.B2(n_96),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_44),
.B(n_26),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_108),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_22),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_29),
.B1(n_19),
.B2(n_34),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_105),
.A2(n_111),
.B1(n_32),
.B2(n_31),
.Y(n_156)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_107),
.A2(n_113),
.B1(n_119),
.B2(n_125),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_44),
.B(n_27),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_117),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_40),
.B(n_38),
.C(n_45),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_120),
.B1(n_58),
.B2(n_20),
.Y(n_154)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_47),
.C(n_67),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_40),
.B1(n_30),
.B2(n_36),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_71),
.A2(n_17),
.B1(n_28),
.B2(n_34),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_119),
.A2(n_98),
.B1(n_88),
.B2(n_83),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_151),
.B1(n_154),
.B2(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_140),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_97),
.C(n_28),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_132),
.B(n_25),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_133),
.A2(n_143),
.B(n_150),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_88),
.B(n_72),
.C(n_77),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_112),
.B(n_47),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_106),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_138),
.A2(n_139),
.B1(n_147),
.B2(n_32),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_95),
.B1(n_76),
.B2(n_75),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_149),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_125),
.B(n_107),
.Y(n_142)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_148),
.B(n_25),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_76),
.B1(n_75),
.B2(n_40),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_30),
.B(n_34),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_31),
.C(n_33),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_30),
.B1(n_58),
.B2(n_54),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_158),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

FAx1_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_112),
.CI(n_110),
.CON(n_159),
.SN(n_159)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_159),
.A2(n_171),
.B(n_176),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_145),
.A2(n_112),
.B1(n_123),
.B2(n_113),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_170),
.B(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_67),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_67),
.Y(n_164)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_167),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_86),
.C(n_112),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_178),
.C(n_131),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_123),
.B1(n_100),
.B2(n_31),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_R g171 ( 
.A(n_143),
.B(n_31),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_33),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

NAND2x1p5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_24),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_86),
.C(n_118),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_54),
.B(n_24),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g210 ( 
.A1(n_181),
.A2(n_24),
.B1(n_32),
.B2(n_129),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_0),
.Y(n_221)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_140),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_151),
.B1(n_134),
.B2(n_138),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_25),
.A3(n_32),
.B1(n_24),
.B2(n_27),
.C1(n_26),
.C2(n_11),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_14),
.Y(n_214)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_158),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_194),
.B(n_200),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_139),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_198),
.C(n_201),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_148),
.Y(n_198)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_163),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_203),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_163),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_206),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_152),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_208),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_149),
.B(n_146),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_172),
.B1(n_168),
.B2(n_181),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_118),
.C(n_27),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_14),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_13),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_13),
.B(n_12),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_179),
.B1(n_187),
.B2(n_184),
.Y(n_227)
);

AOI22x1_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_176),
.B1(n_159),
.B2(n_190),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_223),
.A2(n_227),
.B1(n_237),
.B2(n_238),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_173),
.B1(n_182),
.B2(n_186),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_231),
.B1(n_239),
.B2(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_232),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_176),
.B1(n_174),
.B2(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_159),
.B1(n_165),
.B2(n_181),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_159),
.B1(n_160),
.B2(n_181),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_162),
.B(n_191),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_198),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_196),
.A2(n_170),
.B1(n_180),
.B2(n_183),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_197),
.A2(n_191),
.B1(n_188),
.B2(n_166),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_220),
.B1(n_205),
.B2(n_222),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_195),
.A2(n_167),
.B1(n_1),
.B2(n_3),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_209),
.B1(n_194),
.B2(n_204),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_246),
.B(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_0),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_201),
.C(n_207),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_261),
.C(n_265),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_199),
.B(n_205),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_259),
.B1(n_246),
.B2(n_238),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_211),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_223),
.B(n_216),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_258),
.B(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_243),
.B1(n_235),
.B2(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_218),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_222),
.B1(n_215),
.B2(n_217),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_215),
.B1(n_214),
.B2(n_4),
.Y(n_263)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_224),
.B(n_13),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_12),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_237),
.B(n_244),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_1),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_233),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_236),
.A2(n_1),
.B(n_3),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_270),
.A2(n_226),
.B(n_247),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_272),
.A2(n_273),
.B(n_277),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_227),
.B1(n_225),
.B2(n_240),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_276),
.B1(n_250),
.B2(n_266),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_225),
.B1(n_233),
.B2(n_228),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_10),
.B(n_9),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_10),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

AOI221xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_287),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_261),
.C(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_4),
.C(n_5),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_7),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_254),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_5),
.B(n_6),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_267),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_297),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_293),
.B(n_302),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_258),
.B1(n_249),
.B2(n_264),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_299),
.B1(n_283),
.B2(n_272),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_257),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_254),
.B1(n_9),
.B2(n_6),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_4),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_286),
.C(n_284),
.Y(n_305)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_287),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_311),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_314),
.C(n_304),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_283),
.B1(n_284),
.B2(n_7),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_298),
.B1(n_297),
.B2(n_289),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_7),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_8),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_311),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_309),
.CI(n_314),
.CON(n_317),
.SN(n_317)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_317),
.B(n_321),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_322),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_305),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_324),
.A2(n_319),
.B(n_318),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_323),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

NOR2x1_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_317),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_317),
.Y(n_331)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

NOR3x1_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_330),
.C(n_325),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_334),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_332),
.B(n_331),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_328),
.Y(n_340)
);


endmodule