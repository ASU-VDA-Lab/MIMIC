module fake_jpeg_21498_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_19),
.B(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_31),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_52),
.B(n_53),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_24),
.B1(n_31),
.B2(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_58),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_24),
.B1(n_18),
.B2(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_24),
.B1(n_18),
.B2(n_33),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_27),
.B1(n_32),
.B2(n_17),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_17),
.B1(n_29),
.B2(n_20),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_28),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_38),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_20),
.B(n_29),
.C(n_26),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_38),
.B(n_2),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_25),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_3),
.B(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_66),
.A2(n_68),
.B1(n_64),
.B2(n_61),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_37),
.B1(n_40),
.B2(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_70),
.B(n_79),
.Y(n_117)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_40),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_35),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_83),
.A2(n_100),
.B1(n_101),
.B2(n_64),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_88),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_42),
.B1(n_21),
.B2(n_28),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_89),
.B1(n_92),
.B2(n_97),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_28),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_21),
.B1(n_38),
.B2(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_22),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_22),
.B1(n_32),
.B2(n_21),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_1),
.C(n_2),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_44),
.B(n_3),
.C(n_5),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_15),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_108),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_57),
.B1(n_53),
.B2(n_62),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_68),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_66),
.Y(n_134)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_57),
.B1(n_62),
.B2(n_56),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_126),
.B1(n_83),
.B2(n_72),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_115),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_73),
.B(n_80),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_111),
.B1(n_128),
.B2(n_105),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_134),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_137),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_83),
.B1(n_67),
.B2(n_94),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_77),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_139),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_87),
.B(n_82),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_148),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_92),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_152),
.C(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_79),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_111),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_127),
.B1(n_120),
.B2(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_75),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_96),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_112),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_153),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_69),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_98),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_162),
.B(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_163),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_116),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_154),
.B1(n_137),
.B2(n_148),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_132),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_120),
.B1(n_114),
.B2(n_108),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_143),
.B1(n_136),
.B2(n_129),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_112),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_178),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_114),
.C(n_104),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_159),
.C(n_155),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_182),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_196),
.B1(n_163),
.B2(n_158),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_193),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_154),
.B1(n_131),
.B2(n_151),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_190),
.A2(n_192),
.B1(n_166),
.B2(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_142),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_182),
.B(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_178),
.B(n_164),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_152),
.B1(n_140),
.B2(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_189),
.B(n_169),
.C(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_204),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_176),
.C(n_168),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_179),
.C(n_193),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_177),
.B1(n_170),
.B2(n_158),
.Y(n_203)
);

AOI211xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_157),
.B(n_163),
.C(n_161),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_208),
.A2(n_187),
.B1(n_181),
.B2(n_195),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_140),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_212),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_216),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_196),
.B(n_184),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_173),
.C(n_104),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_204),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_188),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_138),
.B1(n_167),
.B2(n_85),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_81),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_222),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_198),
.B1(n_203),
.B2(n_202),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_215),
.B1(n_212),
.B2(n_211),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_200),
.Y(n_238)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_240),
.B(n_242),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_214),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_217),
.B(n_220),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_216),
.B(n_14),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_228),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_231),
.B1(n_232),
.B2(n_228),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_241),
.B1(n_12),
.B2(n_10),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_250),
.Y(n_252)
);

NOR4xp25_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_15),
.C(n_8),
.D(n_9),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_243),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_7),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.C(n_64),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_81),
.C(n_9),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_8),
.Y(n_256)
);


endmodule