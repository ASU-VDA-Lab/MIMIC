module fake_jpeg_30387_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_23),
.B(n_13),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_1),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_15),
.B1(n_33),
.B2(n_32),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_37),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_14),
.B1(n_31),
.B2(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_2),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_54),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_58),
.B1(n_62),
.B2(n_40),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_43),
.B1(n_39),
.B2(n_41),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_43),
.B1(n_39),
.B2(n_41),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_42),
.B1(n_36),
.B2(n_35),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_40),
.B(n_4),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_46),
.C(n_35),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_6),
.C(n_7),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_77),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_73),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_79),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_4),
.B(n_5),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_19),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_18),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_82),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_7),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_8),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_9),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_10),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_75),
.B(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_100),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_70),
.B(n_26),
.C(n_27),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_89),
.B1(n_85),
.B2(n_88),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_88),
.C(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_101),
.Y(n_106)
);

OAI321xp33_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.A3(n_104),
.B1(n_105),
.B2(n_89),
.C(n_99),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_86),
.B(n_29),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_87),
.Y(n_112)
);


endmodule