module fake_jpeg_27075_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_17),
.Y(n_52)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_32),
.B1(n_27),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_92)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_64),
.Y(n_87)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_27),
.B1(n_30),
.B2(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_72),
.Y(n_113)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_45),
.B1(n_46),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_53),
.B1(n_50),
.B2(n_51),
.Y(n_108)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_45),
.B1(n_48),
.B2(n_32),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_78),
.A2(n_51),
.B1(n_55),
.B2(n_61),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_26),
.B(n_33),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_94),
.B(n_33),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_82),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_30),
.B1(n_21),
.B2(n_32),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_85),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_43),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_75),
.C(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_22),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_86),
.A2(n_92),
.B1(n_26),
.B2(n_34),
.Y(n_126)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_89),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_93),
.Y(n_128)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_31),
.B(n_36),
.C(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_57),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_99),
.Y(n_103)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_104),
.B(n_96),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_105),
.B(n_112),
.Y(n_152)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_109),
.B1(n_100),
.B2(n_99),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_25),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_84),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_54),
.B1(n_55),
.B2(n_61),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_76),
.B1(n_88),
.B2(n_59),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_34),
.B1(n_25),
.B2(n_35),
.Y(n_147)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_129),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_29),
.C(n_17),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_135),
.Y(n_179)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_138),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_155),
.B(n_19),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_84),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_78),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_157),
.C(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_110),
.B1(n_103),
.B2(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_143),
.B(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_78),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_106),
.A2(n_59),
.B1(n_65),
.B2(n_97),
.Y(n_145)
);

NAND2x1_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_78),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_149),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_108),
.B1(n_93),
.B2(n_102),
.Y(n_161)
);

INVx6_ASAP7_75t_SL g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_82),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_40),
.C(n_43),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_130),
.C(n_116),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_59),
.B(n_65),
.C(n_97),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_124),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_74),
.A3(n_70),
.B1(n_31),
.B2(n_36),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_152),
.A3(n_159),
.B1(n_151),
.B2(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_126),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_170),
.B(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_162),
.B1(n_174),
.B2(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_110),
.B1(n_127),
.B2(n_102),
.Y(n_162)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_163),
.A2(n_19),
.B(n_9),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_110),
.B(n_111),
.C(n_28),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_183),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_176),
.B1(n_188),
.B2(n_189),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_169),
.C(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_44),
.C(n_42),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_107),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_142),
.A2(n_114),
.B1(n_123),
.B2(n_103),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_153),
.A2(n_103),
.B1(n_123),
.B2(n_119),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_115),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_182),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_61),
.B1(n_119),
.B2(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_28),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_29),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_187),
.B(n_190),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_28),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_0),
.B(n_1),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_141),
.A2(n_130),
.B1(n_44),
.B2(n_42),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_24),
.B1(n_20),
.B2(n_18),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_194),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g195 ( 
.A1(n_160),
.A2(n_155),
.B1(n_132),
.B2(n_150),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_203),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_143),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_201),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_150),
.B(n_149),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_200),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_133),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_206),
.Y(n_237)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_177),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_210),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_133),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_162),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_0),
.B(n_1),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_131),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_164),
.B(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_219),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_24),
.B1(n_20),
.B2(n_19),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_218),
.B1(n_178),
.B2(n_187),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_170),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_161),
.A2(n_24),
.B1(n_20),
.B2(n_28),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_10),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_9),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_10),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_19),
.C(n_9),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_191),
.C(n_189),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_163),
.C(n_186),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_229),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_194),
.B(n_197),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_188),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_241),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_242),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_213),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_243),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_7),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_250),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_220),
.B(n_3),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_249),
.A2(n_224),
.B1(n_232),
.B2(n_225),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_251),
.A2(n_264),
.B1(n_246),
.B2(n_242),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_252),
.B(n_228),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_204),
.C(n_195),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_261),
.C(n_267),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_246),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_224),
.B1(n_205),
.B2(n_203),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_269),
.B1(n_270),
.B2(n_247),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_195),
.C(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_232),
.A2(n_199),
.B1(n_211),
.B2(n_208),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_197),
.C(n_208),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_198),
.B(n_202),
.C(n_216),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_225),
.A2(n_223),
.B(n_4),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_270),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_255),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_273),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_275),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_298)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_239),
.C(n_235),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_280),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_234),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_269),
.B1(n_259),
.B2(n_2),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_233),
.C(n_229),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_231),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_233),
.C(n_238),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_238),
.C(n_234),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_263),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_250),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_289),
.B(n_269),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_19),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_256),
.B1(n_264),
.B2(n_251),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_12),
.B1(n_16),
.B2(n_6),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_288),
.A2(n_255),
.B(n_258),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_4),
.B(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_292),
.Y(n_316)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_262),
.B(n_253),
.Y(n_293)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_293),
.A2(n_302),
.B(n_4),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_303),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_2),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_269),
.B1(n_281),
.B2(n_277),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_278),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_304),
.A2(n_11),
.B1(n_16),
.B2(n_5),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_274),
.C(n_277),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_305),
.B(n_312),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_314),
.B1(n_297),
.B2(n_299),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_300),
.B1(n_296),
.B2(n_304),
.Y(n_325)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_313),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_268),
.C(n_7),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_16),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_315),
.B(n_7),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_318),
.B(n_322),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_290),
.B1(n_296),
.B2(n_295),
.Y(n_320)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_298),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_294),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_323),
.A2(n_314),
.B(n_306),
.Y(n_326)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_313),
.C(n_293),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_293),
.C(n_294),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_307),
.C(n_11),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_332),
.A2(n_317),
.B1(n_324),
.B2(n_14),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_328),
.C(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_333),
.C(n_329),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_334),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_12),
.C(n_14),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_14),
.C(n_15),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_4),
.Y(n_342)
);


endmodule