module fake_jpeg_26156_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_8),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_21),
.Y(n_43)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_67),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_68),
.Y(n_91)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_69),
.B1(n_36),
.B2(n_43),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_63),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_32),
.Y(n_63)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_33),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_26),
.B1(n_23),
.B2(n_32),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_45),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_102),
.C(n_45),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_54),
.B1(n_30),
.B2(n_72),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_26),
.B1(n_39),
.B2(n_22),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_76),
.A2(n_101),
.B1(n_82),
.B2(n_79),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_80),
.Y(n_137)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_39),
.B1(n_46),
.B2(n_44),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_108),
.B1(n_45),
.B2(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_83),
.B(n_87),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_39),
.B1(n_43),
.B2(n_40),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_86),
.B1(n_40),
.B2(n_29),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_58),
.B1(n_73),
.B2(n_68),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_44),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_98),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_42),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_103),
.B(n_45),
.C(n_40),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_51),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_39),
.B1(n_25),
.B2(n_22),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_28),
.B(n_31),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_42),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_18),
.B1(n_28),
.B2(n_31),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_55),
.A2(n_31),
.B1(n_28),
.B2(n_39),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_65),
.A2(n_45),
.B(n_44),
.C(n_36),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_111),
.A2(n_112),
.B(n_123),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_42),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_120),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_128),
.B1(n_89),
.B2(n_108),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_71),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_124),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_24),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_106),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_134),
.Y(n_147)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_109),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_75),
.A2(n_53),
.B1(n_54),
.B2(n_72),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_138),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_72),
.B1(n_52),
.B2(n_66),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_93),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_56),
.B1(n_62),
.B2(n_30),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_33),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_95),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_94),
.A2(n_56),
.B1(n_62),
.B2(n_33),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_99),
.B1(n_110),
.B2(n_82),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_145),
.B(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_108),
.B1(n_74),
.B2(n_81),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_144),
.B1(n_151),
.B2(n_119),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_123),
.A2(n_81),
.B1(n_78),
.B2(n_107),
.Y(n_144)
);

XOR2x2_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_103),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_78),
.B1(n_90),
.B2(n_87),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_152),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_103),
.C(n_77),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_160),
.C(n_112),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_93),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_114),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_92),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_111),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_98),
.B(n_83),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_170),
.B(n_33),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_99),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_172),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_124),
.B(n_111),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_125),
.B(n_129),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_173),
.A2(n_177),
.B(n_190),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_147),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_187),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_112),
.B(n_128),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_156),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_183),
.B1(n_201),
.B2(n_164),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_115),
.B1(n_121),
.B2(n_89),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_192),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_2),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_140),
.A2(n_89),
.B1(n_22),
.B2(n_34),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_143),
.B1(n_157),
.B2(n_170),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_3),
.B(n_4),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_3),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_191),
.A2(n_199),
.B(n_3),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_33),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_196),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_109),
.C(n_34),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_153),
.C(n_141),
.Y(n_217)
);

BUFx12f_ASAP7_75t_SL g199 ( 
.A(n_167),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_177),
.B(n_190),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_35),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_143),
.Y(n_216)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_158),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_223),
.B(n_224),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_229),
.B1(n_202),
.B2(n_205),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_186),
.B1(n_161),
.B2(n_188),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_211),
.B1(n_214),
.B2(n_218),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_165),
.B1(n_151),
.B2(n_152),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_213),
.C(n_217),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_160),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_219),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_150),
.B1(n_34),
.B2(n_25),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_150),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_109),
.C(n_25),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_230),
.C(n_198),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_197),
.B(n_196),
.C(n_201),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_181),
.B(n_35),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_195),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_21),
.B(n_24),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_176),
.A2(n_21),
.B1(n_24),
.B2(n_5),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_6),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_203),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_187),
.B(n_191),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_180),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_4),
.Y(n_230)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_7),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_235),
.B(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_192),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_241),
.B1(n_245),
.B2(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_204),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_247),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_246),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_175),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_250),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_226),
.B1(n_182),
.B2(n_210),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_197),
.Y(n_266)
);

NAND2x1_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_182),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_207),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_218),
.B1(n_223),
.B2(n_228),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_258),
.B1(n_259),
.B2(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_213),
.C(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_257),
.C(n_260),
.Y(n_275)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_220),
.C(n_230),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_252),
.B1(n_247),
.B2(n_240),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_215),
.C(n_196),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_267),
.Y(n_279)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_197),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_7),
.C(n_8),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_249),
.C(n_245),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_238),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_278),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_269),
.B1(n_239),
.B2(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_282),
.C(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_9),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_236),
.C(n_243),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_284),
.C(n_275),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_239),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_283),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_232),
.C(n_239),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_267),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_287),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_263),
.Y(n_287)
);

OR2x2_ASAP7_75t_SL g290 ( 
.A(n_273),
.B(n_259),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_15),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_294),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_261),
.B(n_268),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_295),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_249),
.C(n_10),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_296),
.B(n_9),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_281),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_302),
.B(n_11),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_279),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_9),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_10),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_291),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_287),
.C(n_295),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_311),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_286),
.C(n_290),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_309),
.A2(n_297),
.B(n_302),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_314),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_306),
.B1(n_299),
.B2(n_15),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_316),
.B(n_315),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_315),
.B1(n_13),
.B2(n_14),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_14),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_320),
.Y(n_321)
);


endmodule