module fake_jpeg_12573_n_575 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_575);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_575;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_5),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_54),
.B(n_75),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_65),
.B(n_66),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_31),
.A2(n_17),
.B(n_16),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g159 ( 
.A(n_72),
.B(n_90),
.CON(n_159),
.SN(n_159)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_77),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_17),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_16),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_25),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_85),
.Y(n_126)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

HAxp5_ASAP7_75t_SL g90 ( 
.A(n_36),
.B(n_0),
.CON(n_90),
.SN(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_101),
.Y(n_150)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_106),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_25),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_36),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_36),
.B(n_0),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_25),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_77),
.B(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_132),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_36),
.B1(n_26),
.B2(n_32),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_112),
.A2(n_162),
.B1(n_95),
.B2(n_94),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_23),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_119),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_63),
.B(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_124),
.B(n_127),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_53),
.A2(n_32),
.B1(n_48),
.B2(n_44),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_131),
.A2(n_84),
.B1(n_78),
.B2(n_73),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_51),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_133),
.B(n_138),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_58),
.B(n_38),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_61),
.B(n_35),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_155),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_55),
.B(n_50),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_55),
.B(n_27),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_35),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_76),
.A2(n_26),
.B1(n_32),
.B2(n_48),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_82),
.B(n_45),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_164),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_81),
.B(n_51),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_56),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_126),
.Y(n_184)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

CKINVDCx12_ASAP7_75t_R g174 ( 
.A(n_135),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_174),
.Y(n_255)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_176),
.B(n_182),
.Y(n_243)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_177),
.Y(n_265)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_178),
.Y(n_249)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_183),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_184),
.B(n_202),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_185),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_96),
.B1(n_98),
.B2(n_25),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_188),
.B(n_205),
.Y(n_250)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_189),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_40),
.B1(n_27),
.B2(n_28),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_190),
.Y(n_273)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_192),
.Y(n_285)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_195),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_122),
.A2(n_45),
.B1(n_28),
.B2(n_33),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_196),
.A2(n_201),
.B1(n_229),
.B2(n_118),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_197),
.Y(n_277)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_127),
.B(n_103),
.C(n_57),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_210),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_141),
.A2(n_40),
.B1(n_50),
.B2(n_34),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_136),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_34),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_0),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_134),
.B(n_113),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_206),
.Y(n_267)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_140),
.B(n_169),
.C(n_149),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_213),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_123),
.B(n_102),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_212),
.B(n_221),
.Y(n_280)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

CKINVDCx6p67_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

NAND2x1_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_230),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_162),
.A2(n_39),
.B1(n_64),
.B2(n_62),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_217),
.B1(n_161),
.B2(n_154),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_112),
.A2(n_39),
.B1(n_60),
.B2(n_91),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_152),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_218),
.B(n_219),
.Y(n_286)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_157),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_131),
.A2(n_100),
.B1(n_99),
.B2(n_59),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_232),
.B1(n_69),
.B2(n_145),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_149),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_223),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_123),
.B(n_33),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_224),
.B(n_227),
.Y(n_283)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_225),
.B(n_228),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_169),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_115),
.A2(n_90),
.B(n_1),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_232),
.A2(n_158),
.B1(n_165),
.B2(n_144),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_233),
.A2(n_221),
.B1(n_177),
.B2(n_229),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_237),
.A2(n_239),
.B1(n_252),
.B2(n_257),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_165),
.B1(n_144),
.B2(n_139),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_242),
.A2(n_263),
.B1(n_270),
.B2(n_275),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_244),
.B(n_6),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_204),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_247),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_171),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_248),
.B(n_269),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_145),
.B1(n_117),
.B2(n_120),
.Y(n_252)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_118),
.B(n_125),
.C(n_115),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_211),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_114),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_272),
.C(n_276),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_172),
.A2(n_117),
.B1(n_154),
.B2(n_129),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_193),
.A2(n_125),
.B1(n_128),
.B2(n_161),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_179),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_210),
.A2(n_139),
.B1(n_128),
.B2(n_52),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_203),
.B(n_39),
.C(n_1),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_195),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_199),
.B(n_48),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_213),
.B1(n_218),
.B2(n_225),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_250),
.B(n_181),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_289),
.B(n_315),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_206),
.C(n_191),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_297),
.C(n_334),
.Y(n_353)
);

BUFx4f_ASAP7_75t_SL g292 ( 
.A(n_255),
.Y(n_292)
);

INVx11_ASAP7_75t_L g363 ( 
.A(n_292),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_242),
.A2(n_266),
.B1(n_270),
.B2(n_273),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_293),
.A2(n_301),
.B1(n_307),
.B2(n_326),
.Y(n_369)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_294),
.Y(n_343)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_296),
.A2(n_306),
.B(n_321),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_189),
.C(n_187),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_246),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_300),
.B(n_303),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_302),
.A2(n_323),
.B1(n_300),
.B2(n_311),
.Y(n_350)
);

AND2x2_ASAP7_75t_SL g303 ( 
.A(n_256),
.B(n_219),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_304),
.B(n_305),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_254),
.B(n_207),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_266),
.A2(n_214),
.B1(n_173),
.B2(n_200),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_222),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_310),
.B(n_325),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_313),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_243),
.B(n_228),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_240),
.Y(n_316)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_316),
.Y(n_379)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_318),
.A2(n_319),
.B1(n_279),
.B2(n_287),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_214),
.Y(n_320)
);

BUFx12_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_280),
.B(n_194),
.Y(n_321)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_255),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_264),
.B(n_244),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_324),
.B(n_327),
.C(n_330),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_6),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_281),
.A2(n_214),
.B1(n_209),
.B2(n_197),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_282),
.B(n_180),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_235),
.B(n_7),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_15),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_249),
.B(n_8),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_249),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_332),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_251),
.B(n_278),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g333 ( 
.A1(n_272),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_337),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_251),
.B(n_8),
.C(n_9),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_8),
.C(n_10),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_286),
.C(n_246),
.Y(n_361)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_260),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_267),
.Y(n_337)
);

AOI22x1_ASAP7_75t_L g341 ( 
.A1(n_293),
.A2(n_239),
.B1(n_246),
.B2(n_286),
.Y(n_341)
);

OA22x2_ASAP7_75t_L g400 ( 
.A1(n_341),
.A2(n_303),
.B1(n_308),
.B2(n_290),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_262),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_344),
.A2(n_364),
.B(n_342),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_314),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_345),
.B(n_357),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_323),
.A2(n_261),
.B1(n_284),
.B2(n_265),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_377),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_311),
.A2(n_306),
.B1(n_296),
.B2(n_312),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_349),
.A2(n_352),
.B(n_358),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_350),
.A2(n_354),
.B1(n_299),
.B2(n_302),
.Y(n_397)
);

AO22x1_ASAP7_75t_L g352 ( 
.A1(n_301),
.A2(n_268),
.B1(n_259),
.B2(n_253),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_288),
.A2(n_265),
.B1(n_274),
.B2(n_268),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_292),
.B(n_278),
.Y(n_357)
);

AO22x1_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_253),
.B1(n_259),
.B2(n_279),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_307),
.A2(n_286),
.B1(n_287),
.B2(n_236),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_359),
.A2(n_380),
.B1(n_15),
.B2(n_373),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_371),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_325),
.A2(n_260),
.B(n_262),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_365),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_236),
.B(n_11),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_321),
.B(n_335),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_10),
.C(n_11),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_290),
.C(n_329),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_292),
.B(n_11),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_303),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_376),
.A2(n_334),
.B1(n_299),
.B2(n_337),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_310),
.B(n_13),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_326),
.A2(n_15),
.B1(n_318),
.B2(n_294),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_375),
.Y(n_382)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

BUFx12f_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_386),
.Y(n_437)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_375),
.Y(n_387)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_388),
.A2(n_405),
.B(n_407),
.Y(n_429)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_320),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_390),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_395),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_321),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_392),
.Y(n_420)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_394),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_297),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_397),
.A2(n_369),
.B1(n_364),
.B2(n_358),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_340),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_417),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_399),
.A2(n_415),
.B1(n_347),
.B2(n_358),
.Y(n_448)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_400),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_402),
.Y(n_428)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_333),
.Y(n_403)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_355),
.B(n_313),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_404),
.B(n_411),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_295),
.Y(n_406)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_349),
.A2(n_322),
.B(n_336),
.Y(n_407)
);

INVx13_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_408),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_353),
.B(n_317),
.C(n_309),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_416),
.C(n_361),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_319),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_412),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_376),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_351),
.B(n_360),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_414),
.B(n_419),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_366),
.B1(n_341),
.B2(n_362),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_353),
.B(n_367),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_342),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_348),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_360),
.B(n_370),
.Y(n_419)
);

NOR3xp33_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_367),
.C(n_356),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_421),
.B(n_440),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_425),
.B(n_441),
.C(n_431),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_367),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_434),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_356),
.Y(n_434)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_435),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_343),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_395),
.B(n_341),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_418),
.B(n_368),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_442),
.B(n_445),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_444),
.A2(n_453),
.B1(n_390),
.B2(n_409),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_393),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_403),
.B(n_389),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_396),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_448),
.A2(n_396),
.B1(n_391),
.B2(n_405),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_343),
.Y(n_450)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_397),
.A2(n_362),
.B1(n_352),
.B2(n_374),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_425),
.B(n_415),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_459),
.Y(n_485)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_400),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_457),
.B(n_460),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_390),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_400),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_447),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_463),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_433),
.B(n_400),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_435),
.Y(n_464)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_464),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_465),
.B(n_451),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_428),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_469),
.Y(n_506)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_423),
.Y(n_467)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_467),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_468),
.A2(n_474),
.B1(n_479),
.B2(n_438),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_427),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_392),
.C(n_390),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_473),
.C(n_429),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_451),
.Y(n_471)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_471),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_392),
.C(n_390),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_448),
.A2(n_407),
.B1(n_388),
.B2(n_417),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_475),
.A2(n_478),
.B1(n_426),
.B2(n_430),
.Y(n_498)
);

A2O1A1O1Ixp25_ASAP7_75t_L g476 ( 
.A1(n_422),
.A2(n_409),
.B(n_399),
.C(n_387),
.D(n_382),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_476),
.B(n_477),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_449),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_453),
.B1(n_441),
.B2(n_443),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_443),
.A2(n_383),
.B1(n_406),
.B2(n_412),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_423),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_481),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_473),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_454),
.B(n_422),
.C(n_420),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_487),
.C(n_491),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_420),
.C(n_429),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_490),
.B(n_503),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_438),
.C(n_446),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_492),
.A2(n_496),
.B1(n_502),
.B2(n_464),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_442),
.CI(n_426),
.CON(n_495),
.SN(n_495)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_480),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_474),
.A2(n_383),
.B1(n_437),
.B2(n_424),
.Y(n_496)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_498),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_478),
.A2(n_452),
.B1(n_430),
.B2(n_437),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_499),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_452),
.C(n_424),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_500),
.B(n_487),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_468),
.A2(n_402),
.B1(n_352),
.B2(n_339),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_459),
.B(n_408),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_475),
.A2(n_385),
.B1(n_339),
.B2(n_381),
.Y(n_504)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_504),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_514),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_518),
.Y(n_531)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_512),
.A2(n_515),
.B1(n_516),
.B2(n_519),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_513),
.A2(n_501),
.B(n_486),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_479),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_492),
.A2(n_458),
.B1(n_456),
.B2(n_471),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_488),
.B(n_472),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

OAI21xp33_ASAP7_75t_SL g520 ( 
.A1(n_497),
.A2(n_482),
.B(n_476),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_513),
.Y(n_536)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_521),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_483),
.B(n_481),
.Y(n_523)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_523),
.Y(n_535)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_525),
.Y(n_530)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_505),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_510),
.A2(n_496),
.B1(n_502),
.B2(n_489),
.Y(n_527)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_527),
.Y(n_544)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_529),
.A2(n_509),
.B(n_514),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_500),
.C(n_490),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_533),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_517),
.B(n_485),
.C(n_484),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_523),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_534),
.B(n_538),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_536),
.B(n_522),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_491),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_522),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_516),
.B(n_498),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_510),
.A2(n_482),
.B1(n_495),
.B2(n_467),
.Y(n_539)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_539),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_511),
.A2(n_495),
.B1(n_504),
.B2(n_503),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_540),
.B(n_386),
.C(n_339),
.Y(n_550)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_542),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_515),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_543),
.B(n_550),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_509),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_545),
.B(n_547),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_541),
.B(n_521),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_549),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_529),
.A2(n_385),
.B1(n_381),
.B2(n_346),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_551),
.A2(n_527),
.B1(n_539),
.B2(n_528),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_553),
.B(n_536),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_557),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_533),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_558),
.B(n_561),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_526),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_532),
.C(n_542),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_563),
.A2(n_560),
.B(n_543),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_561),
.B(n_526),
.Y(n_565)
);

AOI321xp33_ASAP7_75t_SL g567 ( 
.A1(n_565),
.A2(n_555),
.A3(n_548),
.B1(n_537),
.B2(n_552),
.C(n_554),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_566),
.B(n_567),
.C(n_530),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_562),
.A2(n_544),
.B(n_558),
.Y(n_568)
);

AOI322xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_562),
.A3(n_564),
.B1(n_386),
.B2(n_530),
.C1(n_555),
.C2(n_385),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_569),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_570),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_572),
.B(n_346),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_394),
.C(n_408),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_574),
.B(n_394),
.Y(n_575)
);


endmodule