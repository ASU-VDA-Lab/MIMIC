module fake_ibex_1343_n_342 (n_85, n_84, n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_342);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_342;

wire n_151;
wire n_171;
wire n_103;
wire n_204;
wire n_274;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_124;
wire n_256;
wire n_193;
wire n_108;
wire n_165;
wire n_255;
wire n_175;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_239;
wire n_134;
wire n_94;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_176;
wire n_216;
wire n_166;
wire n_163;
wire n_114;
wire n_236;
wire n_189;
wire n_280;
wire n_317;
wire n_340;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_144;
wire n_170;
wire n_270;
wire n_113;
wire n_117;
wire n_265;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_210;
wire n_220;
wire n_287;
wire n_243;
wire n_228;
wire n_147;
wire n_251;
wire n_244;
wire n_310;
wire n_323;
wire n_143;
wire n_106;
wire n_224;
wire n_183;
wire n_333;
wire n_110;
wire n_306;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_109;
wire n_127;
wire n_121;
wire n_325;
wire n_301;
wire n_296;
wire n_120;
wire n_168;
wire n_155;
wire n_315;
wire n_122;
wire n_116;
wire n_289;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_235;
wire n_136;
wire n_261;
wire n_221;
wire n_102;
wire n_99;
wire n_269;
wire n_156;
wire n_126;
wire n_104;
wire n_141;
wire n_222;
wire n_186;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_290;
wire n_174;
wire n_157;
wire n_219;
wire n_246;
wire n_146;
wire n_207;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_205;
wire n_139;
wire n_275;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_335;
wire n_263;
wire n_299;
wire n_262;
wire n_137;
wire n_338;
wire n_173;
wire n_180;
wire n_201;
wire n_257;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_179;
wire n_100;
wire n_206;
wire n_329;
wire n_188;
wire n_200;
wire n_199;
wire n_308;
wire n_135;
wire n_283;
wire n_111;
wire n_322;
wire n_227;
wire n_115;
wire n_248;
wire n_101;
wire n_190;
wire n_138;
wire n_214;
wire n_238;
wire n_332;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_225;
wire n_272;
wire n_223;
wire n_95;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_148;
wire n_233;
wire n_118;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_178;
wire n_303;
wire n_162;
wire n_240;
wire n_282;
wire n_266;
wire n_294;
wire n_112;
wire n_284;
wire n_172;
wire n_250;
wire n_313;
wire n_119;
wire n_319;
wire n_195;
wire n_212;
wire n_311;
wire n_97;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_302;
wire n_297;
wire n_252;
wire n_107;
wire n_149;
wire n_254;
wire n_213;
wire n_271;
wire n_241;
wire n_292;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_160;
wire n_184;
wire n_232;
wire n_281;

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_48),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_91),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_18),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_12),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_33),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_45),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_16),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_7),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g128 ( 
.A(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_26),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_53),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_42),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_1),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_19),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_43),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_27),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_38),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

INVxp33_ASAP7_75t_SL g146 ( 
.A(n_52),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_22),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_14),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_31),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_13),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_3),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_69),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_51),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_20),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_72),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_0),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_46),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_21),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_28),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_2),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_111),
.B(n_9),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_10),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_15),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_17),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_98),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_102),
.B(n_90),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_127),
.B(n_32),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_147),
.B(n_47),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_113),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

AND2x4_ASAP7_75t_L g212 ( 
.A(n_107),
.B(n_55),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_106),
.A2(n_68),
.B1(n_76),
.B2(n_89),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_141),
.B(n_156),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_146),
.B1(n_167),
.B2(n_131),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_156),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_110),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_124),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_125),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_130),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_153),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_135),
.B(n_152),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_120),
.A2(n_128),
.B1(n_144),
.B2(n_141),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_94),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_128),
.A2(n_178),
.B1(n_176),
.B2(n_174),
.Y(n_234)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

NAND2xp33_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_96),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

BUFx6f_ASAP7_75t_SL g240 ( 
.A(n_181),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_144),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

NAND2x1p5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_161),
.Y(n_246)
);

OAI221xp5_ASAP7_75t_L g247 ( 
.A1(n_182),
.A2(n_172),
.B1(n_171),
.B2(n_170),
.C(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

AO22x2_ASAP7_75t_L g250 ( 
.A1(n_201),
.A2(n_154),
.B1(n_169),
.B2(n_168),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g252 ( 
.A1(n_190),
.A2(n_150),
.B1(n_165),
.B2(n_163),
.C(n_139),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_149),
.B1(n_159),
.B2(n_148),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_109),
.Y(n_254)
);

AO22x2_ASAP7_75t_L g255 ( 
.A1(n_185),
.A2(n_145),
.B1(n_143),
.B2(n_122),
.Y(n_255)
);

OAI221xp5_ASAP7_75t_L g256 ( 
.A1(n_193),
.A2(n_119),
.B1(n_157),
.B2(n_158),
.C(n_160),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_227),
.Y(n_260)
);

AO22x2_ASAP7_75t_L g261 ( 
.A1(n_194),
.A2(n_206),
.B1(n_198),
.B2(n_205),
.Y(n_261)
);

AO22x2_ASAP7_75t_L g262 ( 
.A1(n_194),
.A2(n_206),
.B1(n_208),
.B2(n_214),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_215),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_210),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_217),
.B1(n_224),
.B2(n_230),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

OAI221xp5_ASAP7_75t_L g270 ( 
.A1(n_203),
.A2(n_211),
.B1(n_228),
.B2(n_222),
.C(n_219),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_231),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_200),
.B(n_212),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_195),
.Y(n_274)
);

OAI221xp5_ASAP7_75t_L g275 ( 
.A1(n_191),
.A2(n_213),
.B1(n_187),
.B2(n_183),
.C(n_180),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_189),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

AO22x2_ASAP7_75t_L g279 ( 
.A1(n_201),
.A2(n_232),
.B1(n_185),
.B2(n_181),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_201),
.A2(n_232),
.B1(n_185),
.B2(n_181),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_242),
.Y(n_281)
);

NAND2x1p5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_277),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_241),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_260),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_236),
.A2(n_238),
.B1(n_253),
.B2(n_255),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_245),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_254),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_263),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_270),
.A2(n_268),
.B1(n_275),
.B2(n_247),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_280),
.B1(n_252),
.B2(n_250),
.Y(n_293)
);

OR2x6_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_253),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_261),
.A2(n_262),
.B1(n_255),
.B2(n_266),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_251),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_271),
.B(n_265),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_282),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_280),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_279),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_258),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_256),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_237),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_276),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_300),
.A2(n_278),
.B(n_240),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_297),
.Y(n_310)
);

O2A1O1Ixp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_289),
.B(n_298),
.C(n_296),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_285),
.Y(n_312)
);

OR2x6_ASAP7_75t_SL g313 ( 
.A(n_290),
.B(n_293),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_292),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

AND2x2_ASAP7_75t_SL g318 ( 
.A(n_312),
.B(n_295),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_311),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_303),
.A2(n_310),
.B(n_301),
.C(n_304),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_319),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_316),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_325),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_326),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_328),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_331),
.B(n_330),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

OAI221xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_327),
.B1(n_309),
.B2(n_321),
.C(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_313),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_307),
.B(n_334),
.C(n_330),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_305),
.B(n_322),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);


endmodule