module real_aes_2488_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_294;
wire n_393;
wire n_258;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_0), .A2(n_110), .B1(n_414), .B2(n_415), .Y(n_601) );
AOI222xp33_ASAP7_75t_L g381 ( .A1(n_1), .A2(n_105), .B1(n_126), .B2(n_382), .C1(n_383), .C2(n_385), .Y(n_381) );
OAI22x1_ASAP7_75t_L g312 ( .A1(n_2), .A2(n_313), .B1(n_314), .B2(n_353), .Y(n_312) );
INVx1_ASAP7_75t_L g353 ( .A(n_2), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_3), .A2(n_99), .B1(n_281), .B2(n_378), .Y(n_377) );
AO22x2_ASAP7_75t_L g233 ( .A1(n_4), .A2(n_147), .B1(n_230), .B2(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g618 ( .A(n_4), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_5), .A2(n_13), .B1(n_281), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_6), .A2(n_135), .B1(n_279), .B2(n_281), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_7), .A2(n_53), .B1(n_352), .B2(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_8), .A2(n_115), .B1(n_286), .B2(n_376), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_9), .A2(n_102), .B1(n_421), .B2(n_425), .Y(n_488) );
AOI22x1_ASAP7_75t_L g420 ( .A1(n_10), .A2(n_93), .B1(n_421), .B2(n_422), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_11), .A2(n_180), .B1(n_414), .B2(n_415), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_12), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_14), .B(n_530), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_15), .A2(n_91), .B1(n_301), .B2(n_304), .Y(n_300) );
AO22x2_ASAP7_75t_L g229 ( .A1(n_16), .A2(n_50), .B1(n_230), .B2(n_231), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_16), .B(n_617), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_17), .A2(n_191), .B1(n_268), .B2(n_372), .Y(n_371) );
AO222x2_ASAP7_75t_L g626 ( .A1(n_18), .A2(n_49), .B1(n_165), .B2(n_397), .C1(n_407), .C2(n_410), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_19), .A2(n_166), .B1(n_414), .B2(n_415), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_20), .A2(n_65), .B1(n_350), .B2(n_352), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_21), .A2(n_151), .B1(n_226), .B2(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_22), .A2(n_193), .B1(n_424), .B2(n_492), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_23), .A2(n_113), .B1(n_410), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_SL g326 ( .A1(n_24), .A2(n_106), .B1(n_306), .B2(n_327), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_25), .A2(n_168), .B1(n_286), .B2(n_290), .Y(n_285) );
XNOR2xp5_ASAP7_75t_L g391 ( .A(n_26), .B(n_392), .Y(n_391) );
AOI222xp33_ASAP7_75t_L g518 ( .A1(n_27), .A2(n_45), .B1(n_120), .B2(n_397), .C1(n_478), .C2(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g531 ( .A(n_28), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_29), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_30), .A2(n_176), .B1(n_400), .B2(n_403), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_31), .A2(n_152), .B1(n_365), .B2(n_366), .Y(n_364) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_32), .A2(n_127), .B1(n_179), .B2(n_342), .C1(n_383), .C2(n_446), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_33), .A2(n_92), .B1(n_421), .B2(n_425), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_34), .A2(n_183), .B1(n_299), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_SL g405 ( .A1(n_35), .A2(n_195), .B1(n_406), .B2(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_36), .B(n_261), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_37), .A2(n_81), .B1(n_417), .B2(n_418), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_38), .A2(n_141), .B1(n_407), .B2(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_39), .A2(n_88), .B1(n_329), .B2(n_330), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_40), .A2(n_100), .B1(n_443), .B2(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_41), .A2(n_83), .B1(n_409), .B2(n_483), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_42), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_43), .A2(n_201), .B1(n_249), .B2(n_346), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_44), .A2(n_60), .B1(n_345), .B2(n_347), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_46), .A2(n_177), .B1(n_346), .B2(n_505), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_47), .A2(n_134), .B1(n_318), .B2(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_48), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_51), .A2(n_79), .B1(n_409), .B2(n_410), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_52), .A2(n_104), .B1(n_365), .B2(n_366), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_54), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_55), .A2(n_131), .B1(n_421), .B2(n_424), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_56), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g635 ( .A1(n_57), .A2(n_184), .B1(n_418), .B2(n_492), .Y(n_635) );
OAI22x1_ASAP7_75t_L g501 ( .A1(n_58), .A2(n_502), .B1(n_520), .B2(n_521), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_58), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_59), .A2(n_94), .B1(n_409), .B2(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g230 ( .A(n_61), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_62), .A2(n_122), .B1(n_425), .B2(n_606), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_63), .A2(n_125), .B1(n_268), .B2(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_64), .A2(n_143), .B1(n_295), .B2(n_298), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_66), .A2(n_148), .B1(n_366), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_67), .A2(n_85), .B1(n_375), .B2(n_376), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_68), .A2(n_96), .B1(n_268), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_69), .A2(n_98), .B1(n_418), .B2(n_606), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_70), .A2(n_136), .B1(n_346), .B2(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_71), .Y(n_339) );
INVx1_ASAP7_75t_L g470 ( .A(n_72), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_73), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_74), .A2(n_137), .B1(n_415), .B2(n_487), .Y(n_486) );
INVx1_ASAP7_75t_SL g238 ( .A(n_75), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_75), .B(n_103), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_76), .A2(n_129), .B1(n_283), .B2(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_77), .Y(n_398) );
INVx2_ASAP7_75t_L g214 ( .A(n_78), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_80), .A2(n_140), .B1(n_327), .B2(n_376), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_82), .A2(n_175), .B1(n_436), .B2(n_577), .Y(n_576) );
OA22x2_ASAP7_75t_L g221 ( .A1(n_84), .A2(n_222), .B1(n_307), .B2(n_308), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_84), .Y(n_307) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_86), .A2(n_202), .B1(n_439), .B2(n_552), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_87), .A2(n_145), .B1(n_295), .B2(n_331), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g337 ( .A(n_89), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_90), .A2(n_108), .B1(n_439), .B2(n_440), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_95), .Y(n_608) );
OA22x2_ASAP7_75t_L g524 ( .A1(n_97), .A2(n_525), .B1(n_526), .B2(n_559), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_97), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_101), .A2(n_206), .B1(n_406), .B2(n_508), .Y(n_507) );
AO22x2_ASAP7_75t_L g241 ( .A1(n_103), .A2(n_157), .B1(n_230), .B2(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_107), .A2(n_159), .B1(n_298), .B2(n_368), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_109), .A2(n_121), .B1(n_346), .B2(n_452), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g320 ( .A1(n_111), .A2(n_170), .B1(n_321), .B2(n_324), .Y(n_320) );
AOI22xp33_ASAP7_75t_SL g317 ( .A1(n_112), .A2(n_132), .B1(n_318), .B2(n_319), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_114), .A2(n_124), .B1(n_249), .B2(n_255), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_116), .A2(n_181), .B1(n_286), .B2(n_366), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_117), .A2(n_164), .B1(n_268), .B2(n_272), .Y(n_267) );
INVx1_ASAP7_75t_L g239 ( .A(n_118), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_119), .A2(n_172), .B1(n_400), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_123), .A2(n_161), .B1(n_436), .B2(n_437), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_128), .A2(n_155), .B1(n_443), .B2(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_130), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_133), .B(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_138), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_139), .A2(n_173), .B1(n_422), .B2(n_603), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_142), .A2(n_154), .B1(n_226), .B2(n_243), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_144), .A2(n_162), .B1(n_406), .B2(n_407), .Y(n_598) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_146), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_149), .A2(n_171), .B1(n_249), .B2(n_346), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_150), .A2(n_167), .B1(n_424), .B2(n_425), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_153), .A2(n_208), .B(n_215), .C(n_620), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_156), .A2(n_624), .B1(n_643), .B2(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_156), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_158), .A2(n_204), .B1(n_552), .B2(n_553), .C(n_555), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_160), .A2(n_200), .B1(n_400), .B2(n_403), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_163), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g614 ( .A(n_163), .Y(n_614) );
INVx1_ASAP7_75t_L g211 ( .A(n_169), .Y(n_211) );
AND2x2_ASAP7_75t_R g639 ( .A(n_169), .B(n_614), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_174), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_178), .A2(n_197), .B1(n_351), .B2(n_372), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_182), .A2(n_198), .B1(n_226), .B2(n_342), .Y(n_567) );
OA22x2_ASAP7_75t_L g360 ( .A1(n_185), .A2(n_361), .B1(n_362), .B2(n_386), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_185), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_186), .B(n_213), .Y(n_212) );
AO22x2_ASAP7_75t_L g431 ( .A1(n_187), .A2(n_432), .B1(n_453), .B2(n_454), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_187), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_188), .B(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_189), .A2(n_203), .B1(n_346), .B2(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_190), .A2(n_205), .B1(n_417), .B2(n_418), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_192), .B(n_397), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_194), .A2(n_622), .B1(n_623), .B2(n_637), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_194), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_196), .Y(n_532) );
XNOR2x1_ASAP7_75t_L g561 ( .A(n_199), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_209), .B(n_212), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g648 ( .A(n_210), .B(n_212), .Y(n_648) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_211), .B(n_614), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_496), .B1(n_609), .B2(n_610), .C(n_611), .Y(n_215) );
INVx1_ASAP7_75t_L g610 ( .A(n_216), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B1(n_355), .B2(n_356), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_310), .B1(n_311), .B2(n_354), .Y(n_218) );
INVx1_ASAP7_75t_SL g354 ( .A(n_219), .Y(n_354) );
BUFx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_276), .Y(n_222) );
NOR3xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_259), .C(n_266), .Y(n_223) );
NOR4xp25_ASAP7_75t_L g308 ( .A(n_224), .B(n_277), .C(n_293), .D(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_248), .Y(n_224) );
BUFx5_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
BUFx3_ASAP7_75t_L g336 ( .A(n_227), .Y(n_336) );
INVx2_ASAP7_75t_L g384 ( .A(n_227), .Y(n_384) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_235), .Y(n_227) );
AND2x4_ASAP7_75t_L g269 ( .A(n_228), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g306 ( .A(n_228), .B(n_289), .Y(n_306) );
AND2x4_ASAP7_75t_L g400 ( .A(n_228), .B(n_235), .Y(n_400) );
AND2x2_ASAP7_75t_L g406 ( .A(n_228), .B(n_270), .Y(n_406) );
AND2x2_ASAP7_75t_L g483 ( .A(n_228), .B(n_270), .Y(n_483) );
AND2x2_ASAP7_75t_L g492 ( .A(n_228), .B(n_289), .Y(n_492) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_232), .Y(n_228) );
AND2x2_ASAP7_75t_L g246 ( .A(n_229), .B(n_233), .Y(n_246) );
INVx1_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g265 ( .A(n_229), .Y(n_265) );
INVx2_ASAP7_75t_L g231 ( .A(n_230), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_230), .Y(n_234) );
OAI22x1_ASAP7_75t_L g236 ( .A1(n_230), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_230), .Y(n_237) );
INVx1_ASAP7_75t_L g242 ( .A(n_230), .Y(n_242) );
AND2x4_ASAP7_75t_L g264 ( .A(n_232), .B(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g275 ( .A(n_232), .Y(n_275) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g258 ( .A(n_233), .B(n_254), .Y(n_258) );
AND2x2_ASAP7_75t_L g257 ( .A(n_235), .B(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g297 ( .A(n_235), .B(n_264), .Y(n_297) );
AND2x4_ASAP7_75t_L g409 ( .A(n_235), .B(n_258), .Y(n_409) );
AND2x2_ASAP7_75t_L g417 ( .A(n_235), .B(n_264), .Y(n_417) );
AND2x2_ASAP7_75t_L g606 ( .A(n_235), .B(n_264), .Y(n_606) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_236), .Y(n_247) );
AND2x2_ASAP7_75t_L g251 ( .A(n_236), .B(n_241), .Y(n_251) );
INVx2_ASAP7_75t_L g271 ( .A(n_236), .Y(n_271) );
AND2x4_ASAP7_75t_L g289 ( .A(n_240), .B(n_271), .Y(n_289) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g270 ( .A(n_241), .B(n_271), .Y(n_270) );
BUFx2_ASAP7_75t_L g284 ( .A(n_241), .Y(n_284) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g450 ( .A(n_244), .Y(n_450) );
INVx3_ASAP7_75t_L g534 ( .A(n_244), .Y(n_534) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx12f_ASAP7_75t_L g342 ( .A(n_245), .Y(n_342) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x4_ASAP7_75t_L g283 ( .A(n_246), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g299 ( .A(n_246), .B(n_289), .Y(n_299) );
AND2x2_ASAP7_75t_SL g403 ( .A(n_246), .B(n_247), .Y(n_403) );
AND2x4_ASAP7_75t_L g415 ( .A(n_246), .B(n_284), .Y(n_415) );
AND2x4_ASAP7_75t_L g418 ( .A(n_246), .B(n_289), .Y(n_418) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_246), .B(n_247), .Y(n_478) );
BUFx6f_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g348 ( .A(n_250), .Y(n_348) );
BUFx4f_ASAP7_75t_L g452 ( .A(n_250), .Y(n_452) );
INVx2_ASAP7_75t_L g506 ( .A(n_250), .Y(n_506) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g263 ( .A(n_251), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g274 ( .A(n_251), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g397 ( .A(n_251), .B(n_264), .Y(n_397) );
AND2x2_ASAP7_75t_L g407 ( .A(n_251), .B(n_275), .Y(n_407) );
AND2x2_ASAP7_75t_L g410 ( .A(n_251), .B(n_252), .Y(n_410) );
AND2x2_ASAP7_75t_L g481 ( .A(n_251), .B(n_252), .Y(n_481) );
AND2x2_ASAP7_75t_L g508 ( .A(n_251), .B(n_275), .Y(n_508) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx4_ASAP7_75t_L g597 ( .A(n_256), .Y(n_597) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_257), .Y(n_346) );
AND2x2_ASAP7_75t_L g280 ( .A(n_258), .B(n_270), .Y(n_280) );
AND2x4_ASAP7_75t_L g292 ( .A(n_258), .B(n_289), .Y(n_292) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_258), .B(n_270), .Y(n_414) );
AND2x6_ASAP7_75t_L g425 ( .A(n_258), .B(n_289), .Y(n_425) );
AND2x2_ASAP7_75t_L g487 ( .A(n_258), .B(n_270), .Y(n_487) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_260), .B(n_267), .Y(n_309) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g338 ( .A(n_262), .Y(n_338) );
INVx3_ASAP7_75t_L g382 ( .A(n_262), .Y(n_382) );
INVx4_ASAP7_75t_SL g446 ( .A(n_262), .Y(n_446) );
INVx4_ASAP7_75t_SL g530 ( .A(n_262), .Y(n_530) );
INVx6_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g288 ( .A(n_264), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g303 ( .A(n_264), .B(n_270), .Y(n_303) );
AND2x6_ASAP7_75t_L g421 ( .A(n_264), .B(n_270), .Y(n_421) );
AND2x2_ASAP7_75t_L g424 ( .A(n_264), .B(n_289), .Y(n_424) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_269), .Y(n_351) );
BUFx2_ASAP7_75t_L g468 ( .A(n_269), .Y(n_468) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g352 ( .A(n_273), .Y(n_352) );
INVx2_ASAP7_75t_L g372 ( .A(n_273), .Y(n_372) );
INVx1_ASAP7_75t_L g448 ( .A(n_273), .Y(n_448) );
INVx2_ASAP7_75t_SL g571 ( .A(n_273), .Y(n_571) );
INVx6_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_293), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_285), .Y(n_277) );
BUFx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g323 ( .A(n_280), .Y(n_323) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_280), .Y(n_443) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g324 ( .A(n_282), .Y(n_324) );
INVx2_ASAP7_75t_L g463 ( .A(n_282), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_282), .A2(n_540), .B1(n_541), .B2(n_544), .Y(n_539) );
INVx5_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g511 ( .A(n_283), .Y(n_511) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g318 ( .A(n_287), .Y(n_318) );
INVx2_ASAP7_75t_SL g375 ( .A(n_287), .Y(n_375) );
INVx4_ASAP7_75t_L g548 ( .A(n_287), .Y(n_548) );
INVx3_ASAP7_75t_SL g603 ( .A(n_287), .Y(n_603) );
INVx8_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g319 ( .A(n_291), .Y(n_319) );
INVx2_ASAP7_75t_L g376 ( .A(n_291), .Y(n_376) );
INVx1_ASAP7_75t_SL g437 ( .A(n_291), .Y(n_437) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_291), .Y(n_558) );
INVx2_ASAP7_75t_SL g577 ( .A(n_291), .Y(n_577) );
INVx8_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_300), .Y(n_293) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_SL g329 ( .A(n_296), .Y(n_329) );
INVx3_ASAP7_75t_L g368 ( .A(n_296), .Y(n_368) );
INVx2_ASAP7_75t_L g439 ( .A(n_296), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_296), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_555) );
INVx6_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g515 ( .A(n_297), .Y(n_515) );
BUFx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
INVx2_ASAP7_75t_L g441 ( .A(n_299), .Y(n_441) );
BUFx2_ASAP7_75t_SL g552 ( .A(n_299), .Y(n_552) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
INVx2_ASAP7_75t_SL g436 ( .A(n_302), .Y(n_436) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g327 ( .A(n_303), .Y(n_327) );
BUFx2_ASAP7_75t_L g554 ( .A(n_303), .Y(n_554) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g366 ( .A(n_306), .Y(n_366) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_306), .Y(n_422) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_306), .Y(n_517) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_332), .Y(n_314) );
NOR2x1_ASAP7_75t_L g315 ( .A(n_316), .B(n_325), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .Y(n_316) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g380 ( .A(n_323), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2x1_ASAP7_75t_L g332 ( .A(n_333), .B(n_343), .Y(n_332) );
OAI222xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_337), .B1(n_338), .B2(n_339), .C1(n_340), .C2(n_341), .Y(n_333) );
OAI221xp5_ASAP7_75t_L g528 ( .A1(n_334), .A2(n_529), .B1(n_531), .B2(n_532), .C(n_533), .Y(n_528) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx3_ASAP7_75t_L g385 ( .A(n_342), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_349), .Y(n_343) );
BUFx6f_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_427), .B1(n_494), .B2(n_495), .Y(n_356) );
INVx1_ASAP7_75t_L g494 ( .A(n_357), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_359), .B1(n_387), .B2(n_426), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g386 ( .A(n_362), .Y(n_386) );
NAND4xp75_ASAP7_75t_L g362 ( .A(n_363), .B(n_369), .C(n_373), .D(n_381), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_377), .Y(n_373) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g543 ( .A(n_380), .Y(n_543) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_390), .Y(n_426) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_393), .B(n_411), .Y(n_392) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_394), .B(n_404), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_398), .B2(n_399), .C1(n_401), .C2(n_402), .Y(n_394) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_400), .Y(n_519) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
NOR2x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_419), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_423), .Y(n_419) );
INVx2_ASAP7_75t_L g550 ( .A(n_422), .Y(n_550) );
INVx1_ASAP7_75t_L g495 ( .A(n_427), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_471), .B2(n_472), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_431), .B1(n_455), .B2(n_456), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g454 ( .A(n_432), .Y(n_454) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_444), .Y(n_432) );
NAND4xp25_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .C(n_438), .D(n_442), .Y(n_433) );
INVx2_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_445), .B(n_447), .C(n_449), .D(n_451), .Y(n_444) );
INVx1_ASAP7_75t_L g565 ( .A(n_446), .Y(n_565) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
XOR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_470), .Y(n_456) );
NAND4xp75_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .C(n_465), .D(n_469), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
XOR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_493), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_479), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
NOR2x1_ASAP7_75t_L g484 ( .A(n_485), .B(n_489), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_488), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g609 ( .A(n_496), .Y(n_609) );
XNOR2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_587), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_522), .B1(n_584), .B2(n_585), .Y(n_497) );
INVx1_ASAP7_75t_L g584 ( .A(n_498), .Y(n_584) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g502 ( .A(n_503), .B(n_509), .C(n_513), .D(n_518), .Y(n_502) );
AND4x1_ASAP7_75t_L g520 ( .A(n_503), .B(n_509), .C(n_513), .D(n_518), .Y(n_520) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .Y(n_513) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g586 ( .A(n_523), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_560), .B1(n_582), .B2(n_583), .Y(n_523) );
INVx2_ASAP7_75t_L g582 ( .A(n_524), .Y(n_582) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND3x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .C(n_551), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_535), .Y(n_527) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .Y(n_538) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g575 ( .A(n_543), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_549), .B2(n_550), .Y(n_545) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_548), .Y(n_581) );
BUFx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g583 ( .A(n_560), .Y(n_583) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_572), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_566), .B(n_567), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_578), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
XOR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_608), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_591), .B(n_599), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_604), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx3_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_613), .B(n_616), .Y(n_647) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OAI222xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_638), .B1(n_640), .B2(n_644), .C1(n_645), .C2(n_648), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g643 ( .A(n_624), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_625), .B(n_630), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_634), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_646), .Y(n_645) );
CKINVDCx6p67_ASAP7_75t_R g646 ( .A(n_647), .Y(n_646) );
endmodule