module fake_jpeg_237_n_680 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_6),
.B(n_19),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_61),
.Y(n_206)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_63),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g158 ( 
.A(n_64),
.Y(n_158)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_10),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_67),
.B(n_113),
.Y(n_175)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_68),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_70),
.Y(n_207)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_73),
.Y(n_203)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_79),
.Y(n_181)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_82),
.B(n_86),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_83),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_85),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_12),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_87),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_90),
.Y(n_202)
);

BUFx12f_ASAP7_75t_SL g91 ( 
.A(n_41),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_91),
.B(n_128),
.Y(n_186)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_93),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_12),
.B1(n_18),
.B2(n_17),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_94),
.A2(n_21),
.B1(n_55),
.B2(n_32),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_95),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_96),
.B(n_103),
.Y(n_192)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_27),
.B(n_8),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_108),
.Y(n_212)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_109),
.Y(n_219)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_110),
.Y(n_220)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_111),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_44),
.B(n_8),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_112),
.B(n_126),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_116),
.A2(n_119),
.B(n_50),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_21),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_43),
.Y(n_124)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_44),
.B(n_12),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_50),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_48),
.Y(n_129)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_67),
.A2(n_47),
.B(n_45),
.C(n_29),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_134),
.B(n_167),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_128),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g267 ( 
.A1(n_139),
.A2(n_147),
.B1(n_178),
.B2(n_184),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_91),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_151),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_69),
.B(n_45),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_152),
.B(n_157),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_98),
.B(n_47),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_77),
.B(n_22),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_160),
.B(n_162),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_26),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_129),
.B1(n_127),
.B2(n_120),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_66),
.B(n_42),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_166),
.B(n_169),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_113),
.B(n_42),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_61),
.A2(n_21),
.B1(n_55),
.B2(n_32),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_168),
.A2(n_170),
.B1(n_172),
.B2(n_84),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_39),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_63),
.A2(n_55),
.B1(n_32),
.B2(n_33),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_75),
.A2(n_33),
.B1(n_30),
.B2(n_42),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_117),
.B(n_39),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_177),
.B(n_182),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_105),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_64),
.B(n_30),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_100),
.B(n_31),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_183),
.B(n_211),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_124),
.A2(n_31),
.B1(n_33),
.B2(n_53),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_89),
.A2(n_53),
.B1(n_51),
.B2(n_49),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_188),
.A2(n_189),
.B1(n_194),
.B2(n_200),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_87),
.A2(n_53),
.B1(n_51),
.B2(n_49),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_64),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_199),
.A2(n_1),
.B(n_2),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_83),
.A2(n_57),
.B1(n_56),
.B2(n_28),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_83),
.B(n_93),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_104),
.B(n_57),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_214),
.B(n_225),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_114),
.A2(n_56),
.B1(n_28),
.B2(n_13),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_215),
.A2(n_218),
.B1(n_0),
.B2(n_1),
.Y(n_282)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_106),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_116),
.A2(n_28),
.B1(n_12),
.B2(n_13),
.Y(n_218)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_108),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_224),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_118),
.B(n_7),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_119),
.B(n_19),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_186),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_230),
.A2(n_298),
.B1(n_215),
.B2(n_188),
.Y(n_317)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_231),
.Y(n_355)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_232),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_234),
.Y(n_310)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_235),
.Y(n_347)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_237),
.B(n_249),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_135),
.Y(n_239)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_207),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_240),
.B(n_252),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_241),
.A2(n_264),
.B1(n_297),
.B2(n_150),
.Y(n_332)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_242),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_161),
.Y(n_243)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_161),
.Y(n_245)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_245),
.Y(n_341)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_145),
.Y(n_246)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_246),
.Y(n_343)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_247),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_205),
.B(n_65),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_85),
.C(n_88),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_250),
.B(n_296),
.C(n_155),
.Y(n_362)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_251),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_257),
.Y(n_337)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_181),
.Y(n_256)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_208),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_147),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_258),
.B(n_268),
.Y(n_340)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_213),
.Y(n_260)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_260),
.Y(n_323)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_261),
.Y(n_366)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_263),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g264 ( 
.A1(n_189),
.A2(n_178),
.B1(n_184),
.B2(n_139),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_186),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_265),
.B(n_272),
.Y(n_345)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_266),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_176),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_269),
.Y(n_365)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_213),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_270),
.B(n_271),
.Y(n_348)
);

OAI32xp33_ASAP7_75t_L g271 ( 
.A1(n_175),
.A2(n_79),
.A3(n_68),
.B1(n_99),
.B2(n_90),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_208),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_142),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_273),
.B(n_274),
.Y(n_346)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_275),
.Y(n_321)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_146),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_276),
.B(n_277),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_141),
.B(n_95),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

BUFx8_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_279),
.Y(n_315)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_210),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_280),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_192),
.B(n_5),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_281),
.B(n_283),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_282),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_328)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

AOI22x1_ASAP7_75t_SL g284 ( 
.A1(n_134),
.A2(n_222),
.B1(n_220),
.B2(n_219),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_284),
.Y(n_350)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_190),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_285),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_148),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_148),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_154),
.Y(n_288)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_143),
.Y(n_289)
);

AO22x1_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_204),
.B1(n_155),
.B2(n_202),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_153),
.A2(n_5),
.B1(n_16),
.B2(n_15),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_290),
.A2(n_307),
.B(n_200),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_158),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_293),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_156),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_181),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_294),
.A2(n_302),
.B1(n_140),
.B2(n_132),
.Y(n_333)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_143),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_299),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_197),
.B(n_0),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_168),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_149),
.A2(n_14),
.B1(n_16),
.B2(n_15),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_154),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_165),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_304),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_209),
.B(n_14),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_216),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_159),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_306),
.B(n_308),
.Y(n_364)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_202),
.Y(n_308)
);

BUFx8_ASAP7_75t_L g309 ( 
.A(n_158),
.Y(n_309)
);

NAND2x1_ASAP7_75t_SL g358 ( 
.A(n_309),
.B(n_221),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_258),
.A2(n_170),
.B1(n_172),
.B2(n_218),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_312),
.A2(n_317),
.B1(n_332),
.B2(n_335),
.Y(n_389)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_314),
.Y(n_372)
);

OAI22x1_ASAP7_75t_L g316 ( 
.A1(n_267),
.A2(n_140),
.B1(n_150),
.B2(n_203),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_316),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_262),
.B(n_248),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_322),
.B(n_327),
.C(n_352),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_324),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_254),
.B(n_179),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_333),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_233),
.A2(n_156),
.B1(n_194),
.B2(n_201),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_307),
.A2(n_191),
.B(n_180),
.C(n_171),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_336),
.B(n_245),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_284),
.A2(n_203),
.B1(n_196),
.B2(n_173),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_342),
.A2(n_353),
.B1(n_357),
.B2(n_371),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_267),
.A2(n_264),
.B(n_244),
.C(n_241),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_250),
.B(n_296),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_305),
.B(n_136),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_244),
.A2(n_230),
.B1(n_271),
.B2(n_292),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_303),
.A2(n_187),
.B1(n_173),
.B2(n_164),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_300),
.A2(n_221),
.B1(n_164),
.B2(n_158),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_358),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_309),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_297),
.A2(n_296),
.B1(n_267),
.B2(n_256),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_267),
.A2(n_202),
.B1(n_3),
.B2(n_4),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_373),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_263),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_382),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_376),
.B(n_392),
.C(n_396),
.Y(n_421)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_379),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_290),
.B1(n_259),
.B2(n_275),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_380),
.A2(n_393),
.B1(n_410),
.B2(n_411),
.Y(n_454)
);

BUFx5_ASAP7_75t_L g381 ( 
.A(n_326),
.Y(n_381)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_261),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_340),
.A2(n_324),
.B(n_316),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_383),
.A2(n_390),
.B(n_351),
.Y(n_458)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_320),
.B(n_268),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_386),
.Y(n_432)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_329),
.Y(n_387)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_387),
.Y(n_459)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_329),
.Y(n_388)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_309),
.B(n_278),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_274),
.C(n_276),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_348),
.A2(n_231),
.B1(n_286),
.B2(n_287),
.Y(n_393)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_395),
.B(n_397),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_322),
.B(n_273),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_229),
.C(n_228),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_398),
.B(n_418),
.C(n_325),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_319),
.B(n_285),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_406),
.Y(n_431)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_402),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_339),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_401),
.B(n_414),
.Y(n_443)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_404),
.B(n_407),
.Y(n_430)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g444 ( 
.A1(n_405),
.A2(n_310),
.B1(n_326),
.B2(n_365),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_319),
.B(n_260),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_331),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_412),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_348),
.A2(n_232),
.B1(n_294),
.B2(n_269),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_363),
.A2(n_243),
.B1(n_280),
.B2(n_251),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_336),
.B(n_299),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_348),
.A2(n_270),
.B1(n_239),
.B2(n_234),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_413),
.A2(n_419),
.B1(n_314),
.B2(n_334),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_283),
.Y(n_414)
);

AOI32xp33_ASAP7_75t_L g415 ( 
.A1(n_345),
.A2(n_288),
.A3(n_238),
.B1(n_308),
.B2(n_295),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_415),
.A2(n_358),
.B(n_314),
.Y(n_428)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_417),
.Y(n_446)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_340),
.B(n_289),
.C(n_236),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_350),
.A2(n_344),
.B1(n_371),
.B2(n_312),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_339),
.B(n_14),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_349),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_406),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_422),
.B(n_434),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_389),
.A2(n_335),
.B1(n_328),
.B2(n_356),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_423),
.A2(n_425),
.B1(n_428),
.B2(n_435),
.Y(n_481)
);

OAI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_424),
.A2(n_439),
.B1(n_458),
.B2(n_413),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_389),
.A2(n_333),
.B1(n_321),
.B2(n_337),
.Y(n_425)
);

OAI22x1_ASAP7_75t_L g426 ( 
.A1(n_409),
.A2(n_403),
.B1(n_372),
.B2(n_394),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_347),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_429),
.B(n_457),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_399),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_373),
.A2(n_321),
.B1(n_347),
.B2(n_313),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_378),
.A2(n_358),
.B(n_368),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_436),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_403),
.A2(n_313),
.B1(n_368),
.B2(n_343),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_437),
.A2(n_455),
.B1(n_461),
.B2(n_393),
.Y(n_483)
);

AOI22x1_ASAP7_75t_SL g439 ( 
.A1(n_419),
.A2(n_326),
.B1(n_325),
.B2(n_323),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_444),
.A2(n_310),
.B1(n_326),
.B2(n_418),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_374),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_449),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_447),
.B(n_387),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_380),
.A2(n_365),
.B1(n_338),
.B2(n_343),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_448),
.A2(n_409),
.B1(n_372),
.B2(n_411),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_391),
.A2(n_360),
.B(n_359),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_407),
.B(n_359),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_420),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_421),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_383),
.A2(n_360),
.B1(n_338),
.B2(n_351),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_390),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_456),
.B(n_449),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_375),
.B(n_323),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_404),
.A2(n_338),
.B1(n_318),
.B2(n_315),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_433),
.A2(n_408),
.B1(n_401),
.B2(n_412),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_462),
.A2(n_478),
.B1(n_489),
.B2(n_428),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_422),
.B(n_385),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_465),
.B(n_475),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_457),
.C(n_451),
.Y(n_501)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_469),
.A2(n_470),
.B1(n_483),
.B2(n_495),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_434),
.A2(n_379),
.B1(n_409),
.B2(n_376),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_471),
.Y(n_512)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_398),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_473),
.B(n_496),
.Y(n_516)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_446),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_477),
.B(n_482),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_433),
.A2(n_377),
.B1(n_384),
.B2(n_391),
.Y(n_478)
);

CKINVDCx12_ASAP7_75t_R g479 ( 
.A(n_452),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_479),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_421),
.B(n_375),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_429),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_450),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_443),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_484),
.Y(n_505)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_459),
.Y(n_485)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_485),
.Y(n_520)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_459),
.Y(n_486)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_442),
.A2(n_377),
.B1(n_410),
.B2(n_382),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_443),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_490),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_431),
.B(n_392),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_491),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_492),
.Y(n_503)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_493),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_494),
.A2(n_435),
.B1(n_430),
.B2(n_461),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_426),
.A2(n_437),
.B1(n_423),
.B2(n_425),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_431),
.B(n_402),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_497),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_498),
.A2(n_499),
.B1(n_458),
.B2(n_439),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_426),
.A2(n_388),
.B1(n_400),
.B2(n_405),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_501),
.B(n_508),
.C(n_515),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_509),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_507),
.A2(n_514),
.B1(n_518),
.B2(n_532),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_466),
.B(n_427),
.C(n_441),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_430),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_474),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_510),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_467),
.B(n_427),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_513),
.B(n_462),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_467),
.B(n_442),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_470),
.A2(n_448),
.B1(n_441),
.B2(n_453),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_438),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_522),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_523),
.A2(n_474),
.B1(n_478),
.B2(n_469),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_490),
.B(n_447),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g550 ( 
.A(n_527),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_481),
.A2(n_454),
.B1(n_424),
.B2(n_453),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_529),
.A2(n_530),
.B1(n_464),
.B2(n_482),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_481),
.A2(n_454),
.B1(n_445),
.B2(n_456),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_495),
.A2(n_439),
.B1(n_438),
.B2(n_436),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_318),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_533),
.B(n_489),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_488),
.B(n_455),
.C(n_417),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_536),
.C(n_468),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_488),
.B(n_416),
.C(n_330),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_534),
.Y(n_537)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_537),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_538),
.A2(n_546),
.B1(n_518),
.B2(n_519),
.Y(n_586)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_534),
.Y(n_541)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_541),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_542),
.B(n_530),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_557),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_471),
.C(n_472),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_544),
.B(n_562),
.C(n_563),
.Y(n_573)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_525),
.Y(n_545)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_545),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_505),
.A2(n_492),
.B(n_464),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_547),
.A2(n_554),
.B(n_541),
.Y(n_592)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_505),
.B(n_463),
.Y(n_551)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_551),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_516),
.B(n_496),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_552),
.B(n_558),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_511),
.A2(n_463),
.B(n_499),
.Y(n_554)
);

BUFx24_ASAP7_75t_SL g555 ( 
.A(n_511),
.Y(n_555)
);

BUFx24_ASAP7_75t_SL g572 ( 
.A(n_555),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_503),
.A2(n_477),
.B1(n_476),
.B2(n_483),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_556),
.A2(n_567),
.B1(n_512),
.B2(n_519),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_509),
.B(n_497),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_526),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_502),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_559),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_508),
.B(n_465),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_560),
.B(n_564),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_504),
.B(n_475),
.C(n_479),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_521),
.B(n_536),
.C(n_515),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_513),
.B(n_493),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_525),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_565),
.B(n_566),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_395),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_514),
.A2(n_487),
.B1(n_486),
.B2(n_485),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_502),
.Y(n_568)
);

AOI21xp33_ASAP7_75t_L g575 ( 
.A1(n_568),
.A2(n_569),
.B(n_512),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_524),
.B(n_452),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_574),
.B(n_542),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_575),
.B(n_583),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_540),
.B(n_535),
.C(n_517),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_580),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_561),
.A2(n_507),
.B(n_517),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_SL g581 ( 
.A(n_539),
.B(n_526),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_585),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_540),
.B(n_529),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g614 ( 
.A1(n_586),
.A2(n_311),
.B1(n_355),
.B2(n_381),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_500),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_587),
.B(n_593),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_546),
.A2(n_506),
.B1(n_510),
.B2(n_531),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_590),
.A2(n_594),
.B1(n_549),
.B2(n_545),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_551),
.A2(n_531),
.B(n_528),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_591),
.B(n_355),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_592),
.A2(n_553),
.B(n_567),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_539),
.B(n_415),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_538),
.A2(n_528),
.B1(n_520),
.B2(n_524),
.Y(n_594)
);

AOI21x1_ASAP7_75t_L g596 ( 
.A1(n_592),
.A2(n_547),
.B(n_554),
.Y(n_596)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_596),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_544),
.C(n_543),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_597),
.B(n_598),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_563),
.C(n_560),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_582),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_599),
.B(n_602),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_570),
.B(n_556),
.Y(n_600)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_600),
.Y(n_633)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_588),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_603),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_604),
.B(n_607),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_572),
.B(n_557),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_608),
.B(n_609),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_588),
.A2(n_550),
.B(n_549),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_573),
.B(n_564),
.C(n_565),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_610),
.B(n_611),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_585),
.B(n_577),
.C(n_587),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_589),
.B(n_520),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_583),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_577),
.B(n_311),
.C(n_369),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_613),
.B(n_595),
.C(n_581),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_617),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_616),
.A2(n_579),
.B1(n_584),
.B2(n_590),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_595),
.B(n_355),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_610),
.B(n_586),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_618),
.B(n_621),
.Y(n_639)
);

BUFx24_ASAP7_75t_SL g619 ( 
.A(n_601),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_619),
.B(n_366),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_598),
.B(n_576),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_622),
.B(n_623),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_624),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_597),
.B(n_611),
.C(n_605),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_625),
.B(n_626),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_606),
.B(n_571),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_605),
.B(n_574),
.C(n_594),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_635),
.B(n_369),
.Y(n_648)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_635),
.B(n_607),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_636),
.B(n_643),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_629),
.A2(n_606),
.B(n_596),
.Y(n_637)
);

AOI21x1_ASAP7_75t_L g661 ( 
.A1(n_637),
.A2(n_16),
.B(n_18),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_628),
.B(n_609),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_638),
.B(n_644),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_627),
.A2(n_603),
.B(n_600),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_640),
.A2(n_642),
.B(n_647),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_628),
.A2(n_604),
.B(n_602),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_633),
.A2(n_571),
.B1(n_612),
.B2(n_613),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_624),
.A2(n_593),
.B1(n_615),
.B2(n_617),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_634),
.B(n_615),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_648),
.B(n_650),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_630),
.A2(n_366),
.B(n_15),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g656 ( 
.A1(n_649),
.A2(n_16),
.B(n_18),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_639),
.B(n_632),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_652),
.B(n_654),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_636),
.B(n_625),
.C(n_620),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_653),
.B(n_655),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_645),
.B(n_620),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_642),
.B(n_621),
.C(n_631),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_656),
.B(n_659),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_641),
.B(n_631),
.C(n_3),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_661),
.A2(n_649),
.B(n_644),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_653),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_662),
.B(n_665),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_SL g665 ( 
.A(n_660),
.B(n_640),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_655),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_666),
.B(n_669),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_667),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_658),
.A2(n_646),
.B(n_643),
.Y(n_669)
);

A2O1A1O1Ixp25_ASAP7_75t_L g671 ( 
.A1(n_663),
.A2(n_657),
.B(n_659),
.C(n_651),
.D(n_4),
.Y(n_671)
);

AO21x1_ASAP7_75t_L g676 ( 
.A1(n_671),
.A2(n_674),
.B(n_662),
.Y(n_676)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_664),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_672),
.B(n_668),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_675),
.A2(n_676),
.B(n_670),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_677),
.A2(n_673),
.B(n_657),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_SL g679 ( 
.A1(n_678),
.A2(n_2),
.B(n_3),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_2),
.Y(n_680)
);


endmodule