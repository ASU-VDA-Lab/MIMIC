module fake_jpeg_17909_n_85 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_85);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_85;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx4f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_0),
.C(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_24),
.B1(n_16),
.B2(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_16),
.B1(n_17),
.B2(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_13),
.B1(n_10),
.B2(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_13),
.B1(n_1),
.B2(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_21),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_21),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_20),
.B(n_19),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_12),
.B1(n_15),
.B2(n_11),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.C(n_41),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_28),
.B(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_33),
.B1(n_32),
.B2(n_40),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_15),
.B(n_26),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_42),
.C(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_19),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.C(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_46),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_39),
.C(n_19),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_60),
.B1(n_47),
.B2(n_46),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_48),
.B1(n_45),
.B2(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_65),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_18),
.C(n_52),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_68),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_24),
.C(n_19),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_24),
.C(n_3),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_56),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_79),
.Y(n_81)
);

AOI31xp67_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_77),
.A3(n_74),
.B(n_72),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_5),
.B(n_6),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_81),
.B(n_7),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_7),
.Y(n_85)
);


endmodule