module fake_jpeg_19156_n_128 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_128);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_68),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_85),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_47),
.B1(n_40),
.B2(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_82),
.B1(n_53),
.B2(n_52),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_49),
.B1(n_57),
.B2(n_45),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_54),
.Y(n_94)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_83),
.C(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.Y(n_108)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_46),
.C(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_100),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_41),
.B1(n_48),
.B2(n_39),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_39),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_22),
.B(n_38),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_2),
.B(n_3),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_4),
.C(n_5),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_107),
.B(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_26),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_96),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_114),
.B(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_116),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_120),
.A2(n_108),
.B1(n_109),
.B2(n_119),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_111),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_24),
.B1(n_10),
.B2(n_12),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_27),
.C(n_15),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_28),
.B(n_19),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_31),
.Y(n_128)
);


endmodule