module fake_netlist_1_12511_n_727 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_727);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_727;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g101 ( .A(n_67), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_96), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_30), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_75), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_55), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_83), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_58), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_98), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_61), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_22), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_50), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_95), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_3), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_6), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_86), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_88), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_89), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
CKINVDCx14_ASAP7_75t_R g124 ( .A(n_76), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_11), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_99), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_44), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_59), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_43), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_69), .B(n_52), .Y(n_130) );
INVx1_ASAP7_75t_SL g131 ( .A(n_46), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_65), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_39), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_32), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_10), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_42), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_16), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_94), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_20), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_45), .Y(n_141) );
INVx1_ASAP7_75t_SL g142 ( .A(n_53), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_40), .Y(n_143) );
CKINVDCx14_ASAP7_75t_R g144 ( .A(n_64), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g145 ( .A(n_41), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_2), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_101), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_126), .A2(n_0), .B(n_1), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_109), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_143), .B(n_0), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g154 ( .A1(n_105), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_116), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_112), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_140), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_107), .B(n_4), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_104), .B(n_125), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_116), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_116), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_145), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_159), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_159), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_150), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_166), .B(n_111), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_166), .A2(n_105), .B1(n_122), .B2(n_138), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
OR2x6_ASAP7_75t_L g173 ( .A(n_154), .B(n_135), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_166), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_148), .B(n_114), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_148), .B(n_106), .Y(n_178) );
NOR3xp33_ASAP7_75t_L g179 ( .A(n_154), .B(n_118), .C(n_138), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_161), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_161), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_150), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_150), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_149), .B(n_115), .Y(n_189) );
AND2x6_ASAP7_75t_L g190 ( .A(n_152), .B(n_136), .Y(n_190) );
OR2x6_ASAP7_75t_L g191 ( .A(n_152), .B(n_140), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_153), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_149), .B(n_106), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_180), .B(n_151), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_182), .B(n_151), .Y(n_196) );
INVxp67_ASAP7_75t_SL g197 ( .A(n_171), .Y(n_197) );
BUFx12f_ASAP7_75t_L g198 ( .A(n_173), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_194), .B(n_156), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_175), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_190), .B(n_156), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_169), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_174), .B(n_108), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_177), .B(n_157), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_L g205 ( .A1(n_187), .A2(n_157), .B(n_160), .C(n_121), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_191), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_185), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_170), .B(n_108), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_190), .B(n_160), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_187), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
OR2x2_ASAP7_75t_L g214 ( .A(n_173), .B(n_146), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_178), .B(n_113), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_187), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_183), .B(n_113), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_173), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_190), .B(n_132), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_183), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_183), .B(n_132), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_191), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_189), .B(n_133), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_185), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_186), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
OR2x6_ASAP7_75t_L g227 ( .A(n_173), .B(n_130), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_186), .B(n_133), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_191), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_190), .B(n_137), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_190), .B(n_137), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_198), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_200), .A2(n_168), .B(n_167), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_222), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_179), .B(n_167), .C(n_168), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_200), .A2(n_172), .B(n_181), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_206), .A2(n_172), .B(n_181), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_206), .A2(n_176), .B(n_188), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_208), .A2(n_176), .B(n_188), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_196), .B(n_190), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_195), .A2(n_117), .B(n_120), .C(n_129), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_196), .B(n_117), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_196), .B(n_122), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_207), .B(n_141), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_208), .A2(n_192), .B(n_193), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_192), .B(n_193), .Y(n_247) );
NOR2x1p5_ASAP7_75t_SL g248 ( .A(n_210), .B(n_184), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_202), .A2(n_139), .B(n_126), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_141), .B1(n_124), .B2(n_144), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_225), .A2(n_192), .B(n_184), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_196), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_227), .A2(n_123), .B1(n_134), .B2(n_103), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_199), .B(n_119), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_210), .A2(n_128), .B(n_139), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_127), .B1(n_131), .B2(n_142), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_199), .B(n_136), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_216), .B(n_128), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_214), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_210), .A2(n_213), .B(n_220), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_SL g262 ( .A1(n_202), .A2(n_165), .B(n_153), .C(n_162), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_213), .A2(n_147), .B(n_163), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_217), .A2(n_147), .B(n_163), .C(n_158), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_249), .A2(n_202), .B(n_224), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_260), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_261), .A2(n_224), .B(n_213), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_234), .B(n_212), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_253), .B(n_204), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_243), .Y(n_271) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_256), .A2(n_205), .B(n_224), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_244), .B(n_218), .Y(n_273) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_259), .A2(n_201), .B(n_220), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_233), .A2(n_221), .B(n_220), .Y(n_275) );
CKINVDCx11_ASAP7_75t_R g276 ( .A(n_234), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_244), .A2(n_227), .B1(n_198), .B2(n_229), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_255), .B(n_214), .Y(n_279) );
CKINVDCx11_ASAP7_75t_R g280 ( .A(n_257), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_239), .A2(n_228), .B(n_211), .Y(n_281) );
AOI221x1_ASAP7_75t_L g282 ( .A1(n_254), .A2(n_211), .B1(n_230), .B2(n_201), .C(n_226), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_235), .A2(n_223), .B(n_226), .C(n_212), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_246), .A2(n_227), .B(n_231), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_242), .B(n_198), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_247), .A2(n_219), .B(n_230), .Y(n_286) );
INVx5_ASAP7_75t_L g287 ( .A(n_252), .Y(n_287) );
AO31x2_ASAP7_75t_L g288 ( .A1(n_258), .A2(n_147), .A3(n_163), .B(n_158), .Y(n_288) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_263), .A2(n_226), .B(n_147), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_241), .B(n_209), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_267), .B(n_241), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_269), .B(n_248), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_269), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_269), .B(n_212), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_289), .Y(n_295) );
BUFx8_ASAP7_75t_L g296 ( .A(n_271), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_279), .B(n_232), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_266), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_265), .A2(n_259), .B(n_158), .Y(n_299) );
BUFx8_ASAP7_75t_SL g300 ( .A(n_285), .Y(n_300) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_283), .A2(n_251), .B(n_262), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_268), .A2(n_226), .B(n_245), .Y(n_302) );
AOI21x1_ASAP7_75t_L g303 ( .A1(n_282), .A2(n_262), .B(n_203), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_287), .B(n_216), .Y(n_304) );
OAI21x1_ASAP7_75t_SL g305 ( .A1(n_278), .A2(n_207), .B(n_250), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_283), .A2(n_264), .B(n_215), .Y(n_307) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_270), .B(n_207), .Y(n_308) );
INVx6_ASAP7_75t_L g309 ( .A(n_287), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_287), .B(n_216), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_306), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_311), .Y(n_314) );
OA21x2_ASAP7_75t_L g315 ( .A1(n_301), .A2(n_277), .B(n_275), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_311), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_300), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_306), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_292), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_312), .Y(n_320) );
CKINVDCx6p67_ASAP7_75t_R g321 ( .A(n_304), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_311), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_312), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_311), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_296), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_311), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_292), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_311), .Y(n_328) );
AO21x2_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_281), .B(n_284), .Y(n_329) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_307), .A2(n_286), .B(n_290), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_311), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_293), .B(n_273), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_292), .B(n_288), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_295), .Y(n_334) );
AO21x2_ASAP7_75t_L g335 ( .A1(n_307), .A2(n_290), .B(n_273), .Y(n_335) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_302), .A2(n_288), .B(n_274), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
OA21x2_ASAP7_75t_L g338 ( .A1(n_302), .A2(n_274), .B(n_272), .Y(n_338) );
AO21x2_ASAP7_75t_L g339 ( .A1(n_307), .A2(n_272), .B(n_155), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_313), .B(n_292), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_313), .B(n_292), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_318), .B(n_298), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_321), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_313), .B(n_293), .Y(n_346) );
OR2x6_ASAP7_75t_L g347 ( .A(n_319), .B(n_295), .Y(n_347) );
NOR2x1_ASAP7_75t_SL g348 ( .A(n_319), .B(n_307), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_320), .Y(n_349) );
NAND2x1p5_ASAP7_75t_SL g350 ( .A(n_334), .B(n_291), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_320), .B(n_295), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_323), .B(n_295), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_327), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_339), .A2(n_303), .B(n_305), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_323), .B(n_291), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_323), .B(n_298), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_333), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_319), .B(n_293), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_314), .Y(n_364) );
AO21x2_ASAP7_75t_L g365 ( .A1(n_339), .A2(n_303), .B(n_305), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_324), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_293), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_314), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_319), .B(n_293), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_335), .B(n_291), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_333), .B(n_294), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_314), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_322), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_322), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_335), .B(n_308), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_322), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_333), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_333), .B(n_304), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_339), .B(n_299), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_322), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_328), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_339), .B(n_299), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_357), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_341), .B(n_328), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_357), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_359), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_356), .B(n_335), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_356), .B(n_335), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_343), .B(n_335), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_359), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_343), .B(n_335), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_351), .B(n_337), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_341), .B(n_328), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_371), .B(n_328), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_351), .B(n_337), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_373), .B(n_321), .Y(n_400) );
INVx5_ASAP7_75t_L g401 ( .A(n_347), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_346), .B(n_337), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_373), .B(n_321), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_346), .B(n_337), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_341), .B(n_331), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_362), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_342), .B(n_331), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_345), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_345), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_371), .B(n_337), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_359), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_342), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_360), .B(n_331), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_342), .Y(n_414) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_362), .B(n_321), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_363), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_364), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_364), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_363), .B(n_337), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_372), .B(n_331), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_362), .B(n_334), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_372), .B(n_316), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_366), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_378), .B(n_316), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_366), .B(n_332), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_362), .B(n_378), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_364), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_369), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_368), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_380), .B(n_339), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_369), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_380), .B(n_339), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_354), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_352), .B(n_332), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_381), .B(n_334), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_354), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_352), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_360), .B(n_338), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_352), .Y(n_439) );
AND4x1_ASAP7_75t_L g440 ( .A(n_344), .B(n_317), .C(n_297), .D(n_280), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_353), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_368), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_381), .B(n_334), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_353), .B(n_332), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_353), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_358), .B(n_330), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_358), .B(n_330), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_370), .Y(n_448) );
NAND2x1_ASAP7_75t_SL g449 ( .A(n_361), .B(n_317), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_344), .B(n_330), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_344), .A2(n_325), .B1(n_308), .B2(n_297), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_368), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_384), .B(n_338), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_395), .B(n_377), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_440), .B(n_280), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_391), .B(n_377), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_436), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_449), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_390), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_416), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_401), .B(n_370), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_412), .B(n_361), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_428), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_414), .B(n_384), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_431), .Y(n_468) );
OAI21xp33_ASAP7_75t_SL g469 ( .A1(n_400), .A2(n_347), .B(n_367), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_387), .B(n_348), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_392), .B(n_330), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_410), .B(n_350), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_434), .B(n_350), .Y(n_473) );
AND3x2_ASAP7_75t_L g474 ( .A(n_408), .B(n_325), .C(n_382), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_409), .Y(n_475) );
OR2x6_ASAP7_75t_L g476 ( .A(n_403), .B(n_347), .Y(n_476) );
AOI21xp33_ASAP7_75t_L g477 ( .A1(n_446), .A2(n_330), .B(n_365), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_413), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_386), .B(n_382), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_397), .B(n_348), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_401), .B(n_347), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_401), .B(n_347), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_405), .B(n_382), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_453), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_444), .B(n_350), .Y(n_486) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_389), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_398), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_433), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_388), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_405), .B(n_407), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_407), .B(n_385), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_393), .B(n_374), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_393), .B(n_385), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_437), .B(n_374), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_448), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_439), .B(n_385), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_441), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_445), .Y(n_499) );
AND2x2_ASAP7_75t_SL g500 ( .A(n_415), .B(n_308), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_401), .B(n_374), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_435), .B(n_375), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_419), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_396), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_398), .B(n_375), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_435), .B(n_375), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_447), .B(n_376), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_446), .B(n_453), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_435), .B(n_376), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_399), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_425), .B(n_376), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_402), .B(n_379), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_438), .B(n_379), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_443), .B(n_379), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_438), .B(n_430), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_443), .B(n_383), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_404), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_443), .B(n_383), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_430), .B(n_383), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_389), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_394), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_394), .B(n_355), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_411), .B(n_355), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_426), .B(n_355), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_411), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_401), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_426), .B(n_355), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_426), .B(n_365), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_422), .B(n_365), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_417), .Y(n_530) );
NAND2x1_ASAP7_75t_L g531 ( .A(n_406), .B(n_340), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_422), .B(n_365), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_417), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_418), .B(n_340), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_418), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_517), .B(n_432), .Y(n_536) );
AOI32xp33_ASAP7_75t_L g537 ( .A1(n_469), .A2(n_451), .A3(n_406), .B1(n_432), .B2(n_424), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_500), .A2(n_406), .B(n_308), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_488), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_493), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_491), .B(n_424), .Y(n_541) );
INVxp33_ASAP7_75t_L g542 ( .A(n_456), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_475), .Y(n_543) );
AOI21xp33_ASAP7_75t_SL g544 ( .A1(n_462), .A2(n_5), .B(n_6), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_515), .B(n_420), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_515), .B(n_427), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_482), .A2(n_296), .B1(n_421), .B2(n_429), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_489), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_503), .B(n_427), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_476), .B(n_421), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_485), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_429), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_476), .B(n_421), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_505), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_510), .B(n_442), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_525), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_484), .B(n_442), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_508), .B(n_452), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_458), .A2(n_162), .B(n_165), .C(n_452), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_458), .B(n_329), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_467), .B(n_329), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_476), .B(n_340), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_492), .B(n_340), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_467), .A2(n_155), .B(n_164), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_487), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_460), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_520), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_461), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_459), .A2(n_296), .B1(n_309), .B2(n_276), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_464), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_465), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_508), .B(n_315), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_459), .A2(n_309), .B1(n_326), .B2(n_294), .Y(n_574) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_526), .A2(n_296), .B(n_304), .C(n_302), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_468), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_498), .B(n_329), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_499), .B(n_329), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_494), .B(n_329), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_494), .B(n_315), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_490), .B(n_315), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_470), .B(n_338), .Y(n_582) );
OAI211xp5_ASAP7_75t_L g583 ( .A1(n_471), .A2(n_276), .B(n_315), .C(n_165), .Y(n_583) );
NAND3xp33_ASAP7_75t_SL g584 ( .A(n_462), .B(n_310), .C(n_294), .Y(n_584) );
NAND2x1p5_ASAP7_75t_L g585 ( .A(n_526), .B(n_304), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_481), .B(n_483), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_513), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g588 ( .A1(n_481), .A2(n_296), .B(n_222), .C(n_162), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_457), .B(n_315), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_513), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_479), .B(n_5), .Y(n_591) );
AO22x1_ASAP7_75t_L g592 ( .A1(n_483), .A2(n_326), .B1(n_287), .B2(n_207), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_512), .Y(n_593) );
INVxp67_ASAP7_75t_SL g594 ( .A(n_507), .Y(n_594) );
OR2x6_ASAP7_75t_L g595 ( .A(n_531), .B(n_326), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_480), .B(n_338), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_463), .B(n_338), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_502), .B(n_338), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_506), .B(n_326), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_521), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_466), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_507), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_457), .B(n_315), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_479), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_511), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_509), .B(n_326), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_511), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_472), .Y(n_608) );
NOR2x1p5_ASAP7_75t_SL g609 ( .A(n_522), .B(n_315), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_527), .A2(n_309), .B1(n_326), .B2(n_336), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_605), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_608), .B(n_529), .Y(n_612) );
AOI21xp33_ASAP7_75t_SL g613 ( .A1(n_537), .A2(n_486), .B(n_473), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_541), .B(n_532), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_586), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_538), .A2(n_471), .B1(n_455), .B2(n_477), .C(n_497), .Y(n_616) );
XOR2x2_ASAP7_75t_L g617 ( .A(n_570), .B(n_474), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_594), .B(n_455), .Y(n_618) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_538), .A2(n_477), .B1(n_497), .B2(n_528), .C(n_524), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_607), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_544), .A2(n_570), .B(n_584), .C(n_586), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_602), .B(n_454), .Y(n_622) );
AOI221xp5_ASAP7_75t_SL g623 ( .A1(n_604), .A2(n_519), .B1(n_478), .B2(n_514), .C(n_518), .Y(n_623) );
NOR2xp67_ASAP7_75t_SL g624 ( .A(n_583), .B(n_309), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_547), .A2(n_519), .B1(n_501), .B2(n_527), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_567), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g627 ( .A(n_544), .B(n_155), .C(n_164), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_547), .A2(n_501), .B1(n_495), .B2(n_516), .Y(n_628) );
OAI322xp33_ASAP7_75t_L g629 ( .A1(n_591), .A2(n_523), .A3(n_533), .B1(n_530), .B2(n_535), .C1(n_534), .C2(n_155), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_557), .B(n_336), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_539), .B(n_336), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_566), .A2(n_309), .B1(n_326), .B2(n_336), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_554), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_542), .B(n_7), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_561), .A2(n_162), .B1(n_165), .B2(n_164), .C(n_155), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_569), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g637 ( .A1(n_574), .A2(n_7), .B(n_8), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_556), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_597), .B(n_336), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_571), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_572), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_576), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_582), .B(n_336), .Y(n_643) );
OAI21xp33_ASAP7_75t_L g644 ( .A1(n_609), .A2(n_155), .B(n_164), .Y(n_644) );
OAI31xp33_ASAP7_75t_L g645 ( .A1(n_588), .A2(n_294), .A3(n_310), .B(n_222), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_559), .A2(n_310), .B(n_165), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_543), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_550), .B(n_326), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_596), .B(n_336), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_548), .Y(n_650) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_565), .B(n_164), .C(n_155), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_610), .B(n_326), .Y(n_652) );
NOR4xp25_ASAP7_75t_L g653 ( .A(n_560), .B(n_162), .C(n_9), .D(n_10), .Y(n_653) );
AOI32xp33_ASAP7_75t_L g654 ( .A1(n_550), .A2(n_553), .A3(n_601), .B1(n_587), .B2(n_590), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_553), .A2(n_309), .B1(n_299), .B2(n_310), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_593), .B(n_155), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_573), .A2(n_299), .B1(n_164), .B2(n_272), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_573), .A2(n_299), .B1(n_164), .B2(n_216), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_546), .B(n_164), .Y(n_659) );
OAI21xp33_ASAP7_75t_L g660 ( .A1(n_562), .A2(n_8), .B(n_9), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_621), .A2(n_565), .B(n_575), .C(n_579), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_615), .A2(n_545), .B1(n_585), .B2(n_580), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_656), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_623), .B(n_589), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_615), .A2(n_558), .B1(n_595), .B2(n_536), .Y(n_665) );
OA21x2_ASAP7_75t_SL g666 ( .A1(n_652), .A2(n_563), .B(n_603), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_654), .A2(n_563), .B(n_540), .C(n_551), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_613), .A2(n_578), .B1(n_577), .B2(n_581), .C(n_598), .Y(n_668) );
OAI21x1_ASAP7_75t_SL g669 ( .A1(n_625), .A2(n_549), .B(n_552), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g670 ( .A(n_637), .B(n_592), .C(n_555), .Y(n_670) );
OAI221xp5_ASAP7_75t_L g671 ( .A1(n_619), .A2(n_595), .B1(n_600), .B2(n_568), .C(n_564), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_659), .Y(n_672) );
NOR4xp25_ASAP7_75t_L g673 ( .A(n_629), .B(n_606), .C(n_599), .D(n_13), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_629), .A2(n_595), .B(n_216), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_628), .A2(n_216), .B1(n_12), .B2(n_13), .Y(n_675) );
AOI321xp33_ASAP7_75t_L g676 ( .A1(n_616), .A2(n_11), .A3(n_12), .B1(n_14), .B2(n_15), .C(n_16), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_653), .A2(n_14), .B1(n_15), .B2(n_17), .C(n_18), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_633), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_617), .B(n_19), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_618), .B(n_20), .Y(n_680) );
INVx3_ASAP7_75t_L g681 ( .A(n_648), .Y(n_681) );
OAI21xp5_ASAP7_75t_SL g682 ( .A1(n_627), .A2(n_21), .B(n_100), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_650), .A2(n_21), .B1(n_23), .B2(n_24), .C(n_25), .Y(n_683) );
A2O1A1Ixp33_ASAP7_75t_L g684 ( .A1(n_645), .A2(n_26), .B(n_27), .C(n_28), .Y(n_684) );
AOI32xp33_ASAP7_75t_L g685 ( .A1(n_634), .A2(n_29), .A3(n_33), .B1(n_34), .B2(n_35), .Y(n_685) );
NOR4xp25_ASAP7_75t_L g686 ( .A(n_660), .B(n_644), .C(n_636), .D(n_640), .Y(n_686) );
NAND4xp25_ASAP7_75t_L g687 ( .A(n_645), .B(n_36), .C(n_37), .D(n_38), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_627), .B(n_48), .C(n_49), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_655), .A2(n_51), .B(n_54), .C(n_56), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_611), .B(n_57), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_622), .A2(n_60), .B(n_62), .Y(n_691) );
OAI221xp5_ASAP7_75t_SL g692 ( .A1(n_612), .A2(n_63), .B1(n_66), .B2(n_68), .C(n_70), .Y(n_692) );
OAI211xp5_ASAP7_75t_SL g693 ( .A1(n_631), .A2(n_71), .B(n_72), .C(n_73), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g694 ( .A1(n_646), .A2(n_74), .B(n_77), .C(n_78), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_632), .A2(n_79), .B(n_80), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_624), .A2(n_81), .B(n_84), .C(n_87), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_651), .A2(n_91), .B(n_92), .Y(n_697) );
AOI211x1_ASAP7_75t_SL g698 ( .A1(n_638), .A2(n_97), .B(n_651), .C(n_626), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_643), .A2(n_649), .B1(n_639), .B2(n_614), .Y(n_699) );
OAI221xp5_ASAP7_75t_SL g700 ( .A1(n_630), .A2(n_635), .B1(n_620), .B2(n_641), .C(n_642), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_647), .A2(n_658), .B(n_657), .C(n_648), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_623), .B(n_613), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_673), .B(n_686), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_702), .B(n_664), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g705 ( .A1(n_679), .A2(n_670), .B(n_676), .C(n_682), .Y(n_705) );
AOI211xp5_ASAP7_75t_L g706 ( .A1(n_700), .A2(n_661), .B(n_675), .C(n_667), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_668), .A2(n_671), .B1(n_669), .B2(n_672), .C(n_663), .Y(n_707) );
OAI211xp5_ASAP7_75t_SL g708 ( .A1(n_698), .A2(n_677), .B(n_680), .C(n_685), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_662), .Y(n_709) );
NOR4xp25_ASAP7_75t_L g710 ( .A(n_678), .B(n_701), .C(n_699), .D(n_665), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_704), .B(n_709), .Y(n_711) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_703), .B(n_687), .Y(n_712) );
NOR3xp33_ASAP7_75t_SL g713 ( .A(n_705), .B(n_692), .C(n_689), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_707), .Y(n_714) );
AND2x4_ASAP7_75t_L g715 ( .A(n_711), .B(n_681), .Y(n_715) );
NAND3x1_ASAP7_75t_SL g716 ( .A(n_712), .B(n_710), .C(n_706), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_714), .B(n_681), .Y(n_717) );
XNOR2xp5_ASAP7_75t_L g718 ( .A(n_716), .B(n_713), .Y(n_718) );
INVx2_ASAP7_75t_SL g719 ( .A(n_715), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_718), .A2(n_717), .B1(n_708), .B2(n_674), .C(n_683), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_719), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_666), .B1(n_684), .B2(n_696), .Y(n_722) );
OAI21x1_ASAP7_75t_L g723 ( .A1(n_720), .A2(n_697), .B(n_691), .Y(n_723) );
OR2x6_ASAP7_75t_L g724 ( .A(n_723), .B(n_690), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_724), .B(n_722), .Y(n_725) );
NAND2xp33_ASAP7_75t_L g726 ( .A(n_725), .B(n_688), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_695), .B1(n_693), .B2(n_694), .Y(n_727) );
endmodule