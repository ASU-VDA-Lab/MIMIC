module fake_jpeg_24607_n_34 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_34);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_15),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_6),
.B(n_12),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_23),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_5),
.B(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_22),
.B1(n_17),
.B2(n_16),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.C(n_28),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_0),
.B1(n_10),
.B2(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_26),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_13),
.B(n_14),
.Y(n_34)
);


endmodule