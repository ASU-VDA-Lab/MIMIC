module fake_jpeg_18741_n_86 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_86);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_86;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_0),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_22),
.B1(n_26),
.B2(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_15),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_15),
.C(n_22),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_31),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_31),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_23),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_33),
.A3(n_36),
.B1(n_17),
.B2(n_20),
.Y(n_55)
);

NAND5xp2_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_39),
.C(n_10),
.D(n_23),
.E(n_19),
.Y(n_58)
);

XNOR2x2_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_41),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_59),
.B(n_64),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_62),
.B1(n_48),
.B2(n_56),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_37),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_42),
.C(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_11),
.B(n_20),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_70),
.B1(n_59),
.B2(n_49),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_51),
.B(n_16),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_64),
.B(n_65),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_61),
.C(n_70),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_49),
.B1(n_18),
.B2(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_74),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_1),
.Y(n_78)
);

AOI21x1_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_65),
.B(n_1),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_77),
.B(n_75),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_79),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_77),
.B(n_4),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_6),
.C(n_8),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_82),
.C(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_83),
.Y(n_86)
);


endmodule