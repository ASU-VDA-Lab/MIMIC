module real_jpeg_20845_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_0),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_0),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_0),
.A2(n_29),
.B1(n_31),
.B2(n_64),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_1),
.A2(n_47),
.B1(n_59),
.B2(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_29),
.B1(n_31),
.B2(n_47),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_72),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_56),
.B1(n_63),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_67),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_29),
.B1(n_31),
.B2(n_67),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_4),
.A2(n_56),
.B1(n_63),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_4),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_121),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_121),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_4),
.A2(n_29),
.B1(n_31),
.B2(n_121),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_56),
.B1(n_63),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_99),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_5),
.A2(n_29),
.B1(n_31),
.B2(n_99),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_99),
.Y(n_194)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_85)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_10),
.A2(n_29),
.B1(n_31),
.B2(n_49),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_11),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_11),
.B(n_58),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_11),
.A2(n_29),
.B(n_43),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_110),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_11),
.B(n_79),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_11),
.A2(n_60),
.B(n_209),
.Y(n_208)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_13),
.A2(n_29),
.B1(n_31),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_75),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_14),
.A2(n_42),
.A3(n_60),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_100),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_21),
.B(n_100),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_87),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_80),
.B2(n_81),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_50),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_38),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_26),
.B(n_38),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_27),
.A2(n_35),
.B1(n_90),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_27),
.A2(n_35),
.B1(n_113),
.B2(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_27),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_27),
.A2(n_33),
.B1(n_164),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_27),
.A2(n_35),
.B1(n_166),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_27),
.A2(n_35),
.B1(n_153),
.B2(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_28),
.B(n_110),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_31),
.B1(n_43),
.B2(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_31),
.B(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_34),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_161)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_39),
.A2(n_45),
.B1(n_48),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_39),
.A2(n_45),
.B1(n_92),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_39),
.A2(n_45),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_39),
.A2(n_45),
.B1(n_174),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_39),
.A2(n_45),
.B1(n_194),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_39),
.A2(n_45),
.B1(n_132),
.B2(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_41),
.B(n_75),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_42),
.A2(n_44),
.B(n_110),
.C(n_170),
.Y(n_169)
);

CKINVDCx9p33_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_45),
.B(n_110),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_68),
.B2(n_69),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_62),
.B1(n_65),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_53),
.A2(n_65),
.B1(n_98),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_54),
.A2(n_58),
.B1(n_109),
.B2(n_120),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_60),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g109 ( 
.A(n_56),
.B(n_110),
.CON(n_109),
.SN(n_109)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_59),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_59),
.B(n_110),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_73),
.A2(n_79),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_77),
.B1(n_95),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_74),
.A2(n_77),
.B1(n_116),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_74),
.A2(n_77),
.B1(n_148),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_96),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_91),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.C(n_105),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_101),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_105),
.A2(n_106),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.C(n_117),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_112),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_154),
.B(n_237),
.C(n_243),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_139),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_126),
.B(n_139),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_128),
.B(n_129),
.C(n_137),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.C(n_136),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_140),
.B(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_151),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_146),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_150),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_236),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_231),
.B(n_235),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_217),
.B(n_230),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_198),
.B(n_216),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_186),
.B(n_197),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_175),
.B(n_185),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_167),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_171),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_180),
.B(n_184),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_200),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_206),
.B1(n_214),
.B2(n_215),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_201),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_207),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_219),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_227),
.C(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_227),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);


endmodule