module fake_aes_2721_n_402 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_402);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_402;
wire n_117;
wire n_361;
wire n_185;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_391;
wire n_235;
wire n_243;
wire n_394;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_88;
wire n_107;
wire n_254;
wire n_262;
wire n_239;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_396;
wire n_168;
wire n_398;
wire n_134;
wire n_233;
wire n_82;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_350;
wire n_164;
wire n_175;
wire n_145;
wire n_290;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_55), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_65), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_61), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_51), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_67), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_37), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_59), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_42), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_48), .Y(n_93) );
INVxp33_ASAP7_75t_L g94 ( .A(n_49), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_60), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_77), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_76), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_70), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_35), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_72), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_44), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_33), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_62), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_56), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_36), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_32), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_34), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_68), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_31), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_26), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_42), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_63), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_36), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_38), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_35), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_54), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_66), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_18), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_113), .B(n_82), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_113), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_91), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_107), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_96), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_107), .Y(n_135) );
BUFx12f_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_102), .B(n_0), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_117), .B(n_1), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_107), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_94), .B(n_1), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_112), .B(n_2), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_81), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_81), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_83), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g148 ( .A(n_124), .B(n_45), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_124), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_88), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_128), .B(n_108), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_128), .B(n_101), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_128), .B(n_118), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_128), .B(n_101), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_145), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_149), .B(n_106), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_149), .B(n_106), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_130), .A2(n_110), .B1(n_116), .B2(n_114), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_126), .B(n_100), .Y(n_163) );
INVxp67_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_141), .B(n_118), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_145), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_125), .B(n_82), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_130), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_130), .A2(n_110), .B1(n_116), .B2(n_114), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_125), .B(n_100), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
NAND3x1_ASAP7_75t_L g176 ( .A(n_137), .B(n_123), .C(n_122), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_127), .B(n_111), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_146), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_141), .B(n_87), .Y(n_179) );
AND2x4_ASAP7_75t_L g180 ( .A(n_131), .B(n_111), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_151), .B(n_137), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_167), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_166), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_154), .A2(n_138), .B1(n_137), .B2(n_142), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_171), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_172), .Y(n_192) );
NOR2x1p5_ASAP7_75t_L g193 ( .A(n_151), .B(n_136), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_172), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_175), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
AND3x2_ASAP7_75t_SL g201 ( .A(n_167), .B(n_148), .C(n_147), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_161), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_170), .B(n_134), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_164), .B(n_138), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_165), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_177), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_181), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_177), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_180), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_169), .B(n_132), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_152), .B(n_139), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_152), .B(n_143), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
INVx5_ASAP7_75t_L g221 ( .A(n_165), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_181), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_183), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_189), .A2(n_173), .B1(n_162), .B2(n_176), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_217), .B(n_193), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_217), .B(n_165), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_208), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_215), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_186), .B(n_179), .Y(n_230) );
INVx5_ASAP7_75t_L g231 ( .A(n_185), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_185), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_185), .Y(n_233) );
BUFx12f_ASAP7_75t_L g234 ( .A(n_207), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_209), .B(n_174), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_216), .Y(n_236) );
BUFx4_ASAP7_75t_SL g237 ( .A(n_199), .Y(n_237) );
INVx4_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_218), .A2(n_163), .B(n_156), .Y(n_239) );
INVx5_ASAP7_75t_SL g240 ( .A(n_187), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_219), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_223), .B(n_159), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_223), .B(n_159), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_188), .B(n_160), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_221), .B(n_160), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_204), .A2(n_150), .B1(n_147), .B2(n_144), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_191), .Y(n_247) );
AOI21x1_ASAP7_75t_L g248 ( .A1(n_192), .A2(n_196), .B(n_194), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
NOR3xp33_ASAP7_75t_L g250 ( .A(n_211), .B(n_109), .C(n_92), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_194), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_196), .Y(n_252) );
INVx4_ASAP7_75t_L g253 ( .A(n_204), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_197), .A2(n_155), .B(n_153), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_225), .A2(n_214), .B1(n_220), .B2(n_213), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_224), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_232), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_226), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_230), .A2(n_205), .B1(n_222), .B2(n_212), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_234), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_244), .Y(n_261) );
INVx6_ASAP7_75t_L g262 ( .A(n_231), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_250), .A2(n_222), .B1(n_212), .B2(n_184), .Y(n_263) );
INVx4_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_251), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_252), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_227), .A2(n_184), .B1(n_200), .B2(n_120), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_237), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_235), .B(n_184), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_242), .A2(n_200), .B1(n_120), .B2(n_99), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_229), .Y(n_272) );
NOR2x1_ASAP7_75t_SL g273 ( .A(n_238), .B(n_190), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_232), .Y(n_274) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_248), .A2(n_201), .B(n_150), .Y(n_275) );
INVx4_ASAP7_75t_SL g276 ( .A(n_245), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_243), .A2(n_103), .B1(n_105), .B2(n_104), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_241), .B(n_206), .Y(n_279) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_247), .A2(n_115), .B1(n_121), .B2(n_119), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_254), .A2(n_198), .B(n_195), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g282 ( .A1(n_239), .A2(n_203), .B(n_202), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_232), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_249), .A2(n_93), .B1(n_95), .B2(n_84), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_240), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_255), .A2(n_240), .B1(n_246), .B2(n_233), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_256), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_276), .B(n_253), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_265), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_266), .Y(n_290) );
OR2x6_ASAP7_75t_L g291 ( .A(n_268), .B(n_238), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_264), .Y(n_292) );
AOI21xp33_ASAP7_75t_L g293 ( .A1(n_275), .A2(n_98), .B(n_97), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
AO221x2_ASAP7_75t_L g295 ( .A1(n_280), .A2(n_284), .B1(n_261), .B2(n_272), .C(n_278), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_257), .Y(n_296) );
OAI22xp5_ASAP7_75t_SL g297 ( .A1(n_260), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_297) );
INVx4_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
AOI21xp33_ASAP7_75t_L g299 ( .A1(n_259), .A2(n_135), .B(n_133), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_270), .B(n_129), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_258), .B(n_6), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_257), .Y(n_302) );
OR2x6_ASAP7_75t_L g303 ( .A(n_262), .B(n_7), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_257), .Y(n_304) );
OR2x6_ASAP7_75t_L g305 ( .A(n_262), .B(n_8), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
NAND2x1_ASAP7_75t_L g307 ( .A(n_285), .B(n_140), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_277), .A2(n_182), .B1(n_168), .B2(n_12), .C(n_13), .Y(n_308) );
AND2x6_ASAP7_75t_L g309 ( .A(n_274), .B(n_46), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_263), .A2(n_9), .B1(n_14), .B2(n_15), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_263), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_290), .Y(n_313) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_293), .A2(n_282), .B(n_281), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_303), .A2(n_259), .B1(n_271), .B2(n_267), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_287), .Y(n_316) );
AOI222xp33_ASAP7_75t_L g317 ( .A1(n_297), .A2(n_273), .B1(n_20), .B2(n_21), .C1(n_22), .C2(n_23), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_295), .A2(n_283), .B1(n_24), .B2(n_25), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_306), .B(n_27), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_305), .A2(n_28), .B1(n_29), .B2(n_30), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_292), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_286), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
INVx4_ASAP7_75t_SL g326 ( .A(n_309), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_291), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_291), .B(n_50), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_288), .B(n_52), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_296), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_298), .B(n_53), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_312), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_317), .A2(n_308), .B1(n_311), .B2(n_310), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_326), .B(n_309), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_314), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_318), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_323), .Y(n_339) );
AOI22xp33_ASAP7_75t_SL g340 ( .A1(n_324), .A2(n_309), .B1(n_296), .B2(n_302), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_327), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_326), .B(n_302), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_322), .A2(n_307), .B1(n_299), .B2(n_304), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_325), .B(n_302), .Y(n_345) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_329), .B(n_330), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_321), .B(n_304), .Y(n_347) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_319), .B(n_58), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_315), .A2(n_69), .B1(n_71), .B2(n_73), .Y(n_350) );
AND2x2_ASAP7_75t_SL g351 ( .A(n_332), .B(n_74), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_333), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_344), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_336), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_344), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_345), .B(n_331), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_338), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_349), .Y(n_359) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_339), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_349), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_335), .B(n_78), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_341), .B(n_79), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_351), .A2(n_346), .B1(n_334), .B2(n_348), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_352), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_347), .Y(n_366) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_337), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_353), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_355), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_358), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_366), .B(n_340), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_365), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_364), .A2(n_343), .B(n_350), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_360), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_359), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_361), .B(n_342), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_357), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_354), .B(n_356), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_356), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_368), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_369), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_370), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_377), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_374), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_371), .Y(n_385) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_373), .B(n_362), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_372), .B(n_363), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_386), .B(n_383), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_384), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_384), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_389), .Y(n_391) );
NOR3xp33_ASAP7_75t_L g392 ( .A(n_388), .B(n_387), .C(n_385), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_391), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_392), .A2(n_390), .B1(n_389), .B2(n_382), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_394), .B(n_381), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_393), .B(n_380), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_396), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_395), .Y(n_398) );
OR2x2_ASAP7_75t_SL g399 ( .A(n_398), .B(n_397), .Y(n_399) );
OR2x6_ASAP7_75t_L g400 ( .A(n_399), .B(n_376), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_400), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_401), .A2(n_367), .B1(n_375), .B2(n_379), .C(n_378), .Y(n_402) );
endmodule