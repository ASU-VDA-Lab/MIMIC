module real_jpeg_27556_n_12 (n_5, n_4, n_8, n_0, n_280, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_280;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_249;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_131;
wire n_47;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g60 ( 
.A(n_0),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_4),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_4),
.A2(n_41),
.B1(n_43),
.B2(n_95),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_95),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_95),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_6),
.A2(n_41),
.B1(n_43),
.B2(n_182),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_182),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_182),
.Y(n_275)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_79),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_9),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_27),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_27),
.B1(n_41),
.B2(n_43),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_11),
.A2(n_31),
.B(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_11),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_11),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_11),
.B(n_32),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_11),
.A2(n_41),
.B(n_121),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_59),
.B(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_11),
.B(n_40),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_271),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_262),
.B(n_270),
.Y(n_13)
);

OAI321xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_231),
.A3(n_255),
.B1(n_260),
.B2(n_261),
.C(n_280),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_212),
.B(n_230),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_193),
.B(n_211),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_113),
.B(n_174),
.C(n_192),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_99),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_19),
.B(n_99),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_66),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_20),
.B(n_67),
.C(n_85),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_52),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_21)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_22),
.B(n_51),
.C(n_52),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_22),
.A2(n_50),
.B1(n_69),
.B2(n_102),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_22),
.B(n_102),
.C(n_199),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_22),
.A2(n_50),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_22),
.B(n_241),
.C(n_252),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_24),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_26),
.A2(n_30),
.B(n_36),
.C(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_28),
.B(n_32),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_28),
.A2(n_32),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g34 ( 
.A(n_33),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_33),
.A2(n_36),
.B(n_42),
.C(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_35),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_36),
.A2(n_41),
.B(n_79),
.C(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_36),
.B(n_65),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_36),
.B(n_80),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_37),
.B(n_108),
.C(n_111),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_37),
.A2(n_51),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_37),
.A2(n_218),
.B(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_37),
.B(n_218),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_39),
.B(n_40),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_39),
.A2(n_40),
.B1(n_238),
.B2(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_40),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_43),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_49),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_47),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_56),
.A2(n_106),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_56),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_56),
.B(n_158),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_56),
.B(n_135),
.C(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_96),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_58),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_61),
.B(n_62),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_61),
.A2(n_65),
.B1(n_94),
.B2(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_94),
.B(n_96),
.Y(n_93)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_84),
.B2(n_85),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.C(n_81),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_69),
.A2(n_86),
.B1(n_87),
.B2(n_102),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_70),
.Y(n_239)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_76),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_76),
.B1(n_80),
.B2(n_89),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_75),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_76),
.A2(n_80),
.B1(n_204),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_80),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_81),
.A2(n_103),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_81),
.A2(n_103),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_81),
.A2(n_103),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_81),
.B(n_237),
.C(n_240),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_81),
.B(n_247),
.C(n_254),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_82),
.A2(n_83),
.B(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_86),
.A2(n_87),
.B1(n_142),
.B2(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_86),
.B(n_93),
.Y(n_185)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_102),
.C(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_87),
.B(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B(n_91),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_107),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_100),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_103),
.B(n_185),
.C(n_187),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_105),
.B(n_107),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_108),
.B(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_173),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_168),
.B(n_172),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_138),
.B(n_167),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_117),
.B(n_126),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_125),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_135),
.C(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_129),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_137),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_137),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_135),
.B(n_180),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_162),
.B(n_166),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_149),
.B(n_161),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_144),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_142),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_146),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_153),
.B(n_160),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_157),
.B(n_159),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_176),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_190),
.B2(n_191),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_184),
.C(n_191),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_180),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_189),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_190),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_195),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_210),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_202),
.C(n_210),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_206),
.A2(n_207),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_222),
.B(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_213),
.B(n_214),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_228),
.B2(n_229),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_221),
.C(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_233),
.C(n_243),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_233),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_228),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_245),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_241),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_244),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_264),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_264),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_267),
.CI(n_269),
.CON(n_264),
.SN(n_264)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_276),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);


endmodule