module fake_jpeg_6723_n_321 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_33),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_14),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_52),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_58),
.Y(n_94)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_29),
.B1(n_36),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_62),
.B1(n_71),
.B2(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_36),
.B1(n_30),
.B2(n_32),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_49),
.Y(n_64)
);

FAx1_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_50),
.CI(n_43),
.CON(n_88),
.SN(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_36),
.B1(n_18),
.B2(n_20),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_29),
.B1(n_36),
.B2(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_76),
.Y(n_79)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_17),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_43),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_45),
.C(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_52),
.B(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_50),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_55),
.B1(n_48),
.B2(n_40),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_98),
.B1(n_69),
.B2(n_48),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_25),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_22),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_55),
.B1(n_48),
.B2(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_100),
.B(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_67),
.B(n_61),
.C(n_73),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_98),
.B(n_78),
.Y(n_134)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_108),
.Y(n_140)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_110),
.C(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_70),
.C(n_56),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_56),
.C(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_86),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_20),
.Y(n_142)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_57),
.B(n_58),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_55),
.B1(n_58),
.B2(n_57),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_144),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_95),
.B(n_79),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_104),
.B1(n_119),
.B2(n_115),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_29),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_88),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_100),
.B1(n_78),
.B2(n_95),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_88),
.C(n_84),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_141),
.C(n_142),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_110),
.B(n_103),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_45),
.B1(n_86),
.B2(n_55),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_106),
.B1(n_122),
.B2(n_111),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_145),
.B1(n_146),
.B2(n_119),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_56),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_54),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_68),
.C(n_46),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_82),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_121),
.B1(n_123),
.B2(n_114),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_86),
.B1(n_99),
.B2(n_48),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_151),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_153),
.B(n_161),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_129),
.C(n_143),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_162),
.B1(n_175),
.B2(n_23),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_115),
.B1(n_41),
.B2(n_99),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_132),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_125),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_173),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_148),
.B(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_75),
.B1(n_87),
.B2(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_129),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_155),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_160),
.B1(n_173),
.B2(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_164),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_187),
.C(n_167),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_142),
.C(n_139),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_75),
.B1(n_23),
.B2(n_65),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_27),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_191),
.B(n_10),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_196),
.A2(n_202),
.B1(n_149),
.B2(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_23),
.B1(n_27),
.B2(n_21),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_197),
.B(n_199),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_217),
.C(n_218),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_212),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_152),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_220),
.B(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_179),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_210),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_188),
.B1(n_201),
.B2(n_186),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_171),
.C(n_161),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_193),
.CI(n_181),
.CON(n_229),
.SN(n_229)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_150),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_169),
.B1(n_162),
.B2(n_155),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_216),
.B1(n_189),
.B2(n_197),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_41),
.B1(n_21),
.B2(n_19),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_38),
.C(n_37),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_38),
.C(n_37),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_222),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_38),
.B(n_37),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_38),
.C(n_37),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_218),
.C(n_204),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_193),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_235),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_242),
.B(n_237),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_244),
.C(n_245),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_194),
.B1(n_195),
.B2(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_233),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_215),
.A2(n_188),
.B1(n_186),
.B2(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_223),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_202),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_243),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_217),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_199),
.C(n_192),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_191),
.C(n_41),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_224),
.C(n_220),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_253),
.C(n_262),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_230),
.B(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_209),
.C(n_205),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_229),
.B(n_241),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_261),
.B(n_263),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_216),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_259),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_41),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_0),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_10),
.B(n_1),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_51),
.C(n_25),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_235),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_271),
.B(n_256),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_51),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_270),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_239),
.B(n_226),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_269),
.B(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_239),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_246),
.B1(n_254),
.B2(n_262),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_273),
.A2(n_279),
.B1(n_19),
.B2(n_26),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_256),
.A2(n_19),
.B1(n_26),
.B2(n_2),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_0),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_25),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_25),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_26),
.B1(n_19),
.B2(n_24),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_282),
.B(n_285),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_0),
.Y(n_293)
);

FAx1_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_26),
.CI(n_1),
.CON(n_285),
.SN(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_265),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_268),
.B(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_288),
.B(n_292),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_291),
.C(n_276),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_51),
.B(n_35),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_278),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_303),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_298),
.B(n_301),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_279),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_3),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_302),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_24),
.C(n_35),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_35),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_283),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_285),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_308),
.B(n_3),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_285),
.B1(n_290),
.B2(n_24),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_13),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_302),
.A3(n_293),
.B1(n_24),
.B2(n_35),
.C1(n_7),
.C2(n_9),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_313),
.A3(n_314),
.B1(n_304),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_310),
.A2(n_4),
.B(n_5),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_311),
.A2(n_309),
.A3(n_304),
.B1(n_6),
.B2(n_7),
.C1(n_9),
.C2(n_4),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_5),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_316),
.C2(n_306),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_5),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_11),
.B(n_12),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_12),
.B(n_13),
.Y(n_321)
);


endmodule