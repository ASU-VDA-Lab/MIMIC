module fake_jpeg_31386_n_528 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_15),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_54),
.B(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_65),
.Y(n_106)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_31),
.B(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_77),
.Y(n_115)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_81),
.B(n_50),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_30),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_105),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_34),
.B(n_16),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_154),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_30),
.B1(n_37),
.B2(n_33),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_110),
.A2(n_127),
.B1(n_148),
.B2(n_38),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_34),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_114),
.B(n_168),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_65),
.A2(n_48),
.B1(n_37),
.B2(n_33),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_50),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_155),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_77),
.A2(n_30),
.B(n_41),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_18),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_22),
.B1(n_51),
.B2(n_35),
.Y(n_148)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_83),
.B(n_35),
.CON(n_154),
.SN(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_90),
.B(n_41),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_104),
.A2(n_22),
.B1(n_36),
.B2(n_18),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_95),
.B1(n_92),
.B2(n_91),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_97),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_88),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_58),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_170),
.Y(n_254)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_172),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_173),
.B(n_195),
.Y(n_238)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_174),
.Y(n_235)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_177),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_189),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_118),
.A2(n_110),
.B1(n_106),
.B2(n_85),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_179),
.A2(n_222),
.B1(n_226),
.B2(n_209),
.Y(n_269)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_181),
.Y(n_230)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g260 ( 
.A(n_186),
.Y(n_260)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_89),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_190),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_191),
.Y(n_264)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_138),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_115),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_197),
.B(n_201),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_130),
.A2(n_84),
.B(n_79),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_202),
.Y(n_247)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_199),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_150),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_200),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_113),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_141),
.A2(n_32),
.B1(n_67),
.B2(n_62),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_209),
.B1(n_164),
.B2(n_151),
.Y(n_243)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_206),
.B(n_207),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_115),
.B(n_32),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_135),
.A2(n_32),
.B1(n_75),
.B2(n_3),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_211),
.B(n_213),
.Y(n_272)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_153),
.Y(n_212)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_216),
.Y(n_256)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_117),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_224),
.Y(n_239)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_220),
.Y(n_261)
);

INVx6_ASAP7_75t_SL g220 ( 
.A(n_142),
.Y(n_220)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_144),
.A2(n_32),
.B1(n_38),
.B2(n_3),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_134),
.B1(n_157),
.B2(n_144),
.Y(n_246)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_131),
.B(n_124),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_158),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_134),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_122),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_227),
.A2(n_228),
.B1(n_5),
.B2(n_6),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_125),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_184),
.A2(n_167),
.B1(n_112),
.B2(n_128),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_219),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_182),
.B(n_151),
.C(n_124),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_244),
.B(n_252),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_159),
.B(n_2),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_245),
.A2(n_222),
.B(n_191),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_246),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_188),
.A2(n_167),
.B1(n_157),
.B2(n_158),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_250),
.A2(n_220),
.B1(n_212),
.B2(n_186),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_182),
.A2(n_149),
.B1(n_2),
.B2(n_4),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_267),
.B1(n_269),
.B2(n_226),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_179),
.B(n_149),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_192),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_202),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_208),
.B(n_1),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_5),
.Y(n_292)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_273),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_169),
.B(n_190),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_276),
.A2(n_266),
.B(n_231),
.Y(n_326)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_278),
.A2(n_287),
.B1(n_261),
.B2(n_239),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_238),
.B(n_178),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_289),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_204),
.B1(n_185),
.B2(n_174),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_282),
.A2(n_285),
.B1(n_298),
.B2(n_305),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_283),
.A2(n_291),
.B(n_294),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_234),
.A2(n_221),
.B1(n_199),
.B2(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_286),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_227),
.B1(n_181),
.B2(n_200),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_272),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_187),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_292),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_247),
.A2(n_217),
.B(n_216),
.Y(n_291)
);

BUFx24_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_260),
.A2(n_218),
.B1(n_210),
.B2(n_214),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_296),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_229),
.B(n_177),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_262),
.B1(n_251),
.B2(n_241),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_234),
.A2(n_219),
.B1(n_6),
.B2(n_7),
.Y(n_298)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_301),
.Y(n_331)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_302),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_232),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_315),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_246),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_260),
.B1(n_230),
.B2(n_268),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_234),
.A2(n_13),
.B1(n_9),
.B2(n_10),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_7),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_306),
.B(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_231),
.B1(n_266),
.B2(n_230),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_247),
.B(n_244),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_310),
.A2(n_247),
.B(n_255),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_270),
.B(n_10),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_311),
.B(n_312),
.Y(n_334)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_261),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_314),
.B(n_275),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_232),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_326),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_R g319 ( 
.A(n_314),
.B(n_246),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_319),
.B(n_309),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_252),
.C(n_259),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_310),
.C(n_297),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_325),
.A2(n_350),
.B1(n_282),
.B2(n_298),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_328),
.A2(n_284),
.B1(n_281),
.B2(n_293),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_340),
.B(n_348),
.Y(n_352)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_276),
.A2(n_246),
.A3(n_262),
.B1(n_251),
.B2(n_264),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_335),
.A2(n_297),
.B(n_285),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_302),
.B1(n_301),
.B2(n_286),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_346),
.Y(n_355)
);

AO21x2_ASAP7_75t_L g340 ( 
.A1(n_291),
.A2(n_264),
.B(n_268),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_296),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_343),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_313),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_289),
.B(n_275),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_313),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_347),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_283),
.A2(n_233),
.B(n_242),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_278),
.A2(n_233),
.B1(n_249),
.B2(n_242),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_342),
.Y(n_351)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_360),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_327),
.B(n_279),
.Y(n_354)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_312),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_356),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_357),
.A2(n_317),
.B(n_348),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_295),
.Y(n_358)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_337),
.B(n_288),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_316),
.B(n_305),
.Y(n_361)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_361),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_362),
.A2(n_380),
.B1(n_381),
.B2(n_340),
.Y(n_390)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_363),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_326),
.C(n_318),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_319),
.A2(n_300),
.B(n_287),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_365),
.A2(n_367),
.B(n_329),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_308),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_369),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_307),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_370),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_338),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_372),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_315),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_373),
.B(n_377),
.Y(n_400)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_345),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_375),
.Y(n_396)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_325),
.A2(n_284),
.B1(n_300),
.B2(n_303),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_376),
.A2(n_383),
.B1(n_284),
.B2(n_340),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_324),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_334),
.B(n_293),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_379),
.B(n_334),
.Y(n_412)
);

INVx8_ASAP7_75t_L g380 ( 
.A(n_340),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_299),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_340),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_387),
.A2(n_388),
.B(n_352),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_357),
.B(n_370),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_375),
.A2(n_323),
.B1(n_335),
.B2(n_317),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_390),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_392),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_378),
.B(n_320),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_393),
.B(n_402),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_380),
.A2(n_321),
.B1(n_332),
.B2(n_331),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_373),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_403),
.C(n_406),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_332),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_399),
.B(n_413),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_331),
.C(n_321),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_330),
.C(n_322),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_330),
.C(n_322),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_407),
.B(n_369),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_340),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_353),
.Y(n_437)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_412),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_355),
.B(n_328),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_379),
.Y(n_414)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_415),
.Y(n_451)
);

INVx13_ASAP7_75t_L g416 ( 
.A(n_409),
.Y(n_416)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_400),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_417),
.B(n_420),
.Y(n_442)
);

BUFx12f_ASAP7_75t_L g420 ( 
.A(n_388),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_425),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_426),
.A2(n_363),
.B1(n_351),
.B2(n_398),
.Y(n_457)
);

INVx13_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_427),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_407),
.B(n_386),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_405),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_396),
.B(n_372),
.Y(n_430)
);

XOR2x2_ASAP7_75t_SL g432 ( 
.A(n_402),
.B(n_367),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_432),
.B(n_435),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_411),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_433),
.A2(n_389),
.B1(n_391),
.B2(n_410),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_393),
.B(n_397),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_371),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_436),
.B(n_437),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_361),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_438),
.A2(n_439),
.B1(n_423),
.B2(n_384),
.Y(n_445)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_371),
.C(n_358),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_431),
.B(n_403),
.C(n_413),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_441),
.C(n_447),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_387),
.C(n_410),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_418),
.Y(n_467)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_395),
.B1(n_384),
.B2(n_376),
.Y(n_446)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_404),
.C(n_401),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_424),
.A2(n_404),
.B1(n_380),
.B2(n_365),
.Y(n_448)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_437),
.A2(n_392),
.B1(n_383),
.B2(n_366),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_450),
.A2(n_433),
.B1(n_420),
.B2(n_429),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_401),
.C(n_382),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_454),
.C(n_455),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_377),
.C(n_381),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_366),
.C(n_398),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_426),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_293),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_421),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_467),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_469),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_456),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_466),
.B(n_468),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_432),
.Y(n_468)
);

XNOR2x1_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_418),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_472),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_425),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_424),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_474),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_442),
.A2(n_420),
.B(n_427),
.Y(n_475)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_475),
.Y(n_482)
);

AO21x1_ASAP7_75t_L g477 ( 
.A1(n_458),
.A2(n_416),
.B(n_343),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_347),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_458),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_480),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_462),
.B(n_443),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_440),
.C(n_452),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_485),
.A2(n_349),
.B(n_359),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_471),
.A2(n_450),
.B1(n_444),
.B2(n_460),
.Y(n_486)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_477),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_491),
.Y(n_501)
);

AOI31xp33_ASAP7_75t_L g488 ( 
.A1(n_470),
.A2(n_453),
.A3(n_451),
.B(n_459),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_488),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_490),
.A2(n_467),
.B(n_476),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_349),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_333),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_473),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_479),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_SL g494 ( 
.A(n_485),
.B(n_453),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_495),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_489),
.B(n_476),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_500),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_461),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_483),
.C(n_479),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_482),
.A2(n_333),
.B(n_339),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_504),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_508),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_489),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_510),
.B(n_493),
.C(n_499),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_490),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_511),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_498),
.A2(n_486),
.B1(n_484),
.B2(n_277),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_501),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_516),
.Y(n_519)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_509),
.Y(n_517)
);

AO21x1_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_511),
.B(n_507),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_518),
.A2(n_520),
.B(n_515),
.Y(n_521)
);

NOR2x1_ASAP7_75t_SL g520 ( 
.A(n_514),
.B(n_506),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_521),
.A2(n_522),
.B(n_516),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_510),
.C(n_502),
.Y(n_522)
);

AOI322xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_496),
.A3(n_236),
.B1(n_235),
.B2(n_263),
.C1(n_253),
.C2(n_259),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_248),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_235),
.B(n_263),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_248),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_253),
.B(n_13),
.Y(n_528)
);


endmodule