module real_jpeg_4514_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_1),
.A2(n_42),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_42),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_1),
.A2(n_42),
.B1(n_83),
.B2(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_3),
.A2(n_54),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_3),
.A2(n_54),
.B1(n_368),
.B2(n_371),
.Y(n_367)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_5),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_5),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_5),
.Y(n_305)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_6),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_30),
.B1(n_96),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_30),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_7),
.B(n_90),
.Y(n_223)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_7),
.A2(n_247),
.B(n_250),
.C(n_254),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_7),
.B(n_72),
.C(n_161),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_7),
.B(n_118),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_7),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_7),
.B(n_48),
.Y(n_309)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_11),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_11),
.A2(n_104),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_11),
.A2(n_104),
.B1(n_261),
.B2(n_264),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_11),
.A2(n_28),
.B1(n_104),
.B2(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_348),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_214),
.B(n_346),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_182),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_15),
.B(n_182),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g380 ( 
.A(n_15),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_144),
.CI(n_153),
.CON(n_15),
.SN(n_15)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_16),
.B(n_144),
.C(n_153),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_78),
.B2(n_79),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_17),
.B(n_80),
.C(n_112),
.Y(n_377)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_19),
.B(n_46),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_20),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_21),
.A2(n_34),
.B(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_24),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_26),
.A2(n_35),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_26),
.B(n_35),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_29),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_30),
.A2(n_83),
.B(n_86),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_30),
.B(n_87),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_30),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_32),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_33),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_35),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_35),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_36),
.Y(n_303)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_39),
.B(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_44),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B(n_59),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_47),
.A2(n_150),
.B(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_47),
.B(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_48),
.B(n_60),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_48),
.B(n_260),
.Y(n_275)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_51),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_53),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_58),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_58),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_59),
.B(n_275),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_59),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_62),
.Y(n_272)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_66),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_66),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_69),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_112),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_100),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_82),
.B(n_106),
.Y(n_230)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_82),
.Y(n_363)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_90),
.B(n_101),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_90),
.B(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_90),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_90)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_91),
.Y(n_195)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_93),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_94),
.Y(n_211)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_95),
.Y(n_194)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_96),
.Y(n_254)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_100),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_106),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_106),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_111),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_130),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_113),
.B(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_114),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_115),
.Y(n_212)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_118),
.A2(n_131),
.B(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_118),
.B(n_208),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_118),
.A2(n_234),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_119),
.B(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_123),
.Y(n_249)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_130),
.B(n_236),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_141),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_131),
.B(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_132),
.B(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_141),
.Y(n_206)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_145),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_145),
.A2(n_152),
.B1(n_246),
.B2(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_145),
.B(n_149),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_145),
.A2(n_152),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_151),
.B(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_174),
.C(n_176),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_166),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_155),
.B(n_166),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_162),
.B(n_163),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_163),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_163),
.B(n_279),
.Y(n_308)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_167),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_181),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_213),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_183),
.B(n_213),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_186),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_203),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_187),
.B(n_203),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_189),
.B(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_191),
.Y(n_227)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_195),
.A3(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_194),
.Y(n_370)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_330),
.B(n_343),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_265),
.B(n_329),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_241),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_217),
.B(n_241),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_228),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_226),
.B2(n_227),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_220),
.B(n_226),
.C(n_228),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.C(n_224),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_225),
.B(n_296),
.Y(n_306)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_229),
.B(n_232),
.C(n_238),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_255),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_242),
.B(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_245),
.A2(n_255),
.B1(n_256),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_245),
.Y(n_326)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_246),
.Y(n_321)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_258),
.B(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx11_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_323),
.B(n_328),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_313),
.B(n_322),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_290),
.B(n_312),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_276),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_276),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_271),
.B1(n_274),
.B2(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_285),
.Y(n_276)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_297),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_288),
.C(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_299),
.B(n_311),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_294),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_307),
.B(n_310),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_316),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_319),
.C(n_320),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_339),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_333),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_336),
.C(n_337),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_339),
.A2(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_342),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_378),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_350),
.B(n_351),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_377),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_364),
.B2(n_365),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B(n_363),
.Y(n_360)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_374),
.B(n_376),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_366),
.B(n_374),
.Y(n_376)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);


endmodule