module fake_jpeg_2418_n_108 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_13),
.C(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_25),
.C(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.Y(n_39)
);

NOR2xp67_ASAP7_75t_R g50 ( 
.A(n_39),
.B(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_31),
.B1(n_28),
.B2(n_32),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_51),
.B(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_32),
.B(n_29),
.C(n_34),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_26),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_26),
.Y(n_58)
);

NOR2xp67_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_50),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_65),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_76),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_54),
.B(n_50),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_1),
.B(n_3),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_28),
.B1(n_36),
.B2(n_30),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_62),
.B1(n_30),
.B2(n_36),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_SL g87 ( 
.A1(n_83),
.A2(n_48),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

AO221x1_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.C(n_80),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_15),
.Y(n_93)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_94),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_84),
.B1(n_86),
.B2(n_91),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_95),
.B(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_100),
.C(n_93),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);

AOI221xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_74),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_4),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_74),
.C2(n_16),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_17),
.CI(n_18),
.CON(n_108),
.SN(n_108)
);


endmodule