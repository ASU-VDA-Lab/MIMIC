module real_jpeg_17967_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_419),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_0),
.B(n_420),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_1),
.Y(n_420)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_2),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g36 ( 
.A(n_3),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_3),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_3),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_3),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_3),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_3),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_23),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_42),
.Y(n_41)
);

NAND2x1_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_56),
.Y(n_55)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_4),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_4),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_4),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_4),
.B(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_5),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_6),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_6),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_7),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_7),
.Y(n_128)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_10),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_125),
.Y(n_124)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_10),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_10),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_10),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_10),
.B(n_75),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

BUFx4f_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_102),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_60),
.B(n_101),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_17),
.B(n_60),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_50),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.C(n_39),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_19),
.A2(n_20),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_20)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_21),
.A2(n_33),
.B1(n_41),
.B2(n_94),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_22),
.A2(n_41),
.B1(n_49),
.B2(n_94),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_22),
.A2(n_49),
.B1(n_137),
.B2(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_22),
.B(n_143),
.C(n_235),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_22),
.A2(n_93),
.B(n_98),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_22),
.A2(n_49),
.B1(n_235),
.B2(n_238),
.Y(n_304)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_26),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_26),
.A2(n_27),
.B1(n_243),
.B2(n_245),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_30),
.C(n_49),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_27),
.B(n_41),
.Y(n_98)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_30),
.A2(n_34),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_30),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_30),
.B(n_143),
.C(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_30),
.B(n_288),
.C(n_290),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_30),
.B(n_270),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_30),
.A2(n_34),
.B1(n_288),
.B2(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_30),
.A2(n_34),
.B1(n_74),
.B2(n_244),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_30),
.B(n_74),
.C(n_347),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_34),
.B(n_270),
.C(n_292),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.C(n_49),
.Y(n_40)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_R g199 ( 
.A1(n_41),
.A2(n_124),
.B(n_200),
.C(n_206),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_41),
.B(n_124),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_41),
.A2(n_94),
.B1(n_124),
.B2(n_130),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_41),
.B(n_95),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_41),
.B(n_74),
.C(n_96),
.Y(n_261)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_43),
.Y(n_136)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_43),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_43),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_45),
.B(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_45),
.A2(n_127),
.B(n_201),
.Y(n_324)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_49),
.B(n_133),
.C(n_137),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_55),
.A2(n_57),
.B1(n_157),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_55),
.B(n_129),
.C(n_157),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_55),
.A2(n_57),
.B1(n_126),
.B2(n_131),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_55),
.A2(n_57),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_55),
.B(n_113),
.C(n_127),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_57),
.B(n_143),
.C(n_336),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_86),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_61),
.B(n_64),
.Y(n_410)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.C(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_69),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_68),
.Y(n_237)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_69),
.A2(n_247),
.B(n_251),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_69),
.B(n_247),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_69),
.A2(n_91),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_69),
.B(n_95),
.C(n_114),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_138),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_70),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.C(n_81),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_74),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_74),
.A2(n_244),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_76),
.A2(n_95),
.B1(n_96),
.B2(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_76),
.A2(n_96),
.B(n_134),
.C(n_206),
.Y(n_230)
);

AO22x1_ASAP7_75t_L g318 ( 
.A1(n_76),
.A2(n_166),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_76),
.B(n_186),
.C(n_319),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_166),
.Y(n_385)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_80),
.Y(n_341)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_86),
.B(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_87),
.A2(n_88),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_92),
.B(n_99),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B(n_98),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_95),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_95),
.B(n_213),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_95),
.A2(n_96),
.B1(n_113),
.B2(n_114),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_97),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_374),
.B(n_411),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI321xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_282),
.A3(n_362),
.B1(n_367),
.B2(n_368),
.C(n_373),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_254),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_223),
.B(n_253),
.Y(n_106)
);

AOI21x1_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_178),
.B(n_222),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_152),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_109),
.B(n_152),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_132),
.C(n_141),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_123),
.Y(n_110)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_111),
.Y(n_214)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_112),
.A2(n_124),
.B(n_131),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_113),
.A2(n_114),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_127),
.B(n_129),
.Y(n_126)
);

NAND2x1p5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_127),
.Y(n_129)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_117),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_118),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_127),
.A2(n_189),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_127),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_127),
.B(n_201),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_127),
.A2(n_195),
.B1(n_201),
.B2(n_204),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_132),
.A2(n_141),
.B1(n_142),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_134),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_134),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_137),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_137),
.A2(n_157),
.B1(n_160),
.B2(n_186),
.Y(n_262)
);

XNOR2x2_ASAP7_75t_L g317 ( 
.A(n_137),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_151),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_143),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_143),
.A2(n_151),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_148),
.A2(n_171),
.B1(n_234),
.B2(n_239),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_151),
.B(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_163),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_161),
.B2(n_162),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_161),
.C(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_160),
.B(n_186),
.C(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_164),
.B(n_169),
.C(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_171),
.B(n_201),
.C(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_174),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_174),
.A2(n_177),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_174),
.B(n_271),
.C(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_188),
.B(n_189),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_197),
.B(n_221),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_183),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_193),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_193),
.B1(n_194),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_189),
.Y(n_196)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_210),
.B(n_220),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_207),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_204),
.B1(n_235),
.B2(n_238),
.Y(n_234)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_217),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_216),
.B(n_219),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_214),
.B(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_225),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_240),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_228),
.C(n_240),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_233),
.C(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_232),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_252),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_246),
.C(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_251),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_255),
.B(n_256),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_267),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_257),
.B(n_268),
.C(n_281),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_281),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_277),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_279),
.C(n_280),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_350),
.Y(n_282)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_283),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_325),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_284),
.B(n_325),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_305),
.C(n_313),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_285),
.B(n_314),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_298),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_291),
.B1(n_296),
.B2(n_297),
.Y(n_286)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_297),
.C(n_298),
.Y(n_326)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_291),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_302),
.C(n_303),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_299),
.A2(n_300),
.B1(n_302),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

XOR2x2_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_305),
.B(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.C(n_309),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_308),
.Y(n_357)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_315),
.B(n_317),
.C(n_323),
.Y(n_344)
);

XOR2x1_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_328),
.C(n_343),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_343),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_333),
.C(n_342),
.Y(n_387)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_342),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_346),
.C(n_349),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

AOI31xp67_ASAP7_75t_L g368 ( 
.A1(n_350),
.A2(n_363),
.A3(n_369),
.B(n_372),
.Y(n_368)
);

NAND2x1p5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NOR2x1_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_353),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_358),
.C(n_359),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_359),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_366),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NOR3xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_395),
.C(n_406),
.Y(n_375)
);

AND2x4_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_378),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_381),
.C(n_388),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_388),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_386),
.C(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_387),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_391),
.B1(n_392),
.B2(n_393),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_390),
.B(n_393),
.C(n_394),
.Y(n_404)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_396),
.A2(n_414),
.B(n_415),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_405),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_405),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_398),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_404),
.C(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_406),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_409),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_416),
.B(n_417),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);


endmodule