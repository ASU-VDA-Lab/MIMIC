module fake_jpeg_28736_n_355 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_43),
.Y(n_90)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_52),
.Y(n_81)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_58),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_62),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

OR2x4_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_12),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_11),
.Y(n_87)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_22),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_69),
.B(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_71),
.Y(n_123)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_35),
.B1(n_41),
.B2(n_37),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_76),
.A2(n_77),
.B1(n_85),
.B2(n_109),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_35),
.B1(n_41),
.B2(n_37),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_35),
.B1(n_32),
.B2(n_37),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_80),
.A2(n_86),
.B1(n_124),
.B2(n_42),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_38),
.B1(n_30),
.B2(n_37),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_82),
.A2(n_101),
.B1(n_56),
.B2(n_46),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_29),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_94),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_41),
.B1(n_32),
.B2(n_39),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_21),
.B1(n_36),
.B2(n_33),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_43),
.B(n_40),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_50),
.A2(n_30),
.B1(n_38),
.B2(n_23),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_59),
.B(n_18),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_114),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_60),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_48),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_40),
.B1(n_39),
.B2(n_31),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_62),
.A2(n_36),
.B1(n_33),
.B2(n_25),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_25),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_118),
.B(n_114),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_49),
.A2(n_23),
.B1(n_24),
.B2(n_10),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_51),
.B(n_24),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_24),
.B1(n_23),
.B2(n_3),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_125),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_162),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_10),
.C(n_58),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_143),
.Y(n_170)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_78),
.A2(n_54),
.B(n_44),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_121),
.C(n_95),
.Y(n_183)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_67),
.B1(n_66),
.B2(n_55),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_152),
.B1(n_123),
.B2(n_119),
.Y(n_172)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_81),
.B(n_48),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_112),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_153),
.A2(n_159),
.B1(n_124),
.B2(n_104),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_84),
.A2(n_48),
.B(n_43),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_90),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_157),
.Y(n_186)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_79),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_160),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_78),
.A2(n_119),
.B1(n_123),
.B2(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_94),
.B(n_43),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_88),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_96),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_164),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_106),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_129),
.B(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_169),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_117),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_86),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_180),
.B1(n_131),
.B2(n_146),
.Y(n_202)
);

AND2x4_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_153),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_91),
.B1(n_113),
.B2(n_121),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_167),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_88),
.B(n_95),
.C(n_91),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_132),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_134),
.A2(n_89),
.B1(n_105),
.B2(n_92),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_197),
.B1(n_141),
.B2(n_122),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_150),
.B(n_111),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_2),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_111),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_176),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_122),
.B1(n_90),
.B2(n_3),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_210),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_199),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_142),
.B1(n_137),
.B2(n_130),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_218),
.Y(n_233)
);

HB1xp67_ASAP7_75t_SL g231 ( 
.A(n_201),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_144),
.B1(n_161),
.B2(n_140),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_126),
.B1(n_156),
.B2(n_145),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_136),
.B1(n_147),
.B2(n_157),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_138),
.B1(n_125),
.B2(n_133),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_151),
.B1(n_2),
.B2(n_3),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_230),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_151),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_184),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_215),
.A2(n_182),
.B1(n_179),
.B2(n_190),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_190),
.B1(n_179),
.B2(n_182),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_187),
.A2(n_7),
.B1(n_9),
.B2(n_180),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_9),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_170),
.B(n_187),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_167),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g229 ( 
.A1(n_183),
.A2(n_164),
.B1(n_163),
.B2(n_185),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_175),
.B(n_169),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_171),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_209),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_254),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_249),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_202),
.B1(n_221),
.B2(n_207),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_171),
.B1(n_224),
.B2(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_182),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_186),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_252),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_195),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_197),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_199),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_222),
.B(n_195),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_199),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_216),
.C(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_263),
.C(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_208),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_214),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_229),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_239),
.B(n_200),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_265),
.B(n_246),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_201),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_249),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_251),
.B1(n_233),
.B2(n_247),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_SL g270 ( 
.A(n_237),
.B(n_201),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_279),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_209),
.C(n_201),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_278),
.C(n_252),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_206),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_243),
.B(n_225),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_277),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_276),
.B1(n_204),
.B2(n_235),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_233),
.A2(n_205),
.B1(n_219),
.B2(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_210),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_284),
.B(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_275),
.A2(n_246),
.B1(n_235),
.B2(n_251),
.Y(n_286)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_297),
.B1(n_260),
.B2(n_278),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_236),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_257),
.C(n_263),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_236),
.C(n_254),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_271),
.C(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_251),
.B1(n_256),
.B2(n_255),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_302),
.B1(n_311),
.B2(n_309),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_264),
.B1(n_258),
.B2(n_277),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_289),
.Y(n_318)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_304),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_310),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_270),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_295),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_308),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_258),
.C(n_241),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_309),
.A2(n_242),
.B(n_240),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_255),
.C(n_240),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_294),
.A2(n_289),
.B(n_296),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_281),
.B(n_291),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_317),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_238),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_307),
.B1(n_245),
.B2(n_224),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_319),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_298),
.A2(n_295),
.B1(n_281),
.B2(n_238),
.Y(n_319)
);

AND2x2_ASAP7_75t_SL g334 ( 
.A(n_320),
.B(n_322),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_242),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_320),
.B(n_314),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_319),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_313),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_324),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_335),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_312),
.B(n_323),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_333),
.A2(n_322),
.B(n_303),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_318),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_337),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_339),
.B(n_342),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_328),
.B(n_300),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_310),
.C(n_300),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_334),
.C(n_321),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_343),
.A2(n_346),
.B(n_189),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_341),
.B(n_213),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_321),
.A3(n_334),
.B1(n_338),
.B2(n_342),
.C1(n_196),
.C2(n_336),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_181),
.B1(n_345),
.B2(n_196),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_349),
.A2(n_350),
.B(n_346),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_344),
.A2(n_184),
.B(n_181),
.C(n_218),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_352),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_174),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_354),
.B(n_174),
.Y(n_355)
);


endmodule