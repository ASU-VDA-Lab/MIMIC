module fake_netlist_5_1314_n_1130 (n_137, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1130);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1130;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_1126;
wire n_642;
wire n_469;
wire n_615;
wire n_1060;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_1099;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_983;
wire n_1128;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_1112;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_1120;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_1110;
wire n_951;
wire n_1121;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_368;
wire n_247;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_1048;
wire n_946;
wire n_612;
wire n_1001;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_1118;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_1063;
wire n_556;
wire n_1107;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_1124;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_1104;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_1049;
wire n_938;
wire n_1098;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_1108;
wire n_325;
wire n_449;
wire n_1073;
wire n_1100;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_1096;
wire n_976;
wire n_1095;
wire n_234;
wire n_343;
wire n_428;
wire n_308;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_223;
wire n_1114;
wire n_1129;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_1097;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_1020;
wire n_215;
wire n_350;
wire n_798;
wire n_662;
wire n_459;
wire n_1062;
wire n_646;
wire n_897;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_1119;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_1069;
wire n_1075;
wire n_388;
wire n_1127;
wire n_761;
wire n_1012;
wire n_1019;
wire n_1105;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_571;
wire n_477;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_1113;
wire n_652;
wire n_778;
wire n_1111;
wire n_1122;
wire n_306;
wire n_907;
wire n_722;
wire n_1093;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_989;
wire n_852;
wire n_1041;
wire n_1039;
wire n_1102;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_893;
wire n_502;
wire n_892;
wire n_736;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_846;
wire n_586;
wire n_1058;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_748;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_1101;
wire n_273;
wire n_585;
wire n_349;
wire n_1106;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1116;
wire n_767;
wire n_217;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_1103;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_679;
wire n_795;
wire n_695;
wire n_857;
wire n_832;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_1094;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_233;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_1125;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_1109;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_1038;
wire n_409;
wire n_797;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_931;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_870;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_1092;
wire n_238;
wire n_1117;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_890;
wire n_1032;
wire n_764;
wire n_960;
wire n_1056;
wire n_759;
wire n_1018;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_1123;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_12),
.Y(n_209)
);

CKINVDCx11_ASAP7_75t_R g210 ( 
.A(n_144),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_170),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_95),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_62),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_132),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_68),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_131),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_171),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_118),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_117),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_111),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_30),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_197),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_108),
.Y(n_230)
);

CKINVDCx12_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_79),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_125),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_60),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_110),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_35),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_82),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_159),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_156),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_53),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_41),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_172),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_148),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_208),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_21),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_193),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_161),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_2),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_177),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_194),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_198),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_102),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_185),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_23),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_124),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_17),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_89),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_154),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_99),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_50),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_136),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_98),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_3),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_81),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_31),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_73),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_75),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_191),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_47),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_162),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_17),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_123),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_188),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_19),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_174),
.Y(n_281)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_269),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_218),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_210),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_213),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_223),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_210),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_239),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_230),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_218),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_241),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVxp33_ASAP7_75t_SL g310 ( 
.A(n_259),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_221),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_280),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_239),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_209),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_239),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_211),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_0),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_219),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_282),
.A2(n_237),
.B1(n_246),
.B2(n_242),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_214),
.B(n_212),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_278),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_323),
.A2(n_217),
.B(n_216),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_220),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_316),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_298),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_282),
.A2(n_251),
.B1(n_227),
.B2(n_231),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_219),
.Y(n_341)
);

AND2x6_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_219),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_263),
.Y(n_343)
);

BUFx12f_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_294),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_279),
.Y(n_353)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_327),
.A2(n_225),
.B(n_222),
.Y(n_354)
);

AND2x2_ASAP7_75t_R g355 ( 
.A(n_297),
.B(n_263),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_294),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_263),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_283),
.A2(n_276),
.B1(n_275),
.B2(n_273),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_302),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_329),
.B(n_304),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_321),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_228),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_303),
.B(n_232),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_234),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_289),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_307),
.B(n_267),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_289),
.Y(n_371)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_285),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_308),
.B(n_235),
.Y(n_373)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_290),
.A2(n_240),
.B(n_236),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_309),
.B(n_265),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_284),
.Y(n_376)
);

BUFx12f_ASAP7_75t_L g377 ( 
.A(n_297),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_311),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_290),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_320),
.Y(n_380)
);

INVx5_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_313),
.B(n_243),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_292),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_330),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_331),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_331),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_344),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_320),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_344),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_377),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_339),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_R g399 ( 
.A(n_338),
.B(n_380),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_377),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_380),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_372),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_364),
.B(n_314),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_360),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_337),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_353),
.B(n_312),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_341),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_343),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_340),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_368),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_372),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_334),
.B(n_293),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_372),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_R g418 ( 
.A(n_374),
.B(n_244),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_370),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_373),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_375),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_362),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_359),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_R g425 ( 
.A(n_359),
.B(n_291),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_362),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_364),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_334),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_374),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_345),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_364),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_306),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_367),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_367),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_367),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_382),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_355),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_382),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_382),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_358),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_342),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_342),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_365),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_345),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_342),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_374),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_365),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_342),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_348),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_342),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_348),
.Y(n_456)
);

BUFx6f_ASAP7_75t_SL g457 ( 
.A(n_342),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_371),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_301),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_387),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_434),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_286),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_405),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_419),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_317),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_333),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_333),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_L g473 ( 
.A(n_420),
.B(n_421),
.Y(n_473)
);

BUFx4f_ASAP7_75t_L g474 ( 
.A(n_395),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_318),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_398),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_R g477 ( 
.A(n_399),
.B(n_247),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_403),
.B(n_408),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_445),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_430),
.A2(n_333),
.B1(n_336),
.B2(n_354),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_450),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_422),
.B(n_336),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_417),
.B(n_248),
.Y(n_483)
);

AND2x6_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_319),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_413),
.B(n_336),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_410),
.B(n_322),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_398),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_354),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g490 ( 
.A(n_425),
.B(n_250),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_416),
.B(n_354),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_371),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_428),
.B(n_432),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_371),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_430),
.A2(n_295),
.B1(n_296),
.B2(n_315),
.Y(n_495)
);

BUFx6f_ASAP7_75t_SL g496 ( 
.A(n_388),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_366),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_431),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_431),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_391),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_411),
.B(n_254),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_396),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_448),
.B(n_366),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_392),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_391),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_426),
.B(n_295),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_385),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

AND2x2_ASAP7_75t_SL g512 ( 
.A(n_412),
.B(n_296),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_385),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_443),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_385),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_451),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_451),
.B(n_366),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_435),
.B(n_255),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_436),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_437),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_402),
.B(n_0),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_438),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_406),
.B(n_256),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_418),
.A2(n_257),
.B1(n_258),
.B2(n_261),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_388),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_440),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_392),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_441),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_386),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_389),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_390),
.B(n_365),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_423),
.B(n_365),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_433),
.B(n_389),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_423),
.B(n_444),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_394),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_397),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_457),
.B(n_346),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_449),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_453),
.B(n_455),
.C(n_369),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_457),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_400),
.B(n_379),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_498),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_507),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_476),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_475),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g548 ( 
.A(n_501),
.B(n_346),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_501),
.B(n_347),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_495),
.B(n_379),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_467),
.B(n_36),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_464),
.Y(n_552)
);

OR2x2_ASAP7_75t_SL g553 ( 
.A(n_522),
.B(n_1),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_495),
.B(n_379),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_489),
.B(n_482),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_504),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_489),
.B(n_379),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_476),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_460),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_502),
.B(n_508),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_482),
.B(n_366),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_471),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_533),
.B(n_366),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_488),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_466),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_478),
.B(n_37),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_492),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_486),
.B(n_383),
.C(n_369),
.Y(n_569)
);

NOR3xp33_ASAP7_75t_L g570 ( 
.A(n_473),
.B(n_352),
.C(n_347),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_542),
.B(n_457),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_485),
.B(n_369),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_503),
.B(n_524),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_500),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_502),
.B(n_369),
.Y(n_576)
);

NAND2x1p5_ASAP7_75t_L g577 ( 
.A(n_508),
.B(n_369),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_463),
.B(n_383),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_496),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_513),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_469),
.A2(n_383),
.B1(n_352),
.B2(n_381),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_504),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_485),
.B(n_383),
.Y(n_584)
);

OR2x6_ASAP7_75t_L g585 ( 
.A(n_529),
.B(n_383),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_461),
.B(n_351),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_494),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_459),
.B(n_1),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_528),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_468),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_478),
.B(n_38),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_484),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_517),
.A2(n_381),
.B1(n_356),
.B2(n_330),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_511),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_506),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_514),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_513),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_516),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_474),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_497),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_518),
.A2(n_381),
.B1(n_356),
.B2(n_330),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_470),
.A2(n_381),
.B1(n_356),
.B2(n_330),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_487),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_497),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_543),
.B(n_2),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_467),
.B(n_3),
.Y(n_609)
);

AO22x2_ASAP7_75t_L g610 ( 
.A1(n_491),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_515),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_573),
.B(n_469),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_571),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_562),
.A2(n_575),
.B1(n_580),
.B2(n_568),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_562),
.A2(n_469),
.B1(n_535),
.B2(n_512),
.Y(n_615)
);

CKINVDCx10_ASAP7_75t_R g616 ( 
.A(n_579),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_589),
.A2(n_518),
.B1(n_472),
.B2(n_470),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_607),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_578),
.B(n_469),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_555),
.A2(n_542),
.B(n_472),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_590),
.A2(n_519),
.B(n_483),
.C(n_520),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_L g622 ( 
.A(n_571),
.B(n_538),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_585),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_547),
.B(n_474),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_547),
.A2(n_532),
.B1(n_525),
.B2(n_484),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_555),
.A2(n_541),
.B(n_540),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_564),
.B(n_461),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_583),
.B(n_461),
.Y(n_628)
);

AOI21xp33_ASAP7_75t_L g629 ( 
.A1(n_583),
.A2(n_525),
.B(n_527),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_567),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_557),
.A2(n_541),
.B(n_499),
.Y(n_631)
);

BUFx12f_ASAP7_75t_L g632 ( 
.A(n_602),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_567),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_557),
.A2(n_499),
.B(n_487),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_594),
.A2(n_484),
.B1(n_521),
.B2(n_523),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_561),
.A2(n_499),
.B(n_487),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_546),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_561),
.A2(n_505),
.B(n_480),
.Y(n_639)
);

NOR2x1_ASAP7_75t_L g640 ( 
.A(n_551),
.B(n_530),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_550),
.A2(n_480),
.B1(n_462),
.B2(n_493),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_566),
.B(n_462),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_556),
.B(n_493),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_572),
.A2(n_505),
.B(n_539),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_572),
.A2(n_539),
.B(n_356),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_556),
.B(n_529),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_584),
.A2(n_539),
.B(n_356),
.Y(n_647)
);

A2O1A1Ixp33_ASAP7_75t_L g648 ( 
.A1(n_608),
.A2(n_490),
.B(n_529),
.C(n_537),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_587),
.B(n_484),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_584),
.A2(n_465),
.B(n_539),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_544),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_593),
.B(n_477),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_594),
.A2(n_534),
.B(n_465),
.C(n_6),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_550),
.A2(n_531),
.B(n_526),
.C(n_536),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_554),
.A2(n_465),
.B(n_534),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_606),
.A2(n_330),
.B(n_351),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_593),
.B(n_534),
.Y(n_657)
);

NAND2x1p5_ASAP7_75t_L g658 ( 
.A(n_591),
.B(n_351),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_558),
.Y(n_659)
);

O2A1O1Ixp5_ASAP7_75t_L g660 ( 
.A1(n_586),
.A2(n_465),
.B(n_96),
.C(n_207),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_600),
.B(n_592),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_606),
.A2(n_357),
.B(n_351),
.Y(n_662)
);

BUFx4f_ASAP7_75t_L g663 ( 
.A(n_585),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_588),
.B(n_4),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_554),
.A2(n_357),
.B(n_40),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_596),
.B(n_5),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_559),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_597),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_560),
.A2(n_549),
.B(n_548),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_545),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_609),
.A2(n_496),
.B1(n_357),
.B2(n_97),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_585),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_560),
.A2(n_357),
.B(n_42),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_615),
.B(n_598),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_620),
.A2(n_569),
.B(n_604),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_639),
.A2(n_549),
.B(n_548),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_627),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_618),
.B(n_563),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_626),
.A2(n_605),
.B(n_611),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_SL g680 ( 
.A(n_621),
.B(n_570),
.C(n_553),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_643),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_668),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_SL g683 ( 
.A(n_654),
.B(n_610),
.C(n_570),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_617),
.B(n_612),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_634),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_629),
.B(n_599),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_625),
.A2(n_565),
.B(n_574),
.C(n_601),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_661),
.B(n_581),
.Y(n_688)
);

AO32x2_ASAP7_75t_L g689 ( 
.A1(n_641),
.A2(n_610),
.A3(n_595),
.B1(n_577),
.B2(n_576),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_652),
.B(n_581),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_SL g691 ( 
.A(n_648),
.B(n_610),
.C(n_7),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_651),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_614),
.B(n_576),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_613),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_616),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_622),
.A2(n_577),
.B(n_582),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_646),
.B(n_7),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_655),
.A2(n_571),
.B(n_9),
.C(n_10),
.Y(n_698)
);

AOI222xp33_ASAP7_75t_L g699 ( 
.A1(n_657),
.A2(n_571),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_632),
.Y(n_700)
);

AO32x1_ASAP7_75t_L g701 ( 
.A1(n_670),
.A2(n_8),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_624),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_636),
.A2(n_571),
.B(n_13),
.C(n_14),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_SL g704 ( 
.A(n_671),
.B(n_8),
.C(n_15),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_642),
.B(n_16),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_630),
.B(n_16),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_667),
.Y(n_707)
);

O2A1O1Ixp5_ASAP7_75t_L g708 ( 
.A1(n_650),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_630),
.B(n_18),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_638),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_663),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_669),
.A2(n_43),
.B(n_39),
.Y(n_712)
);

O2A1O1Ixp5_ASAP7_75t_L g713 ( 
.A1(n_645),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_713)
);

AOI21x1_ASAP7_75t_L g714 ( 
.A1(n_631),
.A2(n_205),
.B(n_112),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_630),
.B(n_25),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_633),
.B(n_25),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_619),
.A2(n_113),
.B(n_203),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_666),
.A2(n_649),
.B(n_628),
.C(n_664),
.Y(n_718)
);

AOI21x1_ASAP7_75t_L g719 ( 
.A1(n_644),
.A2(n_109),
.B(n_202),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_633),
.B(n_26),
.Y(n_720)
);

CKINVDCx16_ASAP7_75t_R g721 ( 
.A(n_633),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_653),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_659),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_635),
.A2(n_107),
.B(n_201),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_658),
.B(n_27),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_640),
.B(n_28),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_623),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_672),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_672),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_672),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_613),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_665),
.A2(n_204),
.B(n_115),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_660),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_692),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_685),
.Y(n_735)
);

BUFx4f_ASAP7_75t_SL g736 ( 
.A(n_700),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_681),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_729),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_729),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_702),
.Y(n_741)
);

AO21x1_ASAP7_75t_L g742 ( 
.A1(n_674),
.A2(n_647),
.B(n_637),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_707),
.Y(n_743)
);

INVx6_ASAP7_75t_L g744 ( 
.A(n_721),
.Y(n_744)
);

BUFx12f_ASAP7_75t_L g745 ( 
.A(n_695),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_694),
.B(n_613),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_694),
.B(n_673),
.Y(n_747)
);

INVx8_ASAP7_75t_L g748 ( 
.A(n_731),
.Y(n_748)
);

BUFx2_ASAP7_75t_SL g749 ( 
.A(n_681),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_731),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_723),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_727),
.Y(n_752)
);

BUFx2_ASAP7_75t_SL g753 ( 
.A(n_706),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_697),
.B(n_29),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_682),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_690),
.B(n_656),
.Y(n_756)
);

BUFx12f_ASAP7_75t_L g757 ( 
.A(n_725),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_710),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_728),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_709),
.Y(n_760)
);

CKINVDCx14_ASAP7_75t_R g761 ( 
.A(n_720),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_716),
.Y(n_762)
);

CKINVDCx16_ASAP7_75t_R g763 ( 
.A(n_680),
.Y(n_763)
);

BUFx12f_ASAP7_75t_L g764 ( 
.A(n_715),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_693),
.B(n_662),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_714),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_678),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_677),
.Y(n_768)
);

INVx5_ASAP7_75t_L g769 ( 
.A(n_733),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_704),
.B(n_44),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_688),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_683),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_719),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_675),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_686),
.B(n_32),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_726),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_691),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_705),
.Y(n_778)
);

INVx3_ASAP7_75t_SL g779 ( 
.A(n_699),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_684),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_699),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_687),
.Y(n_782)
);

INVx3_ASAP7_75t_SL g783 ( 
.A(n_698),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_718),
.B(n_33),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_722),
.B(n_703),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_730),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_711),
.Y(n_787)
);

INVx3_ASAP7_75t_SL g788 ( 
.A(n_708),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_689),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_689),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_717),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_712),
.Y(n_792)
);

BUFx2_ASAP7_75t_SL g793 ( 
.A(n_724),
.Y(n_793)
);

NAND2x1p5_ASAP7_75t_L g794 ( 
.A(n_676),
.B(n_45),
.Y(n_794)
);

BUFx2_ASAP7_75t_SL g795 ( 
.A(n_696),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_732),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_689),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_732),
.B(n_46),
.Y(n_798)
);

OAI21x1_ASAP7_75t_SL g799 ( 
.A1(n_785),
.A2(n_679),
.B(n_701),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_779),
.A2(n_713),
.B1(n_701),
.B2(n_34),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_735),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_784),
.A2(n_701),
.B(n_49),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_784),
.A2(n_48),
.B(n_51),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_735),
.B(n_52),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_737),
.Y(n_805)
);

AOI21x1_ASAP7_75t_L g806 ( 
.A1(n_782),
.A2(n_54),
.B(n_55),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_737),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_754),
.B(n_56),
.Y(n_808)
);

OAI21x1_ASAP7_75t_L g809 ( 
.A1(n_766),
.A2(n_57),
.B(n_58),
.Y(n_809)
);

INVx6_ASAP7_75t_L g810 ( 
.A(n_744),
.Y(n_810)
);

AO21x2_ASAP7_75t_L g811 ( 
.A1(n_773),
.A2(n_59),
.B(n_61),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_774),
.Y(n_812)
);

BUFx4_ASAP7_75t_SL g813 ( 
.A(n_741),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_766),
.A2(n_63),
.B(n_64),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_745),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_773),
.A2(n_65),
.B(n_66),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_741),
.Y(n_817)
);

OAI21x1_ASAP7_75t_SL g818 ( 
.A1(n_781),
.A2(n_67),
.B(n_69),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_769),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_744),
.Y(n_820)
);

AOI21x1_ASAP7_75t_L g821 ( 
.A1(n_772),
.A2(n_70),
.B(n_71),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_794),
.A2(n_72),
.B(n_74),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_743),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_781),
.A2(n_199),
.B1(n_77),
.B2(n_78),
.Y(n_824)
);

OA21x2_ASAP7_75t_L g825 ( 
.A1(n_742),
.A2(n_76),
.B(n_80),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_737),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_743),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_774),
.Y(n_828)
);

OA21x2_ASAP7_75t_L g829 ( 
.A1(n_797),
.A2(n_83),
.B(n_84),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_760),
.B(n_85),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_795),
.B(n_86),
.Y(n_831)
);

OAI21x1_ASAP7_75t_L g832 ( 
.A1(n_794),
.A2(n_87),
.B(n_88),
.Y(n_832)
);

BUFx8_ASAP7_75t_L g833 ( 
.A(n_745),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_767),
.B(n_90),
.Y(n_834)
);

AOI21x1_ASAP7_75t_L g835 ( 
.A1(n_775),
.A2(n_91),
.B(n_92),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_750),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_765),
.A2(n_93),
.B(n_94),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_763),
.B(n_778),
.Y(n_838)
);

OR2x6_ASAP7_75t_SL g839 ( 
.A(n_792),
.B(n_100),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_780),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_770),
.A2(n_101),
.B(n_103),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_744),
.Y(n_842)
);

BUFx2_ASAP7_75t_SL g843 ( 
.A(n_739),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_780),
.A2(n_104),
.B(n_105),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_787),
.A2(n_106),
.B1(n_114),
.B2(n_119),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_776),
.B(n_120),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_738),
.B(n_121),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_751),
.B(n_126),
.Y(n_848)
);

AO21x2_ASAP7_75t_L g849 ( 
.A1(n_798),
.A2(n_127),
.B(n_128),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_737),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_765),
.A2(n_129),
.B(n_130),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_747),
.A2(n_133),
.B(n_134),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_777),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_853)
);

OA21x2_ASAP7_75t_L g854 ( 
.A1(n_802),
.A2(n_791),
.B(n_798),
.Y(n_854)
);

OAI22xp33_ASAP7_75t_L g855 ( 
.A1(n_839),
.A2(n_777),
.B1(n_783),
.B2(n_787),
.Y(n_855)
);

NOR2x1_ASAP7_75t_SL g856 ( 
.A(n_831),
.B(n_769),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_801),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_819),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_823),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_812),
.B(n_789),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_827),
.Y(n_861)
);

CKINVDCx8_ASAP7_75t_R g862 ( 
.A(n_843),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_819),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_840),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_840),
.B(n_738),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_812),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_838),
.B(n_768),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_829),
.B(n_789),
.Y(n_868)
);

BUFx4f_ASAP7_75t_L g869 ( 
.A(n_829),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_828),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_829),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_799),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_825),
.B(n_789),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_825),
.Y(n_874)
);

AOI21x1_ASAP7_75t_L g875 ( 
.A1(n_800),
.A2(n_751),
.B(n_734),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_811),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_842),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_847),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_825),
.B(n_769),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_836),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_805),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_816),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_816),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_811),
.Y(n_884)
);

INVxp67_ASAP7_75t_SL g885 ( 
.A(n_834),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_836),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_809),
.A2(n_796),
.B(n_747),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_824),
.A2(n_783),
.B1(n_786),
.B2(n_777),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_820),
.B(n_789),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_844),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_833),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_805),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_820),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_804),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_804),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_803),
.A2(n_758),
.B(n_788),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_804),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_831),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_848),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_855),
.A2(n_824),
.B1(n_796),
.B2(n_777),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_867),
.B(n_893),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_857),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_864),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_860),
.B(n_790),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_869),
.B(n_898),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_864),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_878),
.B(n_778),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_889),
.B(n_817),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_858),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_865),
.B(n_771),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_889),
.B(n_817),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_R g912 ( 
.A(n_896),
.B(n_831),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_891),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_885),
.B(n_771),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_888),
.A2(n_786),
.B1(n_818),
.B2(n_841),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_859),
.B(n_762),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_860),
.B(n_790),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_R g918 ( 
.A(n_896),
.B(n_868),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_863),
.B(n_761),
.Y(n_919)
);

CKINVDCx16_ASAP7_75t_R g920 ( 
.A(n_891),
.Y(n_920)
);

INVxp33_ASAP7_75t_SL g921 ( 
.A(n_880),
.Y(n_921)
);

CKINVDCx8_ASAP7_75t_R g922 ( 
.A(n_892),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_854),
.A2(n_761),
.B1(n_788),
.B2(n_845),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_864),
.B(n_790),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_861),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_869),
.A2(n_845),
.B1(n_853),
.B2(n_753),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_866),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_887),
.A2(n_806),
.B(n_814),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_872),
.Y(n_929)
);

INVxp67_ASAP7_75t_SL g930 ( 
.A(n_871),
.Y(n_930)
);

CKINVDCx11_ASAP7_75t_R g931 ( 
.A(n_862),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_866),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_901),
.B(n_868),
.Y(n_933)
);

AO21x2_ASAP7_75t_L g934 ( 
.A1(n_930),
.A2(n_874),
.B(n_876),
.Y(n_934)
);

OAI221xp5_ASAP7_75t_SL g935 ( 
.A1(n_923),
.A2(n_853),
.B1(n_846),
.B2(n_868),
.C(n_830),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_908),
.B(n_868),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_909),
.B(n_873),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_900),
.A2(n_869),
.B(n_846),
.C(n_873),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_914),
.B(n_899),
.Y(n_939)
);

INVx4_ASAP7_75t_R g940 ( 
.A(n_931),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_930),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_927),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_926),
.A2(n_854),
.B1(n_896),
.B2(n_849),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_932),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_902),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_903),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_909),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_911),
.B(n_917),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_906),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_925),
.Y(n_950)
);

AO21x2_ASAP7_75t_L g951 ( 
.A1(n_928),
.A2(n_876),
.B(n_890),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_929),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_929),
.A2(n_890),
.B(n_884),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_904),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_924),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_905),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_938),
.A2(n_923),
.B(n_915),
.C(n_913),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_940),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_940),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_935),
.A2(n_856),
.B(n_915),
.Y(n_960)
);

AO31x2_ASAP7_75t_L g961 ( 
.A1(n_941),
.A2(n_952),
.A3(n_856),
.B(n_950),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_943),
.A2(n_849),
.B(n_898),
.Y(n_962)
);

OAI211xp5_ASAP7_75t_L g963 ( 
.A1(n_943),
.A2(n_931),
.B(n_907),
.C(n_916),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_947),
.A2(n_910),
.B(n_877),
.C(n_919),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_956),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_933),
.B(n_905),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_939),
.B(n_921),
.Y(n_967)
);

AO31x2_ASAP7_75t_L g968 ( 
.A1(n_941),
.A2(n_898),
.A3(n_892),
.B(n_884),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_952),
.A2(n_755),
.B(n_879),
.C(n_886),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_933),
.B(n_917),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_950),
.Y(n_971)
);

AO31x2_ASAP7_75t_L g972 ( 
.A1(n_950),
.A2(n_882),
.A3(n_883),
.B(n_870),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_959),
.B(n_920),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_958),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_971),
.Y(n_975)
);

AO21x2_ASAP7_75t_L g976 ( 
.A1(n_962),
.A2(n_934),
.B(n_953),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_968),
.Y(n_977)
);

AND2x2_ASAP7_75t_SL g978 ( 
.A(n_957),
.B(n_854),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_968),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_967),
.B(n_954),
.Y(n_980)
);

AOI21xp33_ASAP7_75t_SL g981 ( 
.A1(n_963),
.A2(n_815),
.B(n_918),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_961),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_966),
.B(n_936),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_968),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_975),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_974),
.B(n_970),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_980),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_976),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_977),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_983),
.B(n_954),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_973),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_981),
.B(n_937),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_986),
.Y(n_993)
);

NOR2x1_ASAP7_75t_L g994 ( 
.A(n_991),
.B(n_973),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_991),
.B(n_815),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_992),
.B(n_978),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_989),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_987),
.B(n_978),
.Y(n_998)
);

NAND2x1_ASAP7_75t_SL g999 ( 
.A(n_988),
.B(n_977),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_993),
.B(n_998),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_994),
.B(n_985),
.Y(n_1001)
);

AND5x1_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_960),
.C(n_964),
.D(n_969),
.E(n_976),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_996),
.B(n_833),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_997),
.A2(n_988),
.B1(n_990),
.B2(n_956),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_937),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_997),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_993),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_993),
.B(n_961),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_993),
.B(n_945),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_993),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_1007),
.A2(n_982),
.B1(n_956),
.B2(n_979),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1006),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1010),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_1001),
.B(n_945),
.Y(n_1014)
);

NOR2x1p5_ASAP7_75t_L g1015 ( 
.A(n_1000),
.B(n_813),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1003),
.B(n_965),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_1004),
.A2(n_956),
.B1(n_979),
.B2(n_984),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1009),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1005),
.B(n_984),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1013),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1015),
.B(n_1008),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1016),
.A2(n_1008),
.B1(n_1002),
.B2(n_918),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1014),
.Y(n_1023)
);

OA21x2_ASAP7_75t_L g1024 ( 
.A1(n_1012),
.A2(n_755),
.B(n_821),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_1017),
.A2(n_835),
.B(n_822),
.Y(n_1025)
);

OA21x2_ASAP7_75t_L g1026 ( 
.A1(n_1019),
.A2(n_832),
.B(n_852),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1018),
.Y(n_1027)
);

AOI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_1019),
.A2(n_1011),
.B1(n_965),
.B2(n_749),
.C(n_942),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_1027),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1020),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1021),
.B(n_948),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1023),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1022),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_961),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1024),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1028),
.B(n_948),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1031),
.B(n_1026),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1032),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1029),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1029),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_1026),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1030),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1035),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_1036),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_1024),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1043),
.Y(n_1046)
);

NOR3xp33_ASAP7_75t_L g1047 ( 
.A(n_1039),
.B(n_1034),
.C(n_833),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1040),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

NAND4xp25_ASAP7_75t_L g1050 ( 
.A(n_1044),
.B(n_813),
.C(n_736),
.D(n_808),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1038),
.A2(n_759),
.B(n_837),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1042),
.B(n_736),
.C(n_752),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_SL g1053 ( 
.A(n_1041),
.B(n_862),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1045),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_R g1055 ( 
.A(n_1049),
.B(n_1045),
.Y(n_1055)
);

OAI211xp5_ASAP7_75t_L g1056 ( 
.A1(n_1048),
.A2(n_1037),
.B(n_922),
.C(n_752),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1047),
.A2(n_810),
.B1(n_757),
.B2(n_951),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_1054),
.A2(n_739),
.B1(n_740),
.B2(n_942),
.C(n_848),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1053),
.A2(n_810),
.B1(n_764),
.B2(n_912),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1046),
.Y(n_1060)
);

OAI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_1050),
.A2(n_955),
.B(n_936),
.Y(n_1061)
);

OAI21xp33_ASAP7_75t_SL g1062 ( 
.A1(n_1057),
.A2(n_1051),
.B(n_1052),
.Y(n_1062)
);

AOI221xp5_ASAP7_75t_L g1063 ( 
.A1(n_1056),
.A2(n_740),
.B1(n_848),
.B2(n_944),
.C(n_946),
.Y(n_1063)
);

AOI211xp5_ASAP7_75t_L g1064 ( 
.A1(n_1060),
.A2(n_851),
.B(n_750),
.C(n_955),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_1061),
.B(n_955),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1059),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1058),
.A2(n_944),
.B1(n_946),
.B2(n_949),
.C(n_793),
.Y(n_1067)
);

OAI211xp5_ASAP7_75t_SL g1068 ( 
.A1(n_1055),
.A2(n_810),
.B(n_946),
.C(n_949),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1060),
.Y(n_1069)
);

OAI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1060),
.A2(n_748),
.B(n_750),
.C(n_850),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_SL g1071 ( 
.A(n_1069),
.B(n_748),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1065),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1062),
.A2(n_951),
.B(n_748),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1068),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1066),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1070),
.A2(n_912),
.B1(n_953),
.B2(n_951),
.Y(n_1076)
);

AOI321xp33_ASAP7_75t_L g1077 ( 
.A1(n_1067),
.A2(n_894),
.A3(n_899),
.B1(n_897),
.B2(n_895),
.C(n_882),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_1063),
.A2(n_750),
.B1(n_953),
.B2(n_826),
.C(n_805),
.Y(n_1078)
);

OAI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_1064),
.A2(n_756),
.B1(n_746),
.B2(n_879),
.C(n_875),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_1069),
.Y(n_1080)
);

INVx3_ASAP7_75t_SL g1081 ( 
.A(n_1075),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1072),
.B(n_881),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1080),
.B(n_881),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1074),
.B(n_1071),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1073),
.B(n_934),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_1079),
.B(n_934),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_1076),
.B(n_972),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_1078),
.Y(n_1088)
);

NAND3x2_ASAP7_75t_L g1089 ( 
.A(n_1077),
.B(n_140),
.C(n_141),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_L g1090 ( 
.A(n_1075),
.B(n_850),
.C(n_826),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1075),
.B(n_972),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1080),
.B(n_142),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1075),
.B(n_972),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1081),
.A2(n_850),
.B1(n_826),
.B2(n_807),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1082),
.B(n_924),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_1083),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1090),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1092),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1087),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1084),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1088),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1091),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_1101),
.A2(n_1093),
.B1(n_1086),
.B2(n_1085),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_1096),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1101),
.B(n_1089),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1100),
.A2(n_756),
.B(n_887),
.Y(n_1106)
);

XNOR2xp5_ASAP7_75t_L g1107 ( 
.A(n_1098),
.B(n_143),
.Y(n_1107)
);

AO21x2_ASAP7_75t_L g1108 ( 
.A1(n_1099),
.A2(n_145),
.B(n_147),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1094),
.A2(n_807),
.B1(n_826),
.B2(n_850),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1102),
.A2(n_881),
.B1(n_807),
.B2(n_805),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_SL g1111 ( 
.A1(n_1104),
.A2(n_1097),
.B1(n_1095),
.B2(n_807),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1103),
.A2(n_881),
.B1(n_883),
.B2(n_151),
.C(n_152),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1105),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1111),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1114),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_1113),
.B(n_1112),
.Y(n_1116)
);

OAI211xp5_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_1110),
.B(n_1106),
.C(n_1108),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1116),
.A2(n_1107),
.B1(n_1109),
.B2(n_881),
.Y(n_1118)
);

OAI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_1116),
.A2(n_746),
.B1(n_150),
.B2(n_153),
.C(n_158),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1117),
.A2(n_149),
.B(n_160),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1118),
.A2(n_163),
.B(n_164),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1119),
.A2(n_165),
.B(n_166),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_SL g1123 ( 
.A1(n_1120),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1121),
.A2(n_879),
.B1(n_875),
.B2(n_894),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1123),
.A2(n_1124),
.B(n_1125),
.Y(n_1126)
);

AO221x2_ASAP7_75t_L g1127 ( 
.A1(n_1123),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.C(n_182),
.Y(n_1127)
);

NAND3x2_ASAP7_75t_L g1128 ( 
.A(n_1123),
.B(n_183),
.C(n_184),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_1127),
.B(n_1128),
.Y(n_1129)
);

AOI211xp5_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_186),
.B(n_187),
.C(n_189),
.Y(n_1130)
);


endmodule