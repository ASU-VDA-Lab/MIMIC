module real_jpeg_33513_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_0),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_0),
.Y(n_437)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_0),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_537),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_1),
.B(n_538),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_2),
.Y(n_201)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

NAND2x1p5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_4),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_4),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_4),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_4),
.B(n_153),
.Y(n_152)
);

NAND2x1_ASAP7_75t_L g155 ( 
.A(n_4),
.B(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_5),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_5),
.Y(n_213)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_6),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_6),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_6),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_6),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_6),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_6),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_6),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_7),
.B(n_28),
.Y(n_27)
);

NAND2x1_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_R g100 ( 
.A(n_7),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_7),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_7),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_7),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_7),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_7),
.B(n_153),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_8),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_8),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_8),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_8),
.B(n_131),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_8),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_8),
.B(n_303),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_8),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g196 ( 
.A(n_10),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_10),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_10),
.B(n_34),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_10),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_10),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_10),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_10),
.B(n_288),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_11),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_12),
.B(n_104),
.Y(n_251)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_12),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_12),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_12),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_12),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_12),
.B(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_12),
.B(n_478),
.Y(n_477)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_13),
.Y(n_171)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_13),
.Y(n_454)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_14),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_15),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_16),
.B(n_76),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_16),
.B(n_366),
.Y(n_365)
);

BUFx24_ASAP7_75t_L g394 ( 
.A(n_16),
.Y(n_394)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_16),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_17),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_17),
.B(n_131),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_17),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_212),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_17),
.B(n_153),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_183),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_180),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_112),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_23),
.B(n_112),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_85),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_52),
.C(n_70),
.Y(n_24)
);

XNOR2x1_ASAP7_75t_L g113 ( 
.A(n_25),
.B(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_26),
.B(n_42),
.C(n_51),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.C(n_37),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_27),
.A2(n_32),
.B1(n_33),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_27),
.Y(n_141)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_31),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_32),
.A2(n_33),
.B1(n_196),
.B2(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_33),
.B(n_195),
.C(n_196),
.Y(n_194)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_35),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_36),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_37),
.B(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_40),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_40),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_51),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_46),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_46),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_48),
.B(n_194),
.C(n_199),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_48),
.A2(n_49),
.B1(n_199),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_49),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_51),
.B(n_143),
.C(n_155),
.Y(n_142)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_71),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.C(n_65),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_61),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_60),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_61),
.B(n_167),
.C(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_64),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_66),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_65),
.A2(n_66),
.B1(n_319),
.B2(n_390),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_121),
.C(n_125),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_66),
.B(n_121),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_66),
.B(n_319),
.C(n_322),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_69),
.Y(n_253)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_69),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_80),
.C(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_80),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_80),
.B(n_130),
.C(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_80),
.B(n_238),
.Y(n_331)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_84),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B1(n_110),
.B2(n_111),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_130),
.C(n_133),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_94),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_96),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_96),
.A2(n_98),
.B1(n_252),
.B2(n_306),
.Y(n_305)
);

INVx8_ASAP7_75t_L g396 ( 
.A(n_97),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_98),
.B(n_247),
.C(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.C(n_137),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_113),
.B(n_115),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_129),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_116),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_120),
.B(n_129),
.Y(n_224)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_123),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_124),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_146),
.B(n_154),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_126),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_125),
.A2(n_126),
.B1(n_147),
.B2(n_148),
.Y(n_205)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_126),
.B(n_250),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_128),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_133),
.B1(n_134),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_130),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_130),
.A2(n_178),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_132),
.Y(n_325)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_132),
.Y(n_479)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_136),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_142),
.C(n_157),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_144),
.A2(n_145),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_152),
.Y(n_154)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_207),
.C(n_210),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_151),
.B(n_235),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g489 ( 
.A1(n_151),
.A2(n_152),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_151),
.B(n_490),
.Y(n_503)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_152),
.B(n_211),
.Y(n_360)
);

INVx4_ASAP7_75t_SL g316 ( 
.A(n_153),
.Y(n_316)
);

INVx8_ASAP7_75t_L g442 ( 
.A(n_153),
.Y(n_442)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_158),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_163),
.B1(n_174),
.B2(n_179),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_159),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_164),
.B(n_176),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.C(n_172),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_172),
.Y(n_216)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_168),
.A2(n_215),
.B1(n_295),
.B2(n_296),
.Y(n_356)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_266),
.B(n_532),
.Y(n_183)
);

NAND2x1_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_228),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_225),
.Y(n_185)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_186),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.C(n_223),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_191),
.B(n_223),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_202),
.C(n_217),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_192),
.A2(n_193),
.B1(n_218),
.B2(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_194),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_195),
.B(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_196),
.Y(n_244)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_203),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_214),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_204),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_206),
.B(n_214),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_211),
.B(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_211),
.A2(n_236),
.B1(n_314),
.B2(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_225),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_264),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_229),
.B(n_264),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_258),
.C(n_261),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_230),
.B(n_416),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_245),
.B(n_257),
.Y(n_230)
);

HB1xp67_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_232),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.C(n_242),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_237),
.Y(n_338)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_254),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_SL g344 ( 
.A(n_246),
.B(n_254),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.C(n_251),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_251),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_259),
.B(n_262),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_418),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_348),
.B(n_409),
.C(n_410),
.D(n_417),
.Y(n_267)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_268),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_339),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_269),
.B(n_339),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_307),
.C(n_333),
.Y(n_269)
);

INVxp33_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_271),
.A2(n_334),
.B1(n_335),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_271),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_292),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_272),
.B(n_293),
.C(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.C(n_280),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_273),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_275),
.A2(n_276),
.B1(n_280),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g357 ( 
.A1(n_276),
.A2(n_277),
.B(n_279),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_280),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.C(n_291),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_281),
.A2(n_286),
.B1(n_287),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_290),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_304),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.C(n_301),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_297),
.A2(n_298),
.B1(n_301),
.B2(n_302),
.Y(n_327)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_303),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_304),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_307),
.B(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_326),
.C(n_329),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_308),
.B(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.C(n_317),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_312),
.A2(n_313),
.B1(n_317),
.B2(n_318),
.Y(n_385)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_314),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_319),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g388 ( 
.A(n_322),
.B(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_330),
.Y(n_352)
);

XOR2x1_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_345),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

AOI21x1_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_377),
.B(n_408),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_374),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_350),
.B(n_374),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.C(n_369),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_370),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.C(n_358),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_357),
.Y(n_383)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.C(n_365),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_360),
.B(n_519),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_361),
.B(n_365),
.Y(n_519)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_380),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_378),
.B(n_380),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.C(n_386),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_382),
.A2(n_386),
.B1(n_387),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_382),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_384),
.B(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.C(n_405),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_388),
.B(n_514),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_391),
.A2(n_405),
.B1(n_406),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_391),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_397),
.C(n_401),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_392),
.A2(n_393),
.B1(n_401),
.B2(n_402),
.Y(n_499)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_394),
.B(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_394),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_394),
.B(n_481),
.Y(n_480)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_397),
.B(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_400),
.Y(n_449)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_408),
.Y(n_528)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_415),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_415),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.C(n_414),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_528),
.C(n_529),
.Y(n_418)
);

NOR2x1p5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

AOI21x1_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_522),
.B(n_527),
.Y(n_421)
);

OAI21x1_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_511),
.B(n_521),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_493),
.B(n_510),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_472),
.B(n_492),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_426),
.A2(n_455),
.B(n_471),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_438),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_427),
.B(n_438),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_434),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_428),
.A2(n_429),
.B1(n_434),
.B2(n_435),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_428),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

BUFx4f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_447),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_439),
.B(n_448),
.C(n_450),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_443),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_440),
.B(n_443),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_507),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_444),
.B(n_483),
.Y(n_482)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_450),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_453),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_464),
.B(n_470),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_463),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_463),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_474),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_485),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_486),
.C(n_489),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_482),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_480),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_477),
.B(n_480),
.C(n_482),
.Y(n_501)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_490),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_495),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_496),
.A2(n_502),
.B1(n_508),
.B2(n_509),
.Y(n_495)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_496),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_498),
.B1(n_500),
.B2(n_501),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_501),
.C(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_502),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_504),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_505),
.C(n_506),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_520),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_520),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_517),
.C(n_518),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_526),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_533),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_535),
.C(n_536),
.Y(n_533)
);


endmodule