module fake_jpeg_2635_n_535 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_535);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_535;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_56),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_57),
.Y(n_174)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_58),
.Y(n_111)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_64),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_7),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_16),
.C(n_7),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_68),
.B(n_23),
.C(n_39),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_23),
.B(n_6),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_77),
.Y(n_171)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_78),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_94),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_98),
.B(n_110),
.Y(n_161)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_21),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_104),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_32),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_28),
.B(n_6),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_44),
.Y(n_142)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_47),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_52),
.Y(n_122)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_52),
.B1(n_51),
.B2(n_30),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_113),
.A2(n_129),
.B1(n_169),
.B2(n_19),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx4_ASAP7_75t_SL g210 ( 
.A(n_122),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_37),
.B1(n_26),
.B2(n_49),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_36),
.C(n_33),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_88),
.B(n_38),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_131),
.B(n_140),
.Y(n_188)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_133),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_30),
.Y(n_140)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_142),
.B(n_145),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_39),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_155),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_78),
.B(n_51),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_110),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_44),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_95),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_36),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_42),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_101),
.A2(n_51),
.B1(n_26),
.B2(n_19),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_SL g177 ( 
.A(n_166),
.Y(n_177)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_178),
.A2(n_200),
.B1(n_224),
.B2(n_228),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_179),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_33),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_217),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_117),
.A2(n_103),
.B1(n_79),
.B2(n_65),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_182),
.A2(n_187),
.B1(n_205),
.B2(n_229),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_183),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_116),
.B1(n_87),
.B2(n_109),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_214),
.B1(n_227),
.B2(n_171),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_119),
.A2(n_89),
.B1(n_86),
.B2(n_85),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_197),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_191),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_37),
.B1(n_42),
.B2(n_38),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_206),
.Y(n_230)
);

BUFx16f_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_196),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_161),
.A2(n_57),
.B(n_72),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_198),
.B(n_221),
.Y(n_263)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_111),
.A2(n_49),
.B1(n_53),
.B2(n_107),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

BUFx4f_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_125),
.A2(n_82),
.B1(n_63),
.B2(n_71),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_134),
.B(n_92),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_152),
.A2(n_96),
.B(n_22),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_207),
.B(n_174),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_114),
.A2(n_35),
.B(n_41),
.Y(n_209)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_31),
.A3(n_143),
.B1(n_128),
.B2(n_41),
.Y(n_254)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_211),
.Y(n_268)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_129),
.A2(n_135),
.B1(n_170),
.B2(n_168),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_115),
.B(n_106),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_218),
.Y(n_256)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_124),
.B(n_0),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_138),
.B(n_99),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_126),
.B(n_0),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_223),
.Y(n_248)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_1),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_156),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_171),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_172),
.A2(n_93),
.B1(n_90),
.B2(n_83),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_111),
.A2(n_49),
.B1(n_76),
.B2(n_75),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_232),
.A2(n_242),
.B1(n_250),
.B2(n_264),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_153),
.B1(n_144),
.B2(n_157),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_233),
.A2(n_239),
.B1(n_249),
.B2(n_133),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_173),
.C(n_151),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_265),
.C(n_196),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_160),
.B1(n_153),
.B2(n_157),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_210),
.A2(n_175),
.B1(n_172),
.B2(n_160),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_127),
.B1(n_146),
.B2(n_149),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_175),
.B1(n_127),
.B2(n_154),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g252 ( 
.A1(n_227),
.A2(n_146),
.B1(n_128),
.B2(n_143),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_221),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_197),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_259),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_217),
.A2(n_158),
.B1(n_154),
.B2(n_149),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_211),
.C(n_186),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_270),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_278),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_231),
.B(n_188),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_272),
.B(n_279),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_222),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_275),
.B(n_280),
.Y(n_309)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_276),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_232),
.A2(n_219),
.B1(n_202),
.B2(n_225),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_282),
.B1(n_242),
.B2(n_237),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_196),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_231),
.B(n_201),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_216),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

BUFx24_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_262),
.A2(n_213),
.B1(n_199),
.B2(n_193),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_283),
.A2(n_290),
.B1(n_299),
.B2(n_141),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_220),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_224),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_296),
.C(n_298),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_230),
.B(n_192),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_252),
.B1(n_240),
.B2(n_267),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_291),
.Y(n_317)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_212),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_302),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_248),
.B(n_156),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_297),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_183),
.C(n_181),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_228),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_208),
.C(n_190),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_190),
.C(n_226),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_249),
.Y(n_311)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_258),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_239),
.B1(n_257),
.B2(n_233),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_306),
.A2(n_323),
.B1(n_330),
.B2(n_237),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_297),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_307),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_277),
.A2(n_264),
.B1(n_240),
.B2(n_250),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_308),
.A2(n_328),
.B(n_300),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_253),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_261),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_312),
.B(n_334),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_274),
.A2(n_252),
.B1(n_269),
.B2(n_244),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_327),
.Y(n_339)
);

NOR2x1p5_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_274),
.Y(n_319)
);

NAND2x1p5_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_226),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

OAI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_322),
.A2(n_299),
.B(n_294),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_252),
.B1(n_269),
.B2(n_244),
.Y(n_323)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_280),
.Y(n_326)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_266),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_284),
.A2(n_247),
.B(n_245),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_283),
.A2(n_252),
.B1(n_243),
.B2(n_246),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_329),
.A2(n_291),
.B1(n_301),
.B2(n_276),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_266),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_342),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_279),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_336),
.Y(n_368)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_273),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_272),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_296),
.B(n_278),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_341),
.A2(n_344),
.B(n_351),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_328),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_319),
.A2(n_304),
.B(n_305),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_325),
.B(n_286),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_350),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_298),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_353),
.C(n_360),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_303),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_349),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_258),
.Y(n_349)
);

AO22x1_ASAP7_75t_SL g352 ( 
.A1(n_313),
.A2(n_282),
.B1(n_281),
.B2(n_237),
.Y(n_352)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_362),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_308),
.A2(n_307),
.B1(n_329),
.B2(n_305),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_361),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_314),
.B(n_253),
.Y(n_360)
);

AO22x1_ASAP7_75t_L g361 ( 
.A1(n_323),
.A2(n_238),
.B1(n_281),
.B2(n_192),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_306),
.A2(n_243),
.B1(n_246),
.B2(n_281),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_292),
.Y(n_363)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_363),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_364),
.A2(n_334),
.B(n_322),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_364),
.A2(n_311),
.B(n_314),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_384),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_363),
.Y(n_375)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_378),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_355),
.B(n_321),
.Y(n_380)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_382),
.Y(n_412)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_383),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_346),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_388),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_318),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_386),
.B(n_185),
.Y(n_418)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_337),
.Y(n_387)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_332),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_341),
.A2(n_332),
.B1(n_317),
.B2(n_310),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_390),
.A2(n_356),
.B1(n_354),
.B2(n_342),
.Y(n_396)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_392),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_336),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_324),
.C(n_310),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_352),
.C(n_235),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_331),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_389),
.Y(n_427)
);

XNOR2x1_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_343),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_SL g425 ( 
.A(n_397),
.B(n_384),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_382),
.A2(n_359),
.B1(n_358),
.B2(n_364),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_399),
.A2(n_409),
.B1(n_421),
.B2(n_423),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_369),
.B(n_359),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_404),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_380),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_351),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_414),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_388),
.B(n_350),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_407),
.B(n_376),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_383),
.A2(n_352),
.B1(n_362),
.B2(n_347),
.Y(n_409)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_410),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_366),
.B(n_235),
.C(n_176),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_417),
.C(n_419),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_289),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_379),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_204),
.C(n_179),
.Y(n_417)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_212),
.C(n_316),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_368),
.A2(n_361),
.B1(n_302),
.B2(n_316),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_316),
.C(n_361),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_381),
.C(n_374),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_389),
.A2(n_316),
.B1(n_159),
.B2(n_260),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_121),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_387),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_429),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_411),
.B(n_377),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_426),
.B(n_432),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_409),
.B1(n_414),
.B2(n_398),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_390),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_430),
.B(n_397),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_374),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_159),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_400),
.A2(n_377),
.B(n_401),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_444),
.Y(n_450)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_408),
.A2(n_392),
.B1(n_395),
.B2(n_376),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_437),
.A2(n_422),
.B1(n_420),
.B2(n_395),
.Y(n_454)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_440),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_391),
.C(n_370),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_447),
.C(n_448),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_378),
.Y(n_443)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_370),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_445),
.B(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_446),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_375),
.C(n_367),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_367),
.C(n_365),
.Y(n_448)
);

OAI22x1_ASAP7_75t_SL g449 ( 
.A1(n_433),
.A2(n_396),
.B1(n_412),
.B2(n_413),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_449),
.A2(n_454),
.B1(n_461),
.B2(n_464),
.Y(n_478)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_460),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_466),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_439),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_SL g461 ( 
.A1(n_427),
.A2(n_400),
.B(n_423),
.C(n_424),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_436),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_462),
.B(n_15),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_438),
.A2(n_400),
.B1(n_365),
.B2(n_379),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_163),
.C(n_158),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_467),
.B(n_163),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_465),
.B(n_428),
.C(n_448),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_469),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_465),
.B(n_428),
.C(n_441),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_442),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_461),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_447),
.C(n_429),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_473),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_434),
.C(n_431),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_430),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_474),
.B(n_476),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_475),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_444),
.C(n_425),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_479),
.B(n_483),
.Y(n_486)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_482),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_158),
.C(n_154),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_458),
.A2(n_120),
.B(n_238),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_484),
.B(n_456),
.C(n_467),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_466),
.C(n_455),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_491),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_493),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_472),
.C(n_473),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_449),
.C(n_459),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_492),
.B(n_9),
.Y(n_508)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_478),
.B(n_461),
.CI(n_120),
.CON(n_493),
.SN(n_493)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_461),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_496),
.A2(n_10),
.B(n_12),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_77),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_499),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_49),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_31),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_10),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_496),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_501)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_501),
.Y(n_519)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_506),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_1),
.C(n_2),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_508),
.B(n_510),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_491),
.A2(n_490),
.B(n_497),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_509),
.A2(n_511),
.B(n_486),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_488),
.A2(n_10),
.B1(n_2),
.B2(n_5),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_485),
.B(n_6),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_506),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_513),
.B(n_500),
.Y(n_521)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_514),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_495),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_517),
.C(n_503),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_498),
.C(n_499),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_516),
.A2(n_10),
.B(n_12),
.Y(n_526)
);

AO21x1_ASAP7_75t_L g525 ( 
.A1(n_521),
.A2(n_505),
.B(n_493),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_522),
.A2(n_515),
.B(n_520),
.Y(n_527)
);

AOI31xp33_ASAP7_75t_L g524 ( 
.A1(n_519),
.A2(n_513),
.A3(n_507),
.B(n_503),
.Y(n_524)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_524),
.A2(n_525),
.B(n_526),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_527),
.B(n_529),
.Y(n_531)
);

AOI322xp5_ASAP7_75t_L g529 ( 
.A1(n_523),
.A2(n_518),
.A3(n_521),
.B1(n_13),
.B2(n_15),
.C1(n_12),
.C2(n_1),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_524),
.C(n_15),
.Y(n_530)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_530),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_531),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_15),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_1),
.Y(n_535)
);


endmodule