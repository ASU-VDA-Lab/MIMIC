module real_aes_8166_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g513 ( .A1(n_0), .A2(n_156), .B(n_514), .C(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_1), .B(n_175), .Y(n_517) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_3), .A2(n_142), .B(n_147), .C(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_4), .A2(n_137), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_5), .B(n_212), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_6), .A2(n_137), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_7), .B(n_175), .Y(n_241) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_8), .A2(n_160), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g142 ( .A(n_9), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_10), .A2(n_142), .B(n_147), .C(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g154 ( .A(n_11), .Y(n_154) );
INVx1_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_12), .B(n_41), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_13), .B(n_152), .Y(n_189) );
INVx1_ASAP7_75t_L g135 ( .A(n_14), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_15), .B(n_212), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g168 ( .A1(n_16), .A2(n_155), .B(n_169), .C(n_173), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_17), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_18), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_19), .B(n_281), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_20), .A2(n_199), .B(n_200), .C(n_202), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_21), .A2(n_147), .B(n_216), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_22), .B(n_152), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_23), .B(n_152), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_24), .Y(n_223) );
INVx1_ASAP7_75t_L g211 ( .A(n_25), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_26), .A2(n_147), .B(n_216), .C(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_27), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_28), .Y(n_182) );
INVx1_ASAP7_75t_L g277 ( .A(n_29), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_30), .A2(n_137), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g140 ( .A(n_31), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_32), .A2(n_228), .B(n_449), .C(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_33), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_34), .A2(n_199), .B(n_237), .C(n_239), .Y(n_236) );
INVxp67_ASAP7_75t_L g278 ( .A(n_35), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_36), .B(n_473), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_37), .A2(n_147), .B(n_210), .C(n_216), .Y(n_209) );
CKINVDCx14_ASAP7_75t_R g235 ( .A(n_38), .Y(n_235) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_39), .A2(n_46), .B1(n_744), .B2(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_39), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_40), .A2(n_45), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_40), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_41), .B(n_108), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_42), .A2(n_151), .B(n_153), .C(n_156), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_43), .B(n_272), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_44), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_45), .Y(n_728) );
INVx1_ASAP7_75t_L g745 ( .A(n_46), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_47), .B(n_212), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_48), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_49), .B(n_137), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_50), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_51), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_52), .A2(n_228), .B(n_449), .C(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g516 ( .A(n_53), .Y(n_516) );
INVx1_ASAP7_75t_L g451 ( .A(n_54), .Y(n_451) );
INVx1_ASAP7_75t_L g197 ( .A(n_55), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_56), .B(n_137), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_57), .Y(n_497) );
CKINVDCx14_ASAP7_75t_R g145 ( .A(n_58), .Y(n_145) );
INVx1_ASAP7_75t_L g143 ( .A(n_59), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_60), .B(n_137), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_61), .B(n_175), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_62), .A2(n_215), .B(n_462), .C(n_463), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_63), .A2(n_102), .B1(n_116), .B2(n_754), .Y(n_101) );
INVx1_ASAP7_75t_L g134 ( .A(n_64), .Y(n_134) );
INVx1_ASAP7_75t_SL g238 ( .A(n_65), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_66), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_67), .B(n_212), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_68), .B(n_175), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_69), .B(n_155), .Y(n_526) );
INVx1_ASAP7_75t_L g226 ( .A(n_70), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g512 ( .A(n_71), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_72), .B(n_188), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_73), .A2(n_147), .B(n_228), .C(n_502), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_74), .Y(n_460) );
INVx1_ASAP7_75t_L g115 ( .A(n_75), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_76), .A2(n_137), .B(n_144), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_77), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_78), .A2(n_137), .B(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_79), .A2(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g167 ( .A(n_80), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_81), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_82), .B(n_187), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_83), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_84), .A2(n_137), .B(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g170 ( .A(n_85), .Y(n_170) );
INVx2_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g186 ( .A(n_87), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_88), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_89), .B(n_152), .Y(n_527) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
OR2x2_ASAP7_75t_L g440 ( .A(n_90), .B(n_123), .Y(n_440) );
OR2x2_ASAP7_75t_L g747 ( .A(n_90), .B(n_735), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_91), .A2(n_147), .B(n_225), .C(n_228), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_92), .B(n_137), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_93), .Y(n_484) );
INVxp67_ASAP7_75t_L g464 ( .A(n_94), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_95), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_96), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g201 ( .A(n_97), .Y(n_201) );
INVx1_ASAP7_75t_L g503 ( .A(n_98), .Y(n_503) );
INVx1_ASAP7_75t_L g523 ( .A(n_99), .Y(n_523) );
AND2x2_ASAP7_75t_L g454 ( .A(n_100), .B(n_131), .Y(n_454) );
BUFx4f_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g754 ( .A(n_105), .Y(n_754) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .C(n_113), .Y(n_110) );
AND2x2_ASAP7_75t_L g123 ( .A(n_111), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g122 ( .A(n_112), .B(n_123), .Y(n_122) );
NOR2x2_ASAP7_75t_L g734 ( .A(n_112), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO221x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_737), .B1(n_740), .B2(n_748), .C(n_750), .Y(n_116) );
OAI222xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_726), .B1(n_727), .B2(n_730), .C1(n_733), .C2(n_736), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_125), .B1(n_437), .B2(n_441), .Y(n_118) );
AOI22x1_ASAP7_75t_SL g730 ( .A1(n_119), .A2(n_437), .B1(n_731), .B2(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g735 ( .A(n_123), .Y(n_735) );
INVx2_ASAP7_75t_L g731 ( .A(n_125), .Y(n_731) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_367), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_282), .C(n_314), .D(n_331), .E(n_354), .Y(n_126) );
AOI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_205), .B1(n_242), .B2(n_246), .C(n_250), .Y(n_127) );
INVx1_ASAP7_75t_L g394 ( .A(n_128), .Y(n_394) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_177), .Y(n_128) );
AND3x2_ASAP7_75t_L g369 ( .A(n_129), .B(n_179), .C(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_162), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_130), .B(n_248), .Y(n_247) );
BUFx3_ASAP7_75t_L g257 ( .A(n_130), .Y(n_257) );
AND2x2_ASAP7_75t_L g261 ( .A(n_130), .B(n_193), .Y(n_261) );
INVx2_ASAP7_75t_L g291 ( .A(n_130), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_130), .B(n_194), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_130), .B(n_178), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_130), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g381 ( .A(n_130), .B(n_194), .Y(n_381) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_136), .B(n_159), .Y(n_130) );
INVx1_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_131), .A2(n_183), .B(n_208), .C(n_209), .Y(n_207) );
INVx2_ASAP7_75t_L g231 ( .A(n_131), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_131), .A2(n_447), .B(n_448), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_131), .A2(n_481), .B(n_482), .Y(n_480) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_L g161 ( .A(n_132), .B(n_133), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx2_ASAP7_75t_L g272 ( .A(n_137), .Y(n_272) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_138), .B(n_142), .Y(n_183) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g215 ( .A(n_139), .Y(n_215) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx1_ASAP7_75t_L g203 ( .A(n_140), .Y(n_203) );
INVx1_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_141), .Y(n_155) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_141), .Y(n_172) );
INVx1_ASAP7_75t_L g473 ( .A(n_141), .Y(n_473) );
INVx4_ASAP7_75t_SL g158 ( .A(n_142), .Y(n_158) );
BUFx3_ASAP7_75t_L g216 ( .A(n_142), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_146), .B(n_150), .C(n_158), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_SL g166 ( .A1(n_146), .A2(n_158), .B(n_167), .C(n_168), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g196 ( .A1(n_146), .A2(n_158), .B(n_197), .C(n_198), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_146), .A2(n_158), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g273 ( .A1(n_146), .A2(n_158), .B(n_274), .C(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g449 ( .A(n_146), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_146), .A2(n_158), .B(n_460), .C(n_461), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_146), .A2(n_158), .B(n_512), .C(n_513), .Y(n_511) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_148), .Y(n_240) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx5_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
INVx2_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g173 ( .A(n_157), .Y(n_173) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_157), .Y(n_453) );
INVx1_ASAP7_75t_L g228 ( .A(n_158), .Y(n_228) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_160), .Y(n_164) );
INVx4_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_160), .A2(n_469), .B(n_470), .Y(n_468) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g269 ( .A(n_161), .Y(n_269) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_162), .Y(n_260) );
AND2x2_ASAP7_75t_L g322 ( .A(n_162), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_162), .B(n_178), .Y(n_341) );
INVx1_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g249 ( .A(n_163), .B(n_178), .Y(n_249) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_163), .Y(n_256) );
AND2x2_ASAP7_75t_L g308 ( .A(n_163), .B(n_194), .Y(n_308) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_163), .B(n_177), .C(n_291), .Y(n_333) );
AND2x2_ASAP7_75t_L g398 ( .A(n_163), .B(n_179), .Y(n_398) );
AND2x2_ASAP7_75t_L g432 ( .A(n_163), .B(n_178), .Y(n_432) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_174), .Y(n_163) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_164), .A2(n_195), .B(n_204), .Y(n_194) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_164), .A2(n_233), .B(n_241), .Y(n_232) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_164), .A2(n_458), .B(n_465), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_171), .B(n_201), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_171), .A2(n_212), .B1(n_277), .B2(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g462 ( .A(n_171), .Y(n_462) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g188 ( .A(n_172), .Y(n_188) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_175), .A2(n_510), .B(n_517), .Y(n_509) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_176), .B(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_176), .B(n_218), .Y(n_217) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_176), .A2(n_222), .B(n_229), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_176), .B(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g499 ( .A1(n_176), .A2(n_500), .B(n_507), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_176), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_176), .A2(n_522), .B(n_528), .Y(n_521) );
INVxp67_ASAP7_75t_L g258 ( .A(n_177), .Y(n_258) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_178), .B(n_291), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_178), .B(n_322), .Y(n_330) );
AND2x2_ASAP7_75t_L g380 ( .A(n_178), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g408 ( .A(n_178), .Y(n_408) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g315 ( .A(n_179), .B(n_308), .Y(n_315) );
BUFx3_ASAP7_75t_L g347 ( .A(n_179), .Y(n_347) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_191), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_180), .B(n_497), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_184), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_183), .A2(n_223), .B(n_224), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_183), .A2(n_523), .B(n_524), .Y(n_522) );
O2A1O1Ixp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_189), .C(n_190), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_187), .A2(n_190), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_187), .A2(n_451), .B(n_452), .C(n_453), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_187), .A2(n_453), .B(n_484), .C(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g323 ( .A(n_193), .Y(n_323) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_194), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_199), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_199), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g475 ( .A(n_202), .Y(n_475) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_205), .A2(n_383), .B1(n_385), .B2(n_386), .Y(n_382) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_219), .Y(n_205) );
AND2x2_ASAP7_75t_L g242 ( .A(n_206), .B(n_243), .Y(n_242) );
INVx3_ASAP7_75t_SL g253 ( .A(n_206), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_206), .B(n_286), .Y(n_318) );
OR2x2_ASAP7_75t_L g337 ( .A(n_206), .B(n_220), .Y(n_337) );
AND2x2_ASAP7_75t_L g342 ( .A(n_206), .B(n_294), .Y(n_342) );
AND2x2_ASAP7_75t_L g345 ( .A(n_206), .B(n_287), .Y(n_345) );
AND2x2_ASAP7_75t_L g357 ( .A(n_206), .B(n_232), .Y(n_357) );
AND2x2_ASAP7_75t_L g373 ( .A(n_206), .B(n_221), .Y(n_373) );
AND2x4_ASAP7_75t_L g376 ( .A(n_206), .B(n_244), .Y(n_376) );
OR2x2_ASAP7_75t_L g393 ( .A(n_206), .B(n_329), .Y(n_393) );
OR2x2_ASAP7_75t_L g424 ( .A(n_206), .B(n_266), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_206), .B(n_352), .Y(n_426) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .C(n_214), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_212), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g514 ( .A(n_212), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_214), .A2(n_494), .B(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_215), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g300 ( .A(n_219), .B(n_264), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_219), .B(n_287), .Y(n_419) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_232), .Y(n_219) );
AND2x2_ASAP7_75t_L g252 ( .A(n_220), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g286 ( .A(n_220), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g294 ( .A(n_220), .B(n_266), .Y(n_294) );
AND2x2_ASAP7_75t_L g312 ( .A(n_220), .B(n_244), .Y(n_312) );
OR2x2_ASAP7_75t_L g329 ( .A(n_220), .B(n_287), .Y(n_329) );
INVx2_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
BUFx2_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
AND2x2_ASAP7_75t_L g352 ( .A(n_221), .B(n_232), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx1_ASAP7_75t_L g281 ( .A(n_231), .Y(n_281) );
INVx2_ASAP7_75t_L g244 ( .A(n_232), .Y(n_244) );
INVx1_ASAP7_75t_L g364 ( .A(n_232), .Y(n_364) );
AND2x2_ASAP7_75t_L g414 ( .A(n_232), .B(n_253), .Y(n_414) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_240), .Y(n_505) );
AND2x2_ASAP7_75t_L g263 ( .A(n_243), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g298 ( .A(n_243), .B(n_253), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_243), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g285 ( .A(n_244), .B(n_253), .Y(n_285) );
OR2x2_ASAP7_75t_L g401 ( .A(n_245), .B(n_375), .Y(n_401) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_248), .B(n_381), .Y(n_387) );
INVx2_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OAI32xp33_ASAP7_75t_L g343 ( .A1(n_249), .A2(n_344), .A3(n_346), .B1(n_348), .B2(n_349), .Y(n_343) );
OR2x2_ASAP7_75t_L g360 ( .A(n_249), .B(n_302), .Y(n_360) );
OAI21xp33_ASAP7_75t_SL g385 ( .A1(n_249), .A2(n_259), .B(n_290), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_254), .B1(n_259), .B2(n_262), .Y(n_250) );
INVxp33_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_252), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_253), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g311 ( .A(n_253), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g411 ( .A(n_253), .B(n_352), .Y(n_411) );
OR2x2_ASAP7_75t_L g435 ( .A(n_253), .B(n_329), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_254), .A2(n_317), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g295 ( .A(n_256), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_256), .B(n_261), .Y(n_313) );
AND2x2_ASAP7_75t_L g335 ( .A(n_257), .B(n_308), .Y(n_335) );
INVx1_ASAP7_75t_L g348 ( .A(n_257), .Y(n_348) );
OR2x2_ASAP7_75t_L g353 ( .A(n_257), .B(n_287), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_260), .B(n_302), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g283 ( .A1(n_261), .A2(n_284), .B1(n_289), .B2(n_293), .Y(n_283) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_264), .A2(n_326), .B1(n_333), .B2(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g410 ( .A(n_264), .B(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_266), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g429 ( .A(n_266), .B(n_312), .Y(n_429) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B(n_279), .Y(n_266) );
INVx1_ASAP7_75t_L g288 ( .A(n_267), .Y(n_288) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_269), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_271), .A2(n_280), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AOI21xp5_ASAP7_75t_SL g490 ( .A1(n_281), .A2(n_491), .B(n_492), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_295), .B1(n_296), .B2(n_301), .C(n_303), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_285), .B(n_287), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_285), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g304 ( .A(n_286), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_286), .A2(n_392), .B(n_393), .C(n_394), .Y(n_391) );
AND2x2_ASAP7_75t_L g396 ( .A(n_286), .B(n_376), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_SL g434 ( .A1(n_286), .A2(n_375), .B(n_435), .C(n_436), .Y(n_434) );
BUFx3_ASAP7_75t_L g326 ( .A(n_287), .Y(n_326) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_290), .B(n_347), .Y(n_390) );
AOI211xp5_ASAP7_75t_L g409 ( .A1(n_290), .A2(n_410), .B(n_412), .C(n_418), .Y(n_409) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVxp67_ASAP7_75t_L g370 ( .A(n_292), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_294), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
AOI211xp5_ASAP7_75t_L g314 ( .A1(n_298), .A2(n_315), .B(n_316), .C(n_324), .Y(n_314) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g399 ( .A(n_302), .Y(n_399) );
OR2x2_ASAP7_75t_L g416 ( .A(n_302), .B(n_346), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_310), .B2(n_313), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_305), .A2(n_317), .B1(n_318), .B2(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
OR2x2_ASAP7_75t_L g403 ( .A(n_307), .B(n_347), .Y(n_403) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g358 ( .A(n_308), .B(n_348), .Y(n_358) );
INVx1_ASAP7_75t_L g366 ( .A(n_309), .Y(n_366) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_312), .B(n_326), .Y(n_374) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_322), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g431 ( .A(n_323), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B(n_330), .Y(n_324) );
INVx1_ASAP7_75t_L g361 ( .A(n_325), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_326), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_326), .B(n_357), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_326), .B(n_352), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_326), .B(n_373), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g388 ( .A1(n_326), .A2(n_336), .B(n_376), .C(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_336), .B1(n_338), .B2(n_342), .C(n_343), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_340), .B(n_348), .Y(n_422) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g433 ( .A1(n_342), .A2(n_357), .B(n_359), .C(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_345), .B(n_352), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_346), .B(n_399), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_347), .Y(n_346) );
INVxp33_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
AOI21xp33_ASAP7_75t_SL g362 ( .A1(n_351), .A2(n_363), .B(n_365), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_351), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_352), .B(n_406), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_359), .B2(n_361), .C(n_362), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_358), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
NAND5xp2_ASAP7_75t_L g367 ( .A(n_368), .B(n_395), .C(n_409), .D(n_420), .E(n_433), .Y(n_367) );
AOI211xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B(n_378), .C(n_391), .Y(n_368) );
INVx2_ASAP7_75t_SL g415 ( .A(n_369), .Y(n_415) );
NAND4xp25_ASAP7_75t_SL g371 ( .A(n_372), .B(n_374), .C(n_375), .D(n_377), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_377), .A2(n_379), .B(n_382), .C(n_388), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_380), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_421), .B1(n_423), .B2(n_425), .C(n_427), .Y(n_420) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI221xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B1(n_400), .B2(n_402), .C(n_404), .Y(n_395) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_403), .A2(n_426), .B1(n_428), .B2(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx4_ASAP7_75t_L g732 ( .A(n_441), .Y(n_732) );
XOR2xp5_ASAP7_75t_L g742 ( .A(n_441), .B(n_743), .Y(n_742) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR5x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_599), .C(n_677), .D(n_701), .E(n_718), .Y(n_442) );
OAI211xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_476), .B(n_518), .C(n_576), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_455), .Y(n_444) );
AND2x2_ASAP7_75t_L g530 ( .A(n_445), .B(n_457), .Y(n_530) );
INVx5_ASAP7_75t_SL g558 ( .A(n_445), .Y(n_558) );
AND2x2_ASAP7_75t_L g594 ( .A(n_445), .B(n_579), .Y(n_594) );
OR2x2_ASAP7_75t_L g633 ( .A(n_445), .B(n_456), .Y(n_633) );
OR2x2_ASAP7_75t_L g664 ( .A(n_445), .B(n_555), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_445), .B(n_568), .Y(n_700) );
AND2x2_ASAP7_75t_L g712 ( .A(n_445), .B(n_555), .Y(n_712) );
OR2x6_ASAP7_75t_L g445 ( .A(n_446), .B(n_454), .Y(n_445) );
AND2x2_ASAP7_75t_L g711 ( .A(n_455), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g574 ( .A(n_456), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_466), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_457), .B(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_457), .Y(n_567) );
INVx3_ASAP7_75t_L g582 ( .A(n_457), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_457), .B(n_466), .Y(n_606) );
OR2x2_ASAP7_75t_L g615 ( .A(n_457), .B(n_558), .Y(n_615) );
AND2x2_ASAP7_75t_L g619 ( .A(n_457), .B(n_579), .Y(n_619) );
AND2x2_ASAP7_75t_L g625 ( .A(n_457), .B(n_626), .Y(n_625) );
INVxp67_ASAP7_75t_L g662 ( .A(n_457), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_457), .B(n_521), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_462), .A2(n_503), .B(n_504), .C(n_505), .Y(n_502) );
OR2x2_ASAP7_75t_L g568 ( .A(n_466), .B(n_521), .Y(n_568) );
AND2x2_ASAP7_75t_L g579 ( .A(n_466), .B(n_555), .Y(n_579) );
AND2x2_ASAP7_75t_L g591 ( .A(n_466), .B(n_582), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_466), .B(n_521), .Y(n_614) );
INVx1_ASAP7_75t_SL g626 ( .A(n_466), .Y(n_626) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g520 ( .A(n_467), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_467), .B(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .B(n_475), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_475), .A2(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
AND2x2_ASAP7_75t_L g539 ( .A(n_478), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_478), .B(n_498), .Y(n_543) );
AND2x2_ASAP7_75t_L g546 ( .A(n_478), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_478), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_562), .Y(n_571) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_478), .Y(n_590) );
AND2x2_ASAP7_75t_L g611 ( .A(n_478), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g621 ( .A(n_478), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g667 ( .A(n_478), .B(n_550), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_478), .B(n_573), .Y(n_694) );
INVx5_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g564 ( .A(n_479), .Y(n_564) );
AND2x2_ASAP7_75t_L g630 ( .A(n_479), .B(n_562), .Y(n_630) );
AND2x2_ASAP7_75t_L g714 ( .A(n_479), .B(n_582), .Y(n_714) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_488), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_488), .Y(n_703) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_498), .Y(n_488) );
AND2x2_ASAP7_75t_L g533 ( .A(n_489), .B(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g542 ( .A(n_489), .B(n_540), .Y(n_542) );
INVx5_ASAP7_75t_L g550 ( .A(n_489), .Y(n_550) );
AND2x2_ASAP7_75t_L g573 ( .A(n_489), .B(n_509), .Y(n_573) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_489), .Y(n_610) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_496), .Y(n_489) );
INVx1_ASAP7_75t_L g651 ( .A(n_498), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_498), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g684 ( .A(n_498), .B(n_550), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_498), .A2(n_607), .B(n_714), .C(n_715), .Y(n_713) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_509), .Y(n_498) );
BUFx2_ASAP7_75t_L g534 ( .A(n_499), .Y(n_534) );
INVx2_ASAP7_75t_L g538 ( .A(n_499), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
INVx2_ASAP7_75t_L g540 ( .A(n_509), .Y(n_540) );
AND2x2_ASAP7_75t_L g547 ( .A(n_509), .B(n_538), .Y(n_547) );
AND2x2_ASAP7_75t_L g638 ( .A(n_509), .B(n_550), .Y(n_638) );
AOI211x1_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_531), .B(n_544), .C(n_569), .Y(n_518) );
INVx1_ASAP7_75t_L g635 ( .A(n_519), .Y(n_635) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_530), .Y(n_519) );
INVx5_ASAP7_75t_SL g555 ( .A(n_521), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_521), .B(n_625), .Y(n_624) );
AOI311xp33_ASAP7_75t_L g643 ( .A1(n_521), .A2(n_644), .A3(n_646), .B(n_647), .C(n_653), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_521), .A2(n_591), .B(n_679), .C(n_682), .Y(n_678) );
INVxp67_ASAP7_75t_L g598 ( .A(n_530), .Y(n_598) );
NAND4xp25_ASAP7_75t_SL g531 ( .A(n_532), .B(n_535), .C(n_541), .D(n_543), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_532), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g589 ( .A(n_533), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_536), .B(n_542), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_536), .B(n_549), .Y(n_669) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_537), .B(n_550), .Y(n_687) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
INVxp67_ASAP7_75t_L g597 ( .A(n_539), .Y(n_597) );
AND2x4_ASAP7_75t_L g549 ( .A(n_540), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g623 ( .A(n_540), .B(n_562), .Y(n_623) );
INVx1_ASAP7_75t_L g650 ( .A(n_540), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_540), .B(n_637), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_541), .B(n_611), .Y(n_631) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_542), .B(n_564), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_542), .B(n_611), .Y(n_710) );
INVx1_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B(n_551), .C(n_559), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g563 ( .A(n_547), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g601 ( .A(n_547), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g583 ( .A(n_548), .Y(n_583) );
AND2x2_ASAP7_75t_L g560 ( .A(n_549), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_549), .B(n_611), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_549), .B(n_630), .Y(n_654) );
OR2x2_ASAP7_75t_L g570 ( .A(n_550), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g602 ( .A(n_550), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_550), .B(n_562), .Y(n_617) );
AND2x2_ASAP7_75t_L g674 ( .A(n_550), .B(n_630), .Y(n_674) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_550), .Y(n_681) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_552), .A2(n_564), .B1(n_686), .B2(n_688), .C(n_691), .Y(n_685) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g575 ( .A(n_555), .B(n_558), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_555), .B(n_625), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_555), .B(n_582), .Y(n_690) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g675 ( .A(n_557), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g689 ( .A(n_557), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_558), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g586 ( .A(n_558), .B(n_579), .Y(n_586) );
AND2x2_ASAP7_75t_L g656 ( .A(n_558), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_558), .B(n_605), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_558), .B(n_706), .Y(n_705) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_563), .B(n_565), .Y(n_559) );
INVx2_ASAP7_75t_L g592 ( .A(n_560), .Y(n_592) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g612 ( .A(n_562), .Y(n_612) );
OR2x2_ASAP7_75t_L g616 ( .A(n_564), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g719 ( .A(n_564), .B(n_687), .Y(n_719) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AOI21xp33_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_572), .B(n_574), .Y(n_569) );
INVx1_ASAP7_75t_L g723 ( .A(n_570), .Y(n_723) );
INVx2_ASAP7_75t_SL g637 ( .A(n_571), .Y(n_637) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_574), .A2(n_655), .B(n_719), .C(n_720), .Y(n_718) );
OAI322xp33_ASAP7_75t_SL g587 ( .A1(n_575), .A2(n_588), .A3(n_591), .B1(n_592), .B2(n_593), .C1(n_595), .C2(n_598), .Y(n_587) );
INVx2_ASAP7_75t_L g607 ( .A(n_575), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_583), .B1(n_584), .B2(n_586), .C(n_587), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp33_ASAP7_75t_SL g653 ( .A1(n_578), .A2(n_654), .B1(n_655), .B2(n_658), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_579), .B(n_582), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_579), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g652 ( .A(n_581), .B(n_614), .Y(n_652) );
INVx1_ASAP7_75t_L g642 ( .A(n_582), .Y(n_642) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_586), .A2(n_696), .B(n_698), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_588), .A2(n_621), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp67_ASAP7_75t_SL g649 ( .A(n_590), .B(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_590), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g706 ( .A(n_591), .Y(n_706) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND4xp25_ASAP7_75t_L g599 ( .A(n_600), .B(n_627), .C(n_643), .D(n_659), .Y(n_599) );
AOI211xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .B(n_608), .C(n_620), .Y(n_600) );
INVx1_ASAP7_75t_L g692 ( .A(n_601), .Y(n_692) );
AND2x2_ASAP7_75t_L g640 ( .A(n_602), .B(n_623), .Y(n_640) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_607), .B(n_642), .Y(n_641) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_613), .B1(n_616), .B2(n_618), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_610), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g658 ( .A(n_611), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_611), .A2(n_650), .B(n_673), .C(n_675), .Y(n_672) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g657 ( .A(n_614), .Y(n_657) );
INVx1_ASAP7_75t_L g717 ( .A(n_615), .Y(n_717) );
NAND2xp33_ASAP7_75t_SL g707 ( .A(n_616), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g646 ( .A(n_625), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_631), .B(n_632), .C(n_634), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_639), .B2(n_641), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_637), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_642), .B(n_663), .Y(n_725) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI21xp33_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_651), .B(n_652), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_665), .B1(n_668), .B2(n_670), .C(n_672), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_675), .A2(n_692), .B1(n_693), .B2(n_694), .Y(n_691) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_685), .C(n_695), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_704), .C(n_713), .Y(n_701) );
INVx1_ASAP7_75t_L g722 ( .A(n_702), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B1(n_709), .B2(n_711), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g749 ( .A(n_739), .Y(n_749) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_746), .Y(n_741) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g753 ( .A(n_747), .Y(n_753) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule