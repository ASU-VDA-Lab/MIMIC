module fake_ariane_1778_n_2382 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_297, n_503, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_231, n_366, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_514, n_418, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_2382);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_297;
input n_503;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_514;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;

output n_2382;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_1703;
wire n_899;
wire n_2332;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_533;
wire n_1917;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_976;
wire n_712;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_2180;
wire n_1942;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_2101;
wire n_1934;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_548;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g526 ( 
.A(n_247),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_21),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_489),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_92),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_435),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_510),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_189),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_60),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_424),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_194),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_325),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_60),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_241),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_466),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_395),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_462),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_391),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_472),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_338),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_432),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_26),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_193),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_187),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_499),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_119),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_32),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_520),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_518),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_242),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_129),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_356),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_144),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_216),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_457),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_231),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_524),
.Y(n_562)
);

CKINVDCx14_ASAP7_75t_R g563 ( 
.A(n_128),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_449),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_15),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_247),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_124),
.Y(n_567)
);

BUFx2_ASAP7_75t_SL g568 ( 
.A(n_74),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_496),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_458),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_3),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_144),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_446),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_186),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_365),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_500),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_211),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_337),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_0),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_376),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_64),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_181),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_49),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_223),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_305),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_508),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_212),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_289),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_212),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_249),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_423),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_380),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_201),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_228),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_451),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_88),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_372),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_369),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_222),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_319),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_126),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_331),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_157),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_146),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_521),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_155),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_260),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_450),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_350),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_218),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_513),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_504),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_36),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_314),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_124),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_285),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_221),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_321),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_162),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_278),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_204),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_11),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_113),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_430),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_62),
.Y(n_626)
);

BUFx5_ASAP7_75t_L g627 ( 
.A(n_502),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_268),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_100),
.Y(n_629)
);

CKINVDCx16_ASAP7_75t_R g630 ( 
.A(n_503),
.Y(n_630)
);

BUFx8_ASAP7_75t_SL g631 ( 
.A(n_256),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_418),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_208),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_228),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_90),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_127),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_377),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_511),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_269),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_320),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_133),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_154),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_101),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_514),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_238),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_517),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_437),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_273),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_90),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_57),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_401),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_515),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_371),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_87),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_434),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_308),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_525),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_80),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_189),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_222),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_342),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_326),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_484),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_431),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_102),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_202),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_519),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_51),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_133),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_246),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_94),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_501),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_158),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_307),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_522),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_444),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_160),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_217),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_69),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_20),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_438),
.Y(n_681)
);

CKINVDCx14_ASAP7_75t_R g682 ( 
.A(n_47),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_304),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_394),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_99),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_313),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_306),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_523),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_127),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_346),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_261),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_385),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_147),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_136),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_382),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_99),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_13),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_44),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_142),
.Y(n_699)
);

CKINVDCx14_ASAP7_75t_R g700 ( 
.A(n_267),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_101),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_311),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_27),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_9),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_452),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_104),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_126),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_400),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_23),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_192),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_355),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_272),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_440),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_38),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_498),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_251),
.Y(n_716)
);

CKINVDCx16_ASAP7_75t_R g717 ( 
.A(n_287),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_351),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_288),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_378),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_516),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_509),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_96),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_512),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_387),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_18),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_197),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_505),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_317),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_145),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_167),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_209),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_26),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_412),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_493),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_507),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_231),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_105),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_29),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_468),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_125),
.Y(n_741)
);

CKINVDCx16_ASAP7_75t_R g742 ( 
.A(n_153),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_159),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_65),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_448),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_716),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_716),
.Y(n_747)
);

INVxp33_ASAP7_75t_SL g748 ( 
.A(n_672),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_577),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_577),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_563),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_604),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_563),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_604),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_697),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_697),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_701),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_701),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_526),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_532),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_547),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_682),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_682),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_552),
.Y(n_764)
);

INVxp33_ASAP7_75t_SL g765 ( 
.A(n_665),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_556),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_559),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_551),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_565),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_574),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_551),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_700),
.Y(n_772)
);

CKINVDCx16_ASAP7_75t_R g773 ( 
.A(n_700),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_598),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_558),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_744),
.B(n_0),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_631),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_583),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_608),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_618),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_558),
.Y(n_781)
);

INVxp33_ASAP7_75t_SL g782 ( 
.A(n_527),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_628),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_631),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_592),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_635),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_642),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_643),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_650),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_630),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_551),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_660),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_668),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_677),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_703),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_706),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_709),
.Y(n_797)
);

INVxp33_ASAP7_75t_L g798 ( 
.A(n_593),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_733),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_741),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_640),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_593),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_611),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_611),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_551),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_605),
.B(n_1),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_670),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_670),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_685),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_546),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_685),
.Y(n_811)
);

CKINVDCx16_ASAP7_75t_R g812 ( 
.A(n_717),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_738),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_657),
.Y(n_814)
);

INVxp33_ASAP7_75t_L g815 ( 
.A(n_738),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_738),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_738),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_589),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_529),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_671),
.Y(n_820)
);

INVxp33_ASAP7_75t_SL g821 ( 
.A(n_533),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_673),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_531),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_568),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_598),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_694),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_579),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_742),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_591),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_603),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_591),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_591),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_736),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_736),
.Y(n_834)
);

INVxp33_ASAP7_75t_SL g835 ( 
.A(n_535),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_603),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_647),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_543),
.Y(n_839)
);

OR2x2_ASAP7_75t_L g840 ( 
.A(n_581),
.B(n_1),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_579),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_579),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_798),
.B(n_679),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_838),
.B(n_530),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_768),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_748),
.A2(n_531),
.B1(n_725),
.B2(n_595),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_810),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_771),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_798),
.B(n_679),
.Y(n_849)
);

INVx5_ASAP7_75t_L g850 ( 
.A(n_810),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_839),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_828),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_774),
.B(n_647),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_829),
.B(n_536),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_810),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_774),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_810),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_813),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_816),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_775),
.Y(n_860)
);

BUFx8_ASAP7_75t_SL g861 ( 
.A(n_775),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_831),
.B(n_539),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_791),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_832),
.B(n_540),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_773),
.B(n_679),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_776),
.B(n_615),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_805),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_817),
.Y(n_868)
);

AOI22x1_ASAP7_75t_SL g869 ( 
.A1(n_823),
.A2(n_648),
.B1(n_678),
.B2(n_602),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_751),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_825),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_833),
.B(n_541),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_830),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_830),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_837),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_785),
.B(n_595),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_834),
.B(n_836),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_823),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_746),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_747),
.A2(n_553),
.B(n_544),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_785),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_790),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_748),
.A2(n_648),
.B1(n_678),
.B2(n_602),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_759),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_837),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_825),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_760),
.Y(n_887)
);

AND2x2_ASAP7_75t_SL g888 ( 
.A(n_840),
.B(n_615),
.Y(n_888)
);

XNOR2xp5_ASAP7_75t_L g889 ( 
.A(n_781),
.B(n_567),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_802),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_765),
.A2(n_728),
.B1(n_725),
.B2(n_584),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_749),
.Y(n_892)
);

XNOR2x2_ASAP7_75t_L g893 ( 
.A(n_781),
.B(n_594),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_815),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_803),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_752),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_750),
.B(n_664),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_761),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_764),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_804),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_754),
.B(n_730),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_784),
.Y(n_902)
);

CKINVDCx16_ASAP7_75t_R g903 ( 
.A(n_812),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_751),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_841),
.B(n_664),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_753),
.B(n_564),
.Y(n_906)
);

OA21x2_ASAP7_75t_L g907 ( 
.A1(n_807),
.A2(n_596),
.B(n_573),
.Y(n_907)
);

INVx4_ASAP7_75t_L g908 ( 
.A(n_875),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_875),
.Y(n_909)
);

OAI21x1_ASAP7_75t_L g910 ( 
.A1(n_880),
.A2(n_609),
.B(n_599),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_874),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_875),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_875),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_875),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_888),
.A2(n_728),
.B1(n_765),
.B2(n_732),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_880),
.A2(n_719),
.B(n_613),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_885),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_851),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_874),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_855),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_858),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_885),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_858),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_866),
.B(n_753),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_851),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_843),
.B(n_755),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_885),
.Y(n_927)
);

AND2x2_ASAP7_75t_SL g928 ( 
.A(n_866),
.B(n_719),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_885),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_885),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_868),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_868),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_873),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_873),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_904),
.B(n_790),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_873),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_907),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_873),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_907),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_907),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_857),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_888),
.B(n_762),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_897),
.B(n_762),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_857),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_904),
.B(n_782),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_903),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_859),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_856),
.B(n_842),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_859),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_877),
.A2(n_801),
.B1(n_814),
.B2(n_782),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_900),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_843),
.Y(n_952)
);

AND2x6_ASAP7_75t_L g953 ( 
.A(n_901),
.B(n_686),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_900),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_861),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_900),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_855),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_886),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_900),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_859),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_859),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_890),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_890),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_895),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_SL g965 ( 
.A(n_870),
.B(n_777),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_895),
.Y(n_966)
);

OA21x2_ASAP7_75t_L g967 ( 
.A1(n_844),
.A2(n_637),
.B(n_610),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_879),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_845),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_878),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_848),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_855),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_878),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_870),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_847),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_847),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_881),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_L g978 ( 
.A(n_881),
.B(n_882),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_849),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_847),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_847),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_863),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_867),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_886),
.B(n_819),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_856),
.B(n_827),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_882),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_850),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_876),
.Y(n_988)
);

CKINVDCx8_ASAP7_75t_R g989 ( 
.A(n_897),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_850),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_849),
.B(n_756),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_897),
.B(n_763),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_850),
.Y(n_993)
);

BUFx6f_ASAP7_75t_SL g994 ( 
.A(n_905),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_886),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_850),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_952),
.B(n_852),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_994),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_928),
.B(n_901),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_911),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_911),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_928),
.B(n_854),
.Y(n_1002)
);

BUFx10_ASAP7_75t_L g1003 ( 
.A(n_918),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_SL g1004 ( 
.A1(n_928),
.A2(n_883),
.B1(n_893),
.B2(n_869),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_919),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_952),
.B(n_906),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_979),
.A2(n_814),
.B1(n_801),
.B2(n_846),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_918),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_968),
.A2(n_821),
.B(n_819),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_919),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_969),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_969),
.A2(n_971),
.B1(n_983),
.B2(n_982),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_971),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_953),
.Y(n_1014)
);

INVx4_ASAP7_75t_L g1015 ( 
.A(n_994),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_974),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_989),
.B(n_821),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_974),
.B(n_865),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_982),
.A2(n_853),
.B1(n_865),
.B2(n_562),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_983),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_968),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_921),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_962),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_915),
.A2(n_953),
.B1(n_926),
.B2(n_991),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_964),
.B(n_862),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_915),
.A2(n_891),
.B1(n_731),
.B2(n_636),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_950),
.A2(n_587),
.B1(n_835),
.B2(n_806),
.Y(n_1027)
);

OAI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_989),
.A2(n_924),
.B1(n_942),
.B2(n_925),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_977),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_962),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_977),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_921),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_986),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_923),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_923),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_986),
.B(n_889),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_946),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_985),
.B(n_871),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_931),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_931),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_932),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_963),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_963),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_948),
.B(n_871),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_985),
.B(n_871),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_970),
.B(n_777),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_932),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_964),
.B(n_966),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_994),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_941),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_941),
.Y(n_1051)
);

OAI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_943),
.A2(n_864),
.B1(n_872),
.B2(n_824),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_958),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_955),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_945),
.B(n_835),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_988),
.B(n_763),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_966),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_944),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_973),
.B(n_902),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_951),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_953),
.A2(n_967),
.B1(n_991),
.B2(n_926),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_955),
.Y(n_1063)
);

BUFx10_ASAP7_75t_L g1064 ( 
.A(n_985),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_935),
.B(n_772),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_985),
.B(n_853),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_958),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_948),
.B(n_853),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_920),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_992),
.B(n_772),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_984),
.B(n_784),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_948),
.B(n_886),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_965),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_920),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_948),
.B(n_905),
.Y(n_1075)
);

INVx6_ASAP7_75t_L g1076 ( 
.A(n_956),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_956),
.Y(n_1077)
);

NAND2xp33_ASAP7_75t_L g1078 ( 
.A(n_920),
.B(n_537),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_995),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_951),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_954),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_957),
.A2(n_887),
.B1(n_898),
.B2(n_884),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_954),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_959),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_978),
.B(n_905),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_957),
.B(n_892),
.Y(n_1086)
);

INVxp33_ASAP7_75t_L g1087 ( 
.A(n_967),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_953),
.B(n_899),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_953),
.B(n_892),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_933),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_957),
.B(n_896),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_959),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_933),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_972),
.B(n_894),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_995),
.B(n_889),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_972),
.B(n_894),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_953),
.B(n_896),
.Y(n_1097)
);

AND2x6_ASAP7_75t_L g1098 ( 
.A(n_937),
.B(n_686),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_953),
.B(n_894),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_956),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_972),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_947),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_967),
.Y(n_1103)
);

AND3x2_ASAP7_75t_L g1104 ( 
.A(n_947),
.B(n_861),
.C(n_860),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_949),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_967),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_956),
.Y(n_1107)
);

INVxp67_ASAP7_75t_SL g1108 ( 
.A(n_912),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_995),
.B(n_894),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_934),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_934),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_949),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_937),
.B(n_894),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_960),
.B(n_766),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_956),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_975),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_960),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_936),
.B(n_893),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_936),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_908),
.B(n_538),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_975),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_938),
.Y(n_1122)
);

INVx6_ASAP7_75t_L g1123 ( 
.A(n_961),
.Y(n_1123)
);

AND2x2_ASAP7_75t_SL g1124 ( 
.A(n_916),
.B(n_860),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_938),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_909),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_939),
.B(n_676),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_975),
.Y(n_1128)
);

OAI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_939),
.A2(n_549),
.B(n_548),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_909),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_908),
.A2(n_726),
.B1(n_696),
.B2(n_555),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_922),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_940),
.B(n_638),
.Y(n_1133)
);

OAI21xp33_ASAP7_75t_SL g1134 ( 
.A1(n_910),
.A2(n_769),
.B(n_767),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_981),
.B(n_757),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1011),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1005),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1012),
.B(n_940),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_998),
.B(n_770),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1013),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_L g1141 ( 
.A(n_1027),
.B(n_566),
.C(n_561),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_998),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1026),
.A2(n_922),
.B1(n_929),
.B2(n_730),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1050),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1053),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1085),
.A2(n_910),
.B(n_929),
.C(n_981),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1029),
.B(n_908),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1029),
.B(n_908),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1020),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1021),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_1016),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1002),
.B(n_912),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1033),
.B(n_912),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1002),
.B(n_912),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1033),
.B(n_912),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_1018),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1031),
.B(n_758),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_999),
.B(n_913),
.Y(n_1158)
);

OAI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1026),
.A2(n_571),
.B1(n_590),
.B2(n_572),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_1055),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1017),
.B(n_1028),
.Y(n_1161)
);

NOR2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1008),
.B(n_778),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1051),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1004),
.A2(n_730),
.B1(n_961),
.B2(n_740),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1135),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1048),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_999),
.B(n_913),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1027),
.B(n_624),
.C(n_614),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1064),
.B(n_913),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1015),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1054),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1048),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1114),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1024),
.B(n_913),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_1015),
.B(n_961),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1024),
.B(n_1025),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1009),
.A2(n_818),
.B(n_822),
.C(n_820),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_1049),
.B(n_779),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1009),
.B(n_914),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1064),
.B(n_913),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1114),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1068),
.B(n_914),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1025),
.B(n_914),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1052),
.B(n_914),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1056),
.B(n_917),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1059),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1037),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1070),
.B(n_914),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1004),
.A2(n_961),
.B1(n_740),
.B2(n_927),
.Y(n_1189)
);

BUFx5_ASAP7_75t_L g1190 ( 
.A(n_1101),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1006),
.B(n_917),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1023),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1030),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1042),
.Y(n_1194)
);

INVx8_ASAP7_75t_L g1195 ( 
.A(n_1066),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1060),
.B(n_815),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1082),
.B(n_1086),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1082),
.B(n_917),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1036),
.B(n_917),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1068),
.B(n_917),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1049),
.B(n_780),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1043),
.Y(n_1202)
);

NAND2xp33_ASAP7_75t_L g1203 ( 
.A(n_1069),
.B(n_927),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1057),
.B(n_783),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_997),
.B(n_927),
.Y(n_1205)
);

NOR2xp67_ASAP7_75t_L g1206 ( 
.A(n_1063),
.B(n_786),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1044),
.B(n_927),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1095),
.B(n_787),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1091),
.B(n_927),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1044),
.B(n_930),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1003),
.B(n_788),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_SL g1212 ( 
.A(n_1003),
.B(n_542),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1066),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1072),
.B(n_930),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1073),
.B(n_930),
.Y(n_1215)
);

NAND2xp33_ASAP7_75t_L g1216 ( 
.A(n_1069),
.B(n_930),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1053),
.Y(n_1217)
);

AO22x2_ASAP7_75t_L g1218 ( 
.A1(n_1118),
.A2(n_826),
.B1(n_809),
.B2(n_811),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1053),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1061),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1007),
.B(n_789),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1089),
.B(n_930),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1080),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1000),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1022),
.B(n_961),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1032),
.B(n_981),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1046),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1034),
.B(n_976),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1035),
.B(n_1039),
.Y(n_1229)
);

OR2x2_ASAP7_75t_SL g1230 ( 
.A(n_1104),
.B(n_792),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1001),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1066),
.B(n_793),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1081),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1040),
.B(n_976),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1041),
.B(n_980),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1047),
.B(n_980),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1058),
.B(n_582),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1075),
.B(n_597),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1074),
.B(n_600),
.Y(n_1239)
);

OAI21xp33_ASAP7_75t_L g1240 ( 
.A1(n_1129),
.A2(n_633),
.B(n_621),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1019),
.B(n_794),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1124),
.A2(n_729),
.B1(n_651),
.B2(n_656),
.Y(n_1242)
);

NOR2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1089),
.B(n_795),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1074),
.B(n_607),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1014),
.B(n_987),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1083),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1010),
.B(n_616),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1131),
.A2(n_675),
.B1(n_690),
.B2(n_646),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1084),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1131),
.A2(n_705),
.B1(n_711),
.B2(n_692),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1038),
.B(n_796),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1014),
.B(n_987),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1065),
.B(n_617),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_L g1254 ( 
.A(n_1014),
.B(n_990),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1122),
.B(n_620),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1092),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1129),
.B(n_622),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1067),
.B(n_990),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1062),
.B(n_623),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1071),
.B(n_626),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1133),
.B(n_797),
.Y(n_1261)
);

BUFx5_ASAP7_75t_L g1262 ( 
.A(n_1098),
.Y(n_1262)
);

NOR2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1116),
.B(n_799),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1079),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1045),
.A2(n_724),
.B1(n_734),
.B2(n_720),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1067),
.B(n_800),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_L g1267 ( 
.A(n_1078),
.B(n_1120),
.C(n_634),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1127),
.B(n_629),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1128),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1067),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1102),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1076),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1105),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1127),
.B(n_639),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1121),
.B(n_641),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1106),
.A2(n_645),
.B1(n_654),
.B2(n_649),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1088),
.B(n_658),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1112),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1125),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1076),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1126),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1121),
.B(n_659),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1088),
.B(n_993),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1130),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1097),
.B(n_993),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_SL g1286 ( 
.A(n_1097),
.B(n_996),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1077),
.B(n_996),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1098),
.B(n_1132),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1106),
.A2(n_689),
.B(n_707),
.C(n_669),
.Y(n_1289)
);

CKINVDCx20_ASAP7_75t_R g1290 ( 
.A(n_1123),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1090),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1117),
.B(n_666),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1098),
.B(n_680),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1115),
.B(n_691),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1133),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1093),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1098),
.B(n_693),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1110),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1111),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1119),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1115),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1123),
.A2(n_699),
.B1(n_704),
.B2(n_698),
.Y(n_1302)
);

AOI221x1_ASAP7_75t_L g1303 ( 
.A1(n_1113),
.A2(n_808),
.B1(n_653),
.B2(n_687),
.C(n_575),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1077),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1100),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1103),
.B(n_710),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1109),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1100),
.B(n_712),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1107),
.B(n_714),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_1094),
.B(n_1096),
.C(n_1107),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1099),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1103),
.B(n_723),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1108),
.B(n_727),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1099),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1113),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1087),
.B(n_737),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1134),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1011),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1026),
.A2(n_743),
.B1(n_739),
.B2(n_722),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1031),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1011),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1085),
.B(n_528),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1011),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_R g1324 ( 
.A(n_1055),
.B(n_534),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1085),
.B(n_545),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1002),
.A2(n_713),
.B1(n_619),
.B2(n_667),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1012),
.B(n_916),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1053),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1085),
.B(n_550),
.Y(n_1329)
);

BUFx5_ASAP7_75t_L g1330 ( 
.A(n_1101),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1011),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1005),
.Y(n_1332)
);

AO221x1_ASAP7_75t_L g1333 ( 
.A1(n_1026),
.A2(n_653),
.B1(n_687),
.B2(n_575),
.C(n_546),
.Y(n_1333)
);

BUFx6f_ASAP7_75t_L g1334 ( 
.A(n_1053),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1004),
.A2(n_554),
.B1(n_560),
.B2(n_557),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1012),
.B(n_916),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1212),
.B(n_569),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1161),
.B(n_570),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1187),
.B(n_576),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1295),
.B(n_916),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1243),
.B(n_850),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1136),
.Y(n_1342)
);

BUFx4f_ASAP7_75t_L g1343 ( 
.A(n_1195),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1140),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1149),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1260),
.B(n_578),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1151),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1147),
.B(n_1148),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1150),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1220),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1166),
.B(n_2),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1141),
.B(n_585),
.C(n_580),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1318),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1172),
.B(n_2),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1335),
.A2(n_575),
.B1(n_653),
.B2(n_546),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1304),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1320),
.B(n_745),
.Y(n_1357)
);

INVx4_ASAP7_75t_L g1358 ( 
.A(n_1195),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1159),
.B(n_586),
.Y(n_1359)
);

AND2x6_ASAP7_75t_SL g1360 ( 
.A(n_1160),
.B(n_3),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1321),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1319),
.A2(n_1189),
.B1(n_1164),
.B2(n_1181),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1227),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1165),
.B(n_4),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1145),
.Y(n_1365)
);

AO22x1_ASAP7_75t_L g1366 ( 
.A1(n_1270),
.A2(n_601),
.B1(n_606),
.B2(n_588),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1199),
.B(n_4),
.Y(n_1367)
);

OR2x6_ASAP7_75t_L g1368 ( 
.A(n_1139),
.B(n_546),
.Y(n_1368)
);

A2O1A1Ixp33_ASAP7_75t_SL g1369 ( 
.A1(n_1275),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1173),
.A2(n_653),
.B1(n_687),
.B2(n_575),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1176),
.B(n_1156),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1196),
.B(n_5),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1304),
.Y(n_1373)
);

NAND2xp33_ASAP7_75t_SL g1374 ( 
.A(n_1197),
.B(n_612),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1204),
.B(n_6),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1323),
.B(n_7),
.Y(n_1376)
);

BUFx4f_ASAP7_75t_L g1377 ( 
.A(n_1139),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1315),
.A2(n_632),
.B(n_625),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_SL g1379 ( 
.A1(n_1168),
.A2(n_735),
.B1(n_652),
.B2(n_655),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1145),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1331),
.B(n_8),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1224),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1290),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1253),
.B(n_644),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1223),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_SL g1386 ( 
.A(n_1289),
.B(n_662),
.C(n_661),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1208),
.B(n_663),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1185),
.B(n_674),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1162),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1241),
.B(n_8),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1142),
.B(n_9),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1232),
.B(n_10),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1211),
.B(n_681),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1232),
.B(n_10),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1248),
.A2(n_687),
.B1(n_683),
.B2(n_684),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1233),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_L g1397 ( 
.A(n_1178),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1246),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1250),
.A2(n_1326),
.B1(n_1242),
.B2(n_1143),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1157),
.Y(n_1400)
);

INVx5_ASAP7_75t_L g1401 ( 
.A(n_1178),
.Y(n_1401)
);

AO21x1_ASAP7_75t_L g1402 ( 
.A1(n_1198),
.A2(n_627),
.B(n_291),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1324),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1218),
.B(n_11),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1201),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1218),
.B(n_1266),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_SL g1407 ( 
.A(n_1276),
.B(n_695),
.C(n_688),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1231),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1201),
.B(n_12),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1206),
.B(n_702),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1155),
.B(n_721),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1215),
.B(n_708),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1229),
.A2(n_1249),
.B1(n_1256),
.B2(n_1183),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1266),
.B(n_12),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1142),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1137),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1213),
.B(n_715),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1332),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1261),
.B(n_13),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1145),
.B(n_718),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1281),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1219),
.B(n_627),
.Y(n_1422)
);

OAI22x1_ASAP7_75t_SL g1423 ( 
.A1(n_1170),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1423)
);

NAND2x1_ASAP7_75t_L g1424 ( 
.A(n_1304),
.B(n_290),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1284),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1271),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1170),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1144),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1268),
.B(n_14),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1263),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1274),
.B(n_16),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_L g1432 ( 
.A(n_1272),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1273),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1230),
.Y(n_1434)
);

AND2x6_ASAP7_75t_SL g1435 ( 
.A(n_1292),
.B(n_17),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1251),
.B(n_17),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_SL g1437 ( 
.A(n_1179),
.B(n_627),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1219),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_R g1439 ( 
.A(n_1217),
.B(n_292),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1221),
.B(n_18),
.Y(n_1440)
);

O2A1O1Ixp5_ASAP7_75t_L g1441 ( 
.A1(n_1308),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_1441)
);

AND2x4_ASAP7_75t_SL g1442 ( 
.A(n_1272),
.B(n_19),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1251),
.B(n_22),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1278),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1264),
.B(n_1269),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1219),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1282),
.B(n_22),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_SL g1448 ( 
.A(n_1240),
.B(n_23),
.C(n_24),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1328),
.B(n_627),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1312),
.A2(n_627),
.B1(n_27),
.B2(n_24),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1163),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1209),
.A2(n_294),
.B(n_293),
.Y(n_1452)
);

INVxp33_ASAP7_75t_L g1453 ( 
.A(n_1255),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1205),
.A2(n_627),
.B1(n_29),
.B2(n_25),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1171),
.Y(n_1455)
);

INVx5_ASAP7_75t_L g1456 ( 
.A(n_1328),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1328),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1279),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1333),
.A2(n_1257),
.B1(n_1259),
.B2(n_1192),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1291),
.B(n_25),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1186),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1193),
.A2(n_627),
.B1(n_31),
.B2(n_28),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1294),
.B(n_1237),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1247),
.B(n_28),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1238),
.B(n_1152),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1334),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1280),
.B(n_30),
.Y(n_1467)
);

BUFx6f_ASAP7_75t_L g1468 ( 
.A(n_1334),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1334),
.B(n_30),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1239),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1194),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1154),
.B(n_31),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1202),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1272),
.B(n_32),
.Y(n_1474)
);

NAND2x2_ASAP7_75t_L g1475 ( 
.A(n_1244),
.B(n_33),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1174),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1138),
.B(n_34),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1322),
.B(n_1325),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1217),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1301),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1329),
.B(n_35),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1298),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1222),
.B(n_36),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1302),
.B(n_37),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1305),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1296),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1203),
.A2(n_296),
.B(n_295),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1188),
.B(n_37),
.Y(n_1488)
);

O2A1O1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1177),
.A2(n_1309),
.B(n_1153),
.C(n_1313),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1299),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1265),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1300),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1228),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1277),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.C(n_42),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1234),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1235),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1311),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1236),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1306),
.B(n_1158),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1167),
.B(n_41),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1226),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1293),
.B(n_42),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1191),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1307),
.B(n_43),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1175),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1225),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1317),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1207),
.B(n_43),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1190),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1184),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1210),
.B(n_45),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1297),
.B(n_46),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1316),
.B(n_47),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1182),
.B(n_48),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1267),
.B(n_1190),
.Y(n_1515)
);

OR2x6_ASAP7_75t_L g1516 ( 
.A(n_1200),
.B(n_48),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1169),
.B(n_49),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1310),
.B(n_50),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1180),
.B(n_50),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1214),
.B(n_51),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1311),
.B(n_52),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1258),
.Y(n_1522)
);

NOR2xp67_ASAP7_75t_L g1523 ( 
.A(n_1314),
.B(n_297),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1314),
.Y(n_1524)
);

OR2x2_ASAP7_75t_SL g1525 ( 
.A(n_1288),
.B(n_52),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1216),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1283),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1190),
.B(n_53),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1336),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1285),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1190),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1190),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1330),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1330),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1330),
.B(n_58),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1245),
.B(n_59),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1286),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1330),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1330),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1262),
.B(n_1327),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1252),
.B(n_1287),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1146),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1254),
.B(n_61),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1262),
.B(n_63),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1262),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1348),
.B(n_1262),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1413),
.B(n_1262),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1371),
.B(n_1303),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1401),
.B(n_63),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1338),
.B(n_1387),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1401),
.B(n_64),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1401),
.B(n_65),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1377),
.B(n_1397),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1377),
.B(n_66),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_SL g1555 ( 
.A(n_1397),
.B(n_66),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1463),
.B(n_67),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_SL g1557 ( 
.A(n_1415),
.B(n_67),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1497),
.B(n_1399),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1497),
.B(n_68),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1346),
.B(n_68),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1400),
.B(n_69),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1497),
.B(n_70),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1393),
.B(n_1440),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1399),
.B(n_70),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1456),
.B(n_71),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1456),
.B(n_71),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1456),
.B(n_72),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1543),
.B(n_72),
.Y(n_1568)
);

NAND2xp33_ASAP7_75t_SL g1569 ( 
.A(n_1427),
.B(n_73),
.Y(n_1569)
);

NAND2xp33_ASAP7_75t_SL g1570 ( 
.A(n_1427),
.B(n_73),
.Y(n_1570)
);

NAND2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1447),
.B(n_74),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1391),
.B(n_75),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1391),
.B(n_75),
.Y(n_1573)
);

NAND2xp33_ASAP7_75t_SL g1574 ( 
.A(n_1386),
.B(n_76),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1347),
.B(n_76),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_SL g1576 ( 
.A(n_1389),
.B(n_1464),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1405),
.B(n_77),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1478),
.B(n_77),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1374),
.B(n_78),
.Y(n_1579)
);

NAND2xp33_ASAP7_75t_SL g1580 ( 
.A(n_1453),
.B(n_78),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1390),
.B(n_79),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_SL g1582 ( 
.A(n_1351),
.B(n_79),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1470),
.B(n_80),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1483),
.B(n_81),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1354),
.B(n_81),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1384),
.B(n_82),
.Y(n_1586)
);

AND2x4_ASAP7_75t_SL g1587 ( 
.A(n_1358),
.B(n_298),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1483),
.B(n_82),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1365),
.B(n_83),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_SL g1590 ( 
.A(n_1358),
.B(n_83),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_SL g1591 ( 
.A(n_1403),
.B(n_84),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1443),
.B(n_1372),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1392),
.B(n_1394),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1365),
.B(n_84),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1365),
.B(n_85),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1495),
.B(n_85),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1380),
.B(n_86),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_SL g1598 ( 
.A(n_1380),
.B(n_86),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_SL g1599 ( 
.A(n_1380),
.B(n_1457),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1341),
.B(n_299),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1457),
.B(n_87),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1429),
.B(n_88),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1457),
.B(n_89),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1468),
.B(n_89),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1468),
.B(n_91),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1468),
.B(n_91),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1378),
.B(n_92),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1517),
.B(n_93),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1409),
.B(n_93),
.Y(n_1609)
);

NAND2xp33_ASAP7_75t_SL g1610 ( 
.A(n_1431),
.B(n_1376),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1496),
.B(n_1344),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1517),
.B(n_94),
.Y(n_1612)
);

NAND2xp33_ASAP7_75t_SL g1613 ( 
.A(n_1381),
.B(n_95),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1519),
.B(n_95),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1519),
.B(n_96),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1342),
.B(n_97),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1345),
.B(n_97),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1349),
.B(n_98),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1353),
.B(n_98),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_SL g1620 ( 
.A(n_1536),
.B(n_100),
.Y(n_1620)
);

NAND2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1535),
.B(n_1430),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1409),
.B(n_102),
.Y(n_1622)
);

NAND2xp33_ASAP7_75t_SL g1623 ( 
.A(n_1439),
.B(n_103),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1536),
.B(n_103),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1521),
.B(n_104),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1485),
.B(n_105),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1341),
.B(n_106),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1409),
.B(n_106),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1356),
.B(n_107),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1356),
.B(n_107),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1373),
.B(n_1465),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1479),
.B(n_300),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1373),
.B(n_108),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1343),
.B(n_108),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1343),
.B(n_109),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1432),
.B(n_1518),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1361),
.B(n_109),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1432),
.B(n_110),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_SL g1639 ( 
.A(n_1379),
.B(n_110),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1524),
.B(n_111),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1382),
.B(n_111),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1438),
.B(n_112),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1408),
.B(n_1493),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1438),
.B(n_112),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1446),
.B(n_113),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1446),
.B(n_114),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1359),
.B(n_114),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1445),
.B(n_115),
.Y(n_1648)
);

AND2x4_ASAP7_75t_SL g1649 ( 
.A(n_1368),
.B(n_1466),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1445),
.B(n_115),
.Y(n_1650)
);

NAND2xp33_ASAP7_75t_SL g1651 ( 
.A(n_1379),
.B(n_116),
.Y(n_1651)
);

NAND2xp33_ASAP7_75t_SL g1652 ( 
.A(n_1467),
.B(n_1364),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1541),
.B(n_116),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1541),
.B(n_117),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1501),
.B(n_117),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1467),
.B(n_118),
.Y(n_1656)
);

NAND2xp33_ASAP7_75t_SL g1657 ( 
.A(n_1436),
.B(n_118),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1466),
.B(n_119),
.Y(n_1658)
);

NAND2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1383),
.B(n_120),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1363),
.B(n_120),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1337),
.B(n_121),
.Y(n_1661)
);

NAND2xp33_ASAP7_75t_SL g1662 ( 
.A(n_1375),
.B(n_121),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_SL g1663 ( 
.A(n_1367),
.B(n_122),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1350),
.B(n_301),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1498),
.B(n_122),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1385),
.B(n_123),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1504),
.B(n_1414),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1489),
.B(n_123),
.Y(n_1668)
);

NAND2xp33_ASAP7_75t_SL g1669 ( 
.A(n_1534),
.B(n_125),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1506),
.B(n_128),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1412),
.B(n_129),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1499),
.B(n_130),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1339),
.B(n_130),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1396),
.B(n_131),
.Y(n_1674)
);

NAND2xp33_ASAP7_75t_SL g1675 ( 
.A(n_1357),
.B(n_131),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1454),
.B(n_132),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1454),
.B(n_132),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1362),
.B(n_134),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1484),
.B(n_134),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1523),
.B(n_135),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1523),
.B(n_135),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1388),
.B(n_136),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1398),
.B(n_137),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1355),
.B(n_137),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1460),
.B(n_138),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_SL g1686 ( 
.A(n_1538),
.B(n_138),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1421),
.B(n_139),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1514),
.B(n_139),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_1425),
.B(n_140),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_SL g1690 ( 
.A(n_1426),
.B(n_140),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1433),
.B(n_141),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1444),
.B(n_141),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1458),
.B(n_142),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1507),
.B(n_1406),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1417),
.B(n_143),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1434),
.B(n_143),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1368),
.B(n_145),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_SL g1698 ( 
.A(n_1520),
.B(n_146),
.Y(n_1698)
);

NAND2xp33_ASAP7_75t_SL g1699 ( 
.A(n_1538),
.B(n_147),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1352),
.B(n_148),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_SL g1701 ( 
.A(n_1513),
.B(n_148),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1526),
.B(n_149),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1526),
.B(n_149),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1505),
.B(n_150),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1477),
.B(n_150),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1411),
.B(n_151),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1419),
.B(n_151),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1509),
.B(n_152),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1404),
.B(n_152),
.Y(n_1709)
);

NAND2xp33_ASAP7_75t_SL g1710 ( 
.A(n_1481),
.B(n_1508),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1544),
.B(n_153),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1476),
.B(n_154),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1486),
.B(n_155),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_SL g1714 ( 
.A(n_1476),
.B(n_156),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1532),
.B(n_156),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1539),
.B(n_157),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1511),
.B(n_158),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1500),
.B(n_159),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1531),
.B(n_160),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1533),
.B(n_161),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1472),
.B(n_161),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_SL g1722 ( 
.A(n_1480),
.B(n_162),
.Y(n_1722)
);

NAND2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1515),
.B(n_163),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1450),
.B(n_163),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1529),
.B(n_164),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1529),
.B(n_164),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1527),
.B(n_165),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1503),
.B(n_165),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1491),
.B(n_1437),
.Y(n_1729)
);

NAND2xp33_ASAP7_75t_SL g1730 ( 
.A(n_1420),
.B(n_166),
.Y(n_1730)
);

NAND2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1474),
.B(n_166),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1522),
.B(n_1340),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1490),
.B(n_302),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1492),
.B(n_167),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1502),
.B(n_168),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1512),
.B(n_168),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1542),
.B(n_1528),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1410),
.B(n_169),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1563),
.A2(n_1448),
.B1(n_1416),
.B2(n_1428),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1592),
.B(n_1442),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1643),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1558),
.B(n_1418),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1561),
.B(n_1516),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1694),
.B(n_1471),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1611),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1616),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1617),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1550),
.B(n_1473),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1732),
.B(n_1451),
.Y(n_1749)
);

OAI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1647),
.A2(n_1510),
.B(n_1494),
.Y(n_1750)
);

AND2x4_ASAP7_75t_SL g1751 ( 
.A(n_1600),
.B(n_1368),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1636),
.B(n_1435),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1564),
.B(n_1455),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1581),
.B(n_1525),
.Y(n_1754)
);

NAND2x1p5_ASAP7_75t_L g1755 ( 
.A(n_1553),
.B(n_1733),
.Y(n_1755)
);

O2A1O1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1560),
.A2(n_1369),
.B(n_1516),
.C(n_1469),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1666),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1674),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1652),
.B(n_1402),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1683),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1621),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1618),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1679),
.B(n_1516),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1619),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1639),
.A2(n_1423),
.B1(n_1407),
.B2(n_1395),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1667),
.B(n_1461),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1713),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1600),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1596),
.B(n_1583),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1637),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1586),
.B(n_1482),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1696),
.B(n_1366),
.Y(n_1772)
);

CKINVDCx16_ASAP7_75t_R g1773 ( 
.A(n_1609),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1649),
.Y(n_1774)
);

BUFx12f_ASAP7_75t_L g1775 ( 
.A(n_1660),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1676),
.A2(n_1459),
.B1(n_1475),
.B2(n_1462),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1641),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1600),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_1591),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1576),
.Y(n_1780)
);

NOR2xp67_ASAP7_75t_L g1781 ( 
.A(n_1575),
.B(n_1452),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1631),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1622),
.B(n_1628),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1548),
.B(n_1488),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1677),
.A2(n_1537),
.B1(n_1530),
.B2(n_1540),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1687),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1593),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1733),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1733),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1608),
.B(n_1360),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1610),
.B(n_1545),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1664),
.Y(n_1792)
);

AND3x1_ASAP7_75t_SL g1793 ( 
.A(n_1659),
.B(n_169),
.C(n_170),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1664),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1651),
.A2(n_1580),
.B1(n_1656),
.B2(n_1623),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1664),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1709),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1599),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1670),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1655),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1546),
.B(n_1422),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1632),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1728),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1649),
.B(n_1449),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1546),
.B(n_1370),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1587),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1587),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1737),
.B(n_1487),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1632),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1632),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1697),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1712),
.A2(n_1424),
.B1(n_1441),
.B2(n_172),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1584),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1612),
.B(n_1614),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1665),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1737),
.B(n_1725),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1723),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1734),
.Y(n_1818)
);

AOI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1714),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1726),
.B(n_171),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1672),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1689),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1702),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1661),
.B(n_173),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1690),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1626),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1710),
.B(n_174),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1668),
.B(n_175),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1703),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1547),
.B(n_176),
.Y(n_1830)
);

AOI221x1_ASAP7_75t_L g1831 ( 
.A1(n_1571),
.A2(n_1602),
.B1(n_1613),
.B2(n_1585),
.C(n_1582),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1691),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1692),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1625),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1835)
);

NOR3xp33_ASAP7_75t_L g1836 ( 
.A(n_1568),
.B(n_179),
.C(n_180),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1705),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1704),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1574),
.B(n_180),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1718),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1686),
.B(n_181),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1615),
.B(n_182),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1729),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1577),
.B(n_183),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1699),
.B(n_184),
.Y(n_1845)
);

CKINVDCx12_ASAP7_75t_R g1846 ( 
.A(n_1557),
.Y(n_1846)
);

A2O1A1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1657),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1620),
.A2(n_190),
.B1(n_185),
.B2(n_188),
.Y(n_1848)
);

BUFx12f_ASAP7_75t_L g1849 ( 
.A(n_1590),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1554),
.B(n_188),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1569),
.B(n_190),
.Y(n_1851)
);

NOR2xp67_ASAP7_75t_L g1852 ( 
.A(n_1695),
.B(n_303),
.Y(n_1852)
);

AND3x1_ASAP7_75t_SL g1853 ( 
.A(n_1673),
.B(n_191),
.C(n_192),
.Y(n_1853)
);

AND3x1_ASAP7_75t_SL g1854 ( 
.A(n_1570),
.B(n_191),
.C(n_193),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1721),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1693),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1555),
.B(n_194),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1547),
.B(n_195),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1588),
.B(n_195),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1624),
.B(n_196),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1717),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1688),
.B(n_196),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1711),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1648),
.B(n_197),
.Y(n_1864)
);

BUFx2_ASAP7_75t_L g1865 ( 
.A(n_1669),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1650),
.B(n_198),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1678),
.B(n_198),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1578),
.B(n_199),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1607),
.B(n_199),
.Y(n_1869)
);

A2O1A1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1662),
.A2(n_1738),
.B(n_1675),
.C(n_1730),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1719),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1634),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1556),
.B(n_200),
.Y(n_1873)
);

AND3x1_ASAP7_75t_SL g1874 ( 
.A(n_1635),
.B(n_200),
.C(n_201),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1627),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1698),
.B(n_202),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1724),
.A2(n_1684),
.B1(n_1653),
.B2(n_1654),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1720),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1549),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1680),
.B(n_203),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1579),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1559),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1715),
.Y(n_1883)
);

BUFx8_ASAP7_75t_L g1884 ( 
.A(n_1551),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_1731),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1552),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1708),
.B(n_206),
.Y(n_1887)
);

AOI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1727),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1562),
.B(n_210),
.Y(n_1889)
);

BUFx8_ASAP7_75t_SL g1890 ( 
.A(n_1638),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1681),
.B(n_210),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1716),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1682),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_SL g1894 ( 
.A1(n_1685),
.A2(n_1701),
.B1(n_1663),
.B2(n_1722),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1565),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1640),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1707),
.A2(n_214),
.B1(n_211),
.B2(n_213),
.Y(n_1897)
);

INVxp67_ASAP7_75t_SL g1898 ( 
.A(n_1629),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1642),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1671),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1706),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1566),
.B(n_213),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1735),
.Y(n_1903)
);

AO21x2_ASAP7_75t_L g1904 ( 
.A1(n_1759),
.A2(n_1700),
.B(n_1736),
.Y(n_1904)
);

OAI21x1_ASAP7_75t_L g1905 ( 
.A1(n_1808),
.A2(n_1594),
.B(n_1589),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1787),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1745),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1749),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1741),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1744),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1774),
.Y(n_1911)
);

NOR2xp67_ASAP7_75t_SL g1912 ( 
.A(n_1849),
.B(n_1567),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1808),
.A2(n_1597),
.B(n_1595),
.Y(n_1913)
);

OR2x6_ASAP7_75t_L g1914 ( 
.A(n_1802),
.B(n_1658),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1744),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1740),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1761),
.B(n_1748),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1780),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1750),
.B(n_1598),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1749),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1766),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1775),
.Y(n_1922)
);

OA21x2_ASAP7_75t_L g1923 ( 
.A1(n_1784),
.A2(n_1603),
.B(n_1601),
.Y(n_1923)
);

OAI21x1_ASAP7_75t_L g1924 ( 
.A1(n_1830),
.A2(n_1605),
.B(n_1604),
.Y(n_1924)
);

OAI21x1_ASAP7_75t_L g1925 ( 
.A1(n_1830),
.A2(n_1606),
.B(n_1644),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1782),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1778),
.Y(n_1927)
);

CKINVDCx11_ASAP7_75t_R g1928 ( 
.A(n_1779),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1806),
.Y(n_1929)
);

OAI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1750),
.A2(n_1633),
.B(n_1630),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1792),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1807),
.Y(n_1932)
);

AO21x2_ASAP7_75t_L g1933 ( 
.A1(n_1784),
.A2(n_1646),
.B(n_1645),
.Y(n_1933)
);

OAI21x1_ASAP7_75t_L g1934 ( 
.A1(n_1858),
.A2(n_310),
.B(n_309),
.Y(n_1934)
);

OAI21x1_ASAP7_75t_L g1935 ( 
.A1(n_1858),
.A2(n_315),
.B(n_312),
.Y(n_1935)
);

BUFx12f_ASAP7_75t_L g1936 ( 
.A(n_1826),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1742),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1791),
.A2(n_214),
.B(n_215),
.Y(n_1938)
);

NAND2x1p5_ASAP7_75t_L g1939 ( 
.A(n_1768),
.B(n_316),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1768),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1742),
.Y(n_1941)
);

INVx6_ASAP7_75t_L g1942 ( 
.A(n_1768),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1751),
.B(n_318),
.Y(n_1943)
);

AO21x2_ASAP7_75t_L g1944 ( 
.A1(n_1805),
.A2(n_1781),
.B(n_1801),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1767),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1757),
.Y(n_1946)
);

OAI21x1_ASAP7_75t_SL g1947 ( 
.A1(n_1816),
.A2(n_215),
.B(n_216),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1801),
.A2(n_323),
.B(n_322),
.Y(n_1948)
);

INVx4_ASAP7_75t_L g1949 ( 
.A(n_1882),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_L g1950 ( 
.A1(n_1805),
.A2(n_327),
.B(n_324),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1783),
.B(n_217),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1794),
.Y(n_1952)
);

BUFx12f_ASAP7_75t_L g1953 ( 
.A(n_1872),
.Y(n_1953)
);

INVx5_ASAP7_75t_L g1954 ( 
.A(n_1778),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1811),
.B(n_218),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1809),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1816),
.A2(n_329),
.B(n_328),
.Y(n_1957)
);

NAND2x1p5_ASAP7_75t_L g1958 ( 
.A(n_1810),
.B(n_330),
.Y(n_1958)
);

BUFx2_ASAP7_75t_SL g1959 ( 
.A(n_1885),
.Y(n_1959)
);

OA21x2_ASAP7_75t_L g1960 ( 
.A1(n_1796),
.A2(n_333),
.B(n_332),
.Y(n_1960)
);

BUFx6f_ASAP7_75t_L g1961 ( 
.A(n_1755),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1895),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1798),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_SL g1964 ( 
.A1(n_1773),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1753),
.A2(n_335),
.B(n_334),
.Y(n_1965)
);

BUFx12f_ASAP7_75t_L g1966 ( 
.A(n_1884),
.Y(n_1966)
);

OAI21x1_ASAP7_75t_SL g1967 ( 
.A1(n_1756),
.A2(n_1795),
.B(n_1820),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1788),
.B(n_336),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1755),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1758),
.Y(n_1970)
);

NAND2x1p5_ASAP7_75t_L g1971 ( 
.A(n_1865),
.B(n_339),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1743),
.B(n_219),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1824),
.B(n_220),
.Y(n_1973)
);

BUFx2_ASAP7_75t_SL g1974 ( 
.A(n_1838),
.Y(n_1974)
);

OAI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1753),
.A2(n_341),
.B(n_340),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1804),
.Y(n_1976)
);

AO21x2_ASAP7_75t_L g1977 ( 
.A1(n_1746),
.A2(n_344),
.B(n_343),
.Y(n_1977)
);

INVx6_ASAP7_75t_L g1978 ( 
.A(n_1884),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1760),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1748),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1895),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1804),
.Y(n_1982)
);

CKINVDCx16_ASAP7_75t_R g1983 ( 
.A(n_1772),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1789),
.B(n_345),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1882),
.Y(n_1985)
);

BUFx12f_ASAP7_75t_L g1986 ( 
.A(n_1879),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1841),
.A2(n_223),
.B(n_224),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1747),
.Y(n_1988)
);

OAI21x1_ASAP7_75t_L g1989 ( 
.A1(n_1817),
.A2(n_348),
.B(n_347),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1762),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1882),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1813),
.Y(n_1992)
);

INVx6_ASAP7_75t_SL g1993 ( 
.A(n_1846),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1813),
.B(n_349),
.Y(n_1994)
);

BUFx3_ASAP7_75t_L g1995 ( 
.A(n_1813),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1786),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1817),
.Y(n_1997)
);

OAI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1883),
.A2(n_353),
.B(n_352),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1764),
.Y(n_1999)
);

OR2x6_ASAP7_75t_L g2000 ( 
.A(n_1763),
.B(n_354),
.Y(n_2000)
);

AO21x2_ASAP7_75t_L g2001 ( 
.A1(n_1770),
.A2(n_358),
.B(n_357),
.Y(n_2001)
);

BUFx8_ASAP7_75t_L g2002 ( 
.A(n_1754),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1777),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1771),
.Y(n_2004)
);

AO21x2_ASAP7_75t_L g2005 ( 
.A1(n_1799),
.A2(n_360),
.B(n_359),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1797),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1863),
.Y(n_2007)
);

BUFx12f_ASAP7_75t_L g2008 ( 
.A(n_1900),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1896),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1821),
.Y(n_2010)
);

BUFx8_ASAP7_75t_L g2011 ( 
.A(n_1966),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_SL g2012 ( 
.A1(n_1983),
.A2(n_1769),
.B1(n_1765),
.B2(n_1790),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1999),
.Y(n_2013)
);

INVx6_ASAP7_75t_L g2014 ( 
.A(n_1966),
.Y(n_2014)
);

CKINVDCx6p67_ASAP7_75t_R g2015 ( 
.A(n_1932),
.Y(n_2015)
);

AO22x1_ASAP7_75t_L g2016 ( 
.A1(n_2002),
.A2(n_1752),
.B1(n_1898),
.B2(n_1850),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1932),
.Y(n_2017)
);

BUFx10_ASAP7_75t_L g2018 ( 
.A(n_1978),
.Y(n_2018)
);

INVx6_ASAP7_75t_L g2019 ( 
.A(n_1978),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1911),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1999),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_2010),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2006),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1964),
.A2(n_1867),
.B1(n_1776),
.B2(n_1836),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1964),
.A2(n_1843),
.B1(n_1870),
.B2(n_1819),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1917),
.B(n_1820),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_2010),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1904),
.A2(n_1861),
.B1(n_1894),
.B2(n_1893),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1908),
.Y(n_2029)
);

INVx6_ASAP7_75t_L g2030 ( 
.A(n_1978),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2007),
.Y(n_2031)
);

OAI21xp5_ASAP7_75t_SL g2032 ( 
.A1(n_1987),
.A2(n_1831),
.B(n_1834),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_SL g2033 ( 
.A1(n_1960),
.A2(n_1967),
.B1(n_2001),
.B2(n_1977),
.Y(n_2033)
);

INVx6_ASAP7_75t_L g2034 ( 
.A(n_2002),
.Y(n_2034)
);

INVxp67_ASAP7_75t_L g2035 ( 
.A(n_2009),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_1904),
.A2(n_1897),
.B1(n_1800),
.B2(n_1815),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1929),
.Y(n_2037)
);

INVx8_ASAP7_75t_L g2038 ( 
.A(n_1929),
.Y(n_2038)
);

AOI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1919),
.A2(n_1793),
.B1(n_1875),
.B2(n_1827),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1906),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1918),
.B(n_1835),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1928),
.Y(n_2042)
);

BUFx8_ASAP7_75t_L g2043 ( 
.A(n_1936),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1937),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_SL g2045 ( 
.A1(n_1960),
.A2(n_1823),
.B1(n_1829),
.B2(n_1834),
.Y(n_2045)
);

OAI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_2000),
.A2(n_1848),
.B1(n_1823),
.B2(n_1829),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1908),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1941),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1928),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_1959),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_SL g2051 ( 
.A1(n_1960),
.A2(n_1860),
.B1(n_1862),
.B2(n_1864),
.Y(n_2051)
);

BUFx12f_ASAP7_75t_L g2052 ( 
.A(n_1936),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1909),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1920),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1920),
.Y(n_2055)
);

INVx6_ASAP7_75t_L g2056 ( 
.A(n_1911),
.Y(n_2056)
);

OAI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_2000),
.A2(n_1814),
.B1(n_1886),
.B2(n_1828),
.Y(n_2057)
);

CKINVDCx6p67_ASAP7_75t_R g2058 ( 
.A(n_1953),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_SL g2059 ( 
.A1(n_1977),
.A2(n_1866),
.B1(n_1876),
.B2(n_1844),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_1919),
.A2(n_1877),
.B1(n_1840),
.B2(n_1855),
.Y(n_2060)
);

INVx6_ASAP7_75t_L g2061 ( 
.A(n_2008),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1921),
.Y(n_2062)
);

BUFx4f_ASAP7_75t_SL g2063 ( 
.A(n_1993),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1988),
.Y(n_2064)
);

INVx6_ASAP7_75t_L g2065 ( 
.A(n_2008),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1990),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1918),
.A2(n_1847),
.B1(n_1851),
.B2(n_1881),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2003),
.Y(n_2068)
);

INVx6_ASAP7_75t_L g2069 ( 
.A(n_1953),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2023),
.Y(n_2070)
);

A2O1A1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_2032),
.A2(n_1987),
.B(n_1938),
.C(n_1852),
.Y(n_2071)
);

AO22x1_ASAP7_75t_L g2072 ( 
.A1(n_2043),
.A2(n_1962),
.B1(n_1981),
.B2(n_1917),
.Y(n_2072)
);

AOI222xp33_ASAP7_75t_L g2073 ( 
.A1(n_2025),
.A2(n_1868),
.B1(n_1973),
.B2(n_1842),
.C1(n_1859),
.C2(n_1857),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2046),
.A2(n_1845),
.B(n_1938),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2044),
.B(n_1980),
.Y(n_2075)
);

NAND2x1p5_ASAP7_75t_L g2076 ( 
.A(n_2020),
.B(n_1997),
.Y(n_2076)
);

OAI21x1_ASAP7_75t_SL g2077 ( 
.A1(n_2031),
.A2(n_1947),
.B(n_2053),
.Y(n_2077)
);

AOI21xp5_ASAP7_75t_L g2078 ( 
.A1(n_2045),
.A2(n_2057),
.B(n_2033),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2022),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_2056),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2013),
.Y(n_2081)
);

AO31x2_ASAP7_75t_L g2082 ( 
.A1(n_2027),
.A2(n_1931),
.A3(n_1952),
.B(n_2004),
.Y(n_2082)
);

INVx1_ASAP7_75t_SL g2083 ( 
.A(n_2040),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_2035),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2029),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2048),
.B(n_2026),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2021),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2064),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2040),
.B(n_1962),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_2056),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2067),
.A2(n_1930),
.B(n_1971),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_2066),
.B(n_1926),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_2015),
.B(n_1986),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_2059),
.A2(n_2001),
.B1(n_1996),
.B2(n_1944),
.Y(n_2094)
);

OAI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_2039),
.A2(n_2000),
.B1(n_1914),
.B2(n_1971),
.Y(n_2095)
);

INVxp67_ASAP7_75t_L g2096 ( 
.A(n_2041),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2068),
.B(n_1981),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2047),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2062),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2054),
.B(n_1944),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_L g2101 ( 
.A1(n_2016),
.A2(n_1930),
.B(n_2005),
.Y(n_2101)
);

AOI21xp33_ASAP7_75t_SL g2102 ( 
.A1(n_2038),
.A2(n_1922),
.B(n_1951),
.Y(n_2102)
);

AOI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_2036),
.A2(n_2005),
.B(n_1828),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2051),
.A2(n_2012),
.B1(n_2024),
.B2(n_2028),
.Y(n_2104)
);

OA21x2_ASAP7_75t_L g2105 ( 
.A1(n_2055),
.A2(n_1915),
.B(n_1910),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_2060),
.A2(n_1914),
.B(n_1997),
.Y(n_2106)
);

AOI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_2050),
.A2(n_1914),
.B(n_1957),
.Y(n_2107)
);

AOI21xp33_ASAP7_75t_SL g2108 ( 
.A1(n_2038),
.A2(n_1916),
.B(n_1955),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2082),
.Y(n_2109)
);

OAI221xp5_ASAP7_75t_SL g2110 ( 
.A1(n_2078),
.A2(n_1888),
.B1(n_1869),
.B2(n_1873),
.C(n_1880),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2104),
.A2(n_1869),
.B1(n_1901),
.B2(n_1880),
.C(n_1996),
.Y(n_2111)
);

INVxp67_ASAP7_75t_L g2112 ( 
.A(n_2084),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2081),
.Y(n_2113)
);

A2O1A1Ixp33_ASAP7_75t_L g2114 ( 
.A1(n_2091),
.A2(n_1912),
.B(n_1974),
.C(n_1972),
.Y(n_2114)
);

OAI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_2074),
.A2(n_2063),
.B1(n_2034),
.B2(n_2061),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2071),
.A2(n_2034),
.B1(n_2019),
.B2(n_2030),
.Y(n_2116)
);

OAI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2103),
.A2(n_2061),
.B1(n_2065),
.B2(n_1993),
.Y(n_2117)
);

A2O1A1Ixp33_ASAP7_75t_L g2118 ( 
.A1(n_2101),
.A2(n_1994),
.B(n_1995),
.C(n_1839),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2083),
.B(n_1963),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2083),
.B(n_2096),
.Y(n_2120)
);

BUFx4f_ASAP7_75t_SL g2121 ( 
.A(n_2080),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2087),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_SL g2123 ( 
.A1(n_2106),
.A2(n_1986),
.B1(n_2065),
.B2(n_1995),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2073),
.A2(n_1993),
.B1(n_1803),
.B2(n_1837),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2086),
.B(n_1963),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2073),
.A2(n_1903),
.B1(n_1818),
.B2(n_1825),
.Y(n_2126)
);

OAI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_2095),
.A2(n_2107),
.B1(n_2094),
.B2(n_2080),
.Y(n_2127)
);

OAI211xp5_ASAP7_75t_L g2128 ( 
.A1(n_2108),
.A2(n_2102),
.B(n_2089),
.C(n_2088),
.Y(n_2128)
);

AOI222xp33_ASAP7_75t_L g2129 ( 
.A1(n_2072),
.A2(n_2086),
.B1(n_1822),
.B2(n_1832),
.C1(n_1833),
.C2(n_1856),
.Y(n_2129)
);

BUFx3_ASAP7_75t_L g2130 ( 
.A(n_2093),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2082),
.Y(n_2131)
);

AOI221xp5_ASAP7_75t_L g2132 ( 
.A1(n_2099),
.A2(n_1946),
.B1(n_1979),
.B2(n_1970),
.C(n_1945),
.Y(n_2132)
);

AO21x2_ASAP7_75t_L g2133 ( 
.A1(n_2109),
.A2(n_2100),
.B(n_2077),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_2121),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_2121),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2112),
.B(n_2129),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2113),
.B(n_2097),
.Y(n_2137)
);

NOR2x1_ASAP7_75t_L g2138 ( 
.A(n_2130),
.B(n_2037),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2131),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2122),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2125),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2140),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2137),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_2134),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2136),
.A2(n_2115),
.B(n_2127),
.Y(n_2145)
);

INVx4_ASAP7_75t_L g2146 ( 
.A(n_2134),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2138),
.A2(n_2124),
.B1(n_2126),
.B2(n_2114),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_2146),
.B(n_2135),
.Y(n_2148)
);

OAI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2147),
.A2(n_2117),
.B1(n_2111),
.B2(n_2141),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2142),
.Y(n_2150)
);

HB1xp67_ASAP7_75t_L g2151 ( 
.A(n_2144),
.Y(n_2151)
);

AOI221xp5_ASAP7_75t_L g2152 ( 
.A1(n_2145),
.A2(n_2110),
.B1(n_2126),
.B2(n_2124),
.C(n_2117),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2143),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2146),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_2147),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2144),
.B(n_2135),
.Y(n_2156)
);

OAI31xp33_ASAP7_75t_SL g2157 ( 
.A1(n_2147),
.A2(n_2115),
.A3(n_2128),
.B(n_2116),
.Y(n_2157)
);

NOR4xp25_ASAP7_75t_SL g2158 ( 
.A(n_2155),
.B(n_2042),
.C(n_2049),
.D(n_2011),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2155),
.B(n_2141),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2150),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2151),
.B(n_2133),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2156),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2153),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2154),
.B(n_2092),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_2157),
.B(n_2123),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2155),
.B(n_2133),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2148),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2157),
.B(n_2058),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2158),
.B(n_2120),
.Y(n_2169)
);

XOR2x2_ASAP7_75t_L g2170 ( 
.A(n_2165),
.B(n_2152),
.Y(n_2170)
);

AND2x4_ASAP7_75t_L g2171 ( 
.A(n_2162),
.B(n_2167),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2158),
.B(n_2017),
.Y(n_2172)
);

NOR4xp25_ASAP7_75t_L g2173 ( 
.A(n_2163),
.B(n_2149),
.C(n_1889),
.D(n_1902),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_2168),
.B(n_2160),
.Y(n_2174)
);

XOR2x2_ASAP7_75t_L g2175 ( 
.A(n_2159),
.B(n_2166),
.Y(n_2175)
);

OAI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2159),
.A2(n_2118),
.B(n_2119),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2171),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2171),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2169),
.B(n_2164),
.Y(n_2179)
);

OAI21xp33_ASAP7_75t_SL g2180 ( 
.A1(n_2173),
.A2(n_2161),
.B(n_2043),
.Y(n_2180)
);

OAI21xp33_ASAP7_75t_L g2181 ( 
.A1(n_2179),
.A2(n_2173),
.B(n_2174),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2178),
.Y(n_2182)
);

AOI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2180),
.A2(n_2170),
.B1(n_2175),
.B2(n_2174),
.Y(n_2183)
);

INVxp67_ASAP7_75t_L g2184 ( 
.A(n_2177),
.Y(n_2184)
);

NAND2x1_ASAP7_75t_L g2185 ( 
.A(n_2182),
.B(n_2172),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2184),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2181),
.B(n_2180),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2183),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2182),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_L g2190 ( 
.A1(n_2188),
.A2(n_2176),
.B1(n_2139),
.B2(n_2133),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2187),
.B(n_2069),
.Y(n_2191)
);

OAI21xp5_ASAP7_75t_SL g2192 ( 
.A1(n_2189),
.A2(n_2011),
.B(n_2017),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2186),
.Y(n_2193)
);

OAI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_2185),
.A2(n_1887),
.B(n_1891),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2187),
.B(n_2069),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2187),
.A2(n_2052),
.B1(n_2014),
.B2(n_2030),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2187),
.B(n_2014),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2186),
.Y(n_2198)
);

NAND3xp33_ASAP7_75t_SL g2199 ( 
.A(n_2185),
.B(n_1939),
.C(n_2090),
.Y(n_2199)
);

AO22x2_ASAP7_75t_L g2200 ( 
.A1(n_2193),
.A2(n_2139),
.B1(n_1994),
.B2(n_1943),
.Y(n_2200)
);

AOI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_2192),
.A2(n_2020),
.B(n_2070),
.Y(n_2201)
);

AOI211x1_ASAP7_75t_SL g2202 ( 
.A1(n_2199),
.A2(n_1874),
.B(n_2075),
.C(n_1853),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2198),
.B(n_2019),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2197),
.B(n_2191),
.Y(n_2204)
);

AOI221x1_ASAP7_75t_L g2205 ( 
.A1(n_2195),
.A2(n_1899),
.B1(n_2075),
.B2(n_1878),
.C(n_1871),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2194),
.B(n_2018),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2190),
.B(n_2132),
.Y(n_2207)
);

AOI21xp5_ASAP7_75t_L g2208 ( 
.A1(n_2192),
.A2(n_1989),
.B(n_1943),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2196),
.B(n_1890),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2193),
.B(n_224),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_2196),
.B(n_2076),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2192),
.A2(n_225),
.B(n_226),
.Y(n_2212)
);

INVxp67_ASAP7_75t_L g2213 ( 
.A(n_2204),
.Y(n_2213)
);

OAI21xp33_ASAP7_75t_SL g2214 ( 
.A1(n_2206),
.A2(n_1924),
.B(n_1925),
.Y(n_2214)
);

NOR2xp67_ASAP7_75t_L g2215 ( 
.A(n_2212),
.B(n_225),
.Y(n_2215)
);

NAND4xp25_ASAP7_75t_L g2216 ( 
.A(n_2203),
.B(n_1812),
.C(n_229),
.D(n_226),
.Y(n_2216)
);

OAI221xp5_ASAP7_75t_L g2217 ( 
.A1(n_2210),
.A2(n_1739),
.B1(n_2076),
.B2(n_1892),
.C(n_1939),
.Y(n_2217)
);

AOI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2207),
.A2(n_1854),
.B1(n_2100),
.B2(n_1907),
.C(n_1968),
.Y(n_2218)
);

AOI21xp33_ASAP7_75t_L g2219 ( 
.A1(n_2209),
.A2(n_227),
.B(n_229),
.Y(n_2219)
);

AOI21xp33_ASAP7_75t_L g2220 ( 
.A1(n_2200),
.A2(n_227),
.B(n_230),
.Y(n_2220)
);

OAI211xp5_ASAP7_75t_SL g2221 ( 
.A1(n_2211),
.A2(n_233),
.B(n_230),
.C(n_232),
.Y(n_2221)
);

NOR2x1_ASAP7_75t_L g2222 ( 
.A(n_2201),
.B(n_232),
.Y(n_2222)
);

AOI221xp5_ASAP7_75t_SL g2223 ( 
.A1(n_2208),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.C(n_236),
.Y(n_2223)
);

OAI21xp33_ASAP7_75t_SL g2224 ( 
.A1(n_2202),
.A2(n_1949),
.B(n_1913),
.Y(n_2224)
);

AOI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_2205),
.A2(n_234),
.B(n_235),
.Y(n_2225)
);

AOI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_2215),
.A2(n_2200),
.B1(n_1933),
.B2(n_1923),
.Y(n_2226)
);

O2A1O1Ixp33_ASAP7_75t_L g2227 ( 
.A1(n_2213),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_2227)
);

OAI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2222),
.A2(n_1949),
.B1(n_1991),
.B2(n_1985),
.Y(n_2228)
);

AO22x1_ASAP7_75t_L g2229 ( 
.A1(n_2223),
.A2(n_240),
.B1(n_237),
.B2(n_239),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2225),
.Y(n_2230)
);

INVxp67_ASAP7_75t_L g2231 ( 
.A(n_2220),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2217),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2221),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2218),
.A2(n_2219),
.B1(n_2224),
.B2(n_2214),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2216),
.Y(n_2235)
);

AOI22xp33_ASAP7_75t_SL g2236 ( 
.A1(n_2213),
.A2(n_1923),
.B1(n_1992),
.B2(n_1991),
.Y(n_2236)
);

AOI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2220),
.A2(n_1968),
.B1(n_1984),
.B2(n_1985),
.C(n_1785),
.Y(n_2237)
);

OAI211xp5_ASAP7_75t_SL g2238 ( 
.A1(n_2230),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_2231),
.B(n_242),
.Y(n_2239)
);

AOI211xp5_ASAP7_75t_L g2240 ( 
.A1(n_2229),
.A2(n_1957),
.B(n_1998),
.C(n_1935),
.Y(n_2240)
);

AOI221xp5_ASAP7_75t_L g2241 ( 
.A1(n_2234),
.A2(n_1984),
.B1(n_244),
.B2(n_245),
.C(n_246),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2233),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_2232),
.A2(n_1992),
.B1(n_1933),
.B2(n_2105),
.Y(n_2243)
);

AOI321xp33_ASAP7_75t_L g2244 ( 
.A1(n_2235),
.A2(n_243),
.A3(n_244),
.B1(n_245),
.B2(n_248),
.C(n_249),
.Y(n_2244)
);

AOI211xp5_ASAP7_75t_L g2245 ( 
.A1(n_2227),
.A2(n_1934),
.B(n_1948),
.C(n_250),
.Y(n_2245)
);

OAI211xp5_ASAP7_75t_L g2246 ( 
.A1(n_2226),
.A2(n_250),
.B(n_243),
.C(n_248),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2237),
.A2(n_1923),
.B1(n_1992),
.B2(n_2105),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2228),
.B(n_251),
.Y(n_2248)
);

O2A1O1Ixp33_ASAP7_75t_L g2249 ( 
.A1(n_2236),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_2249)
);

OAI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_2230),
.A2(n_1992),
.B1(n_1958),
.B2(n_1961),
.Y(n_2250)
);

O2A1O1Ixp33_ASAP7_75t_L g2251 ( 
.A1(n_2230),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_2251)
);

O2A1O1Ixp33_ASAP7_75t_L g2252 ( 
.A1(n_2230),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_2252)
);

AOI222xp33_ASAP7_75t_L g2253 ( 
.A1(n_2231),
.A2(n_1950),
.B1(n_1965),
.B2(n_1975),
.C1(n_259),
.C2(n_260),
.Y(n_2253)
);

O2A1O1Ixp33_ASAP7_75t_L g2254 ( 
.A1(n_2251),
.A2(n_258),
.B(n_255),
.C(n_257),
.Y(n_2254)
);

NAND3xp33_ASAP7_75t_L g2255 ( 
.A(n_2239),
.B(n_258),
.C(n_259),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2244),
.Y(n_2256)
);

OAI211xp5_ASAP7_75t_SL g2257 ( 
.A1(n_2242),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_2257)
);

AOI211xp5_ASAP7_75t_L g2258 ( 
.A1(n_2238),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_2258)
);

AOI222xp33_ASAP7_75t_L g2259 ( 
.A1(n_2246),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.C1(n_267),
.C2(n_268),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2252),
.A2(n_265),
.B(n_266),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2241),
.A2(n_1905),
.B1(n_1958),
.B2(n_1942),
.Y(n_2261)
);

INVx2_ASAP7_75t_SL g2262 ( 
.A(n_2248),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2247),
.Y(n_2263)
);

AOI221xp5_ASAP7_75t_L g2264 ( 
.A1(n_2249),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.C(n_272),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2245),
.Y(n_2265)
);

INVx1_ASAP7_75t_SL g2266 ( 
.A(n_2250),
.Y(n_2266)
);

XNOR2xp5_ASAP7_75t_L g2267 ( 
.A(n_2240),
.B(n_270),
.Y(n_2267)
);

NAND3xp33_ASAP7_75t_L g2268 ( 
.A(n_2243),
.B(n_271),
.C(n_273),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2253),
.B(n_274),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2244),
.Y(n_2270)
);

AOI211x1_ASAP7_75t_L g2271 ( 
.A1(n_2246),
.A2(n_274),
.B(n_275),
.C(n_276),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_2242),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_2242),
.Y(n_2273)
);

AOI221xp5_ASAP7_75t_L g2274 ( 
.A1(n_2249),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.C(n_278),
.Y(n_2274)
);

NOR3xp33_ASAP7_75t_L g2275 ( 
.A(n_2242),
.B(n_277),
.C(n_279),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2242),
.Y(n_2276)
);

NAND3xp33_ASAP7_75t_L g2277 ( 
.A(n_2239),
.B(n_279),
.C(n_280),
.Y(n_2277)
);

AOI221xp5_ASAP7_75t_L g2278 ( 
.A1(n_2249),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.C(n_283),
.Y(n_2278)
);

NOR2x1_ASAP7_75t_L g2279 ( 
.A(n_2272),
.B(n_2276),
.Y(n_2279)
);

AOI321xp33_ASAP7_75t_L g2280 ( 
.A1(n_2256),
.A2(n_281),
.A3(n_282),
.B1(n_283),
.B2(n_284),
.C(n_285),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2270),
.Y(n_2281)
);

OAI32xp33_ASAP7_75t_L g2282 ( 
.A1(n_2269),
.A2(n_284),
.A3(n_286),
.B1(n_287),
.B2(n_1927),
.Y(n_2282)
);

OAI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_2273),
.A2(n_1961),
.B1(n_1982),
.B2(n_1976),
.Y(n_2283)
);

BUFx3_ASAP7_75t_L g2284 ( 
.A(n_2262),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2271),
.Y(n_2285)
);

INVxp67_ASAP7_75t_SL g2286 ( 
.A(n_2275),
.Y(n_2286)
);

OR2x2_ASAP7_75t_L g2287 ( 
.A(n_2255),
.B(n_286),
.Y(n_2287)
);

O2A1O1Ixp33_ASAP7_75t_L g2288 ( 
.A1(n_2265),
.A2(n_1969),
.B(n_362),
.C(n_363),
.Y(n_2288)
);

AND3x2_ASAP7_75t_L g2289 ( 
.A(n_2258),
.B(n_361),
.C(n_364),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2259),
.B(n_2082),
.Y(n_2290)
);

OAI211xp5_ASAP7_75t_L g2291 ( 
.A1(n_2264),
.A2(n_366),
.B(n_367),
.C(n_368),
.Y(n_2291)
);

OA22x2_ASAP7_75t_L g2292 ( 
.A1(n_2267),
.A2(n_1927),
.B1(n_1969),
.B2(n_2098),
.Y(n_2292)
);

AOI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2274),
.A2(n_1942),
.B1(n_1961),
.B2(n_2085),
.Y(n_2293)
);

AOI222xp33_ASAP7_75t_L g2294 ( 
.A1(n_2266),
.A2(n_1961),
.B1(n_2079),
.B2(n_1976),
.C1(n_1982),
.C2(n_1942),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2277),
.B(n_370),
.Y(n_2295)
);

NAND4xp75_ASAP7_75t_L g2296 ( 
.A(n_2260),
.B(n_373),
.C(n_374),
.D(n_375),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2263),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_2284),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2285),
.B(n_2257),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2289),
.B(n_2278),
.Y(n_2300)
);

AND3x4_ASAP7_75t_L g2301 ( 
.A(n_2279),
.B(n_2254),
.C(n_2268),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2281),
.B(n_2261),
.Y(n_2302)
);

OAI221xp5_ASAP7_75t_L g2303 ( 
.A1(n_2280),
.A2(n_2286),
.B1(n_2287),
.B2(n_2291),
.C(n_2297),
.Y(n_2303)
);

OAI211xp5_ASAP7_75t_SL g2304 ( 
.A1(n_2295),
.A2(n_2290),
.B(n_2288),
.C(n_2294),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2282),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2296),
.B(n_2292),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2293),
.Y(n_2307)
);

NOR2x1_ASAP7_75t_L g2308 ( 
.A(n_2283),
.B(n_379),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2285),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_2285),
.B(n_381),
.Y(n_2310)
);

NOR4xp25_ASAP7_75t_L g2311 ( 
.A(n_2286),
.B(n_383),
.C(n_384),
.D(n_386),
.Y(n_2311)
);

OAI221xp5_ASAP7_75t_L g2312 ( 
.A1(n_2279),
.A2(n_1982),
.B1(n_1976),
.B2(n_1940),
.C(n_1954),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2284),
.Y(n_2313)
);

HB1xp67_ASAP7_75t_L g2314 ( 
.A(n_2285),
.Y(n_2314)
);

OAI221xp5_ASAP7_75t_SL g2315 ( 
.A1(n_2281),
.A2(n_1952),
.B1(n_1931),
.B2(n_390),
.C(n_392),
.Y(n_2315)
);

XOR2xp5_ASAP7_75t_L g2316 ( 
.A(n_2281),
.B(n_388),
.Y(n_2316)
);

CKINVDCx16_ASAP7_75t_R g2317 ( 
.A(n_2284),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2317),
.Y(n_2318)
);

AND2x4_ASAP7_75t_L g2319 ( 
.A(n_2298),
.B(n_1976),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2314),
.Y(n_2320)
);

NOR4xp25_ASAP7_75t_L g2321 ( 
.A(n_2309),
.B(n_389),
.C(n_393),
.D(n_396),
.Y(n_2321)
);

NAND4xp25_ASAP7_75t_L g2322 ( 
.A(n_2299),
.B(n_397),
.C(n_398),
.D(n_399),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2313),
.B(n_1982),
.Y(n_2323)
);

AOI211xp5_ASAP7_75t_L g2324 ( 
.A1(n_2303),
.A2(n_402),
.B(n_403),
.C(n_404),
.Y(n_2324)
);

AOI211xp5_ASAP7_75t_L g2325 ( 
.A1(n_2302),
.A2(n_405),
.B(n_406),
.C(n_407),
.Y(n_2325)
);

NOR2x1p5_ASAP7_75t_L g2326 ( 
.A(n_2305),
.B(n_1940),
.Y(n_2326)
);

NAND4xp25_ASAP7_75t_L g2327 ( 
.A(n_2310),
.B(n_408),
.C(n_409),
.D(n_410),
.Y(n_2327)
);

OAI21xp33_ASAP7_75t_SL g2328 ( 
.A1(n_2300),
.A2(n_411),
.B(n_413),
.Y(n_2328)
);

AOI22x1_ASAP7_75t_SL g2329 ( 
.A1(n_2307),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_2329)
);

NOR4xp25_ASAP7_75t_L g2330 ( 
.A(n_2304),
.B(n_417),
.C(n_419),
.D(n_420),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2301),
.A2(n_1954),
.B1(n_1940),
.B2(n_1956),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2316),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2311),
.B(n_421),
.Y(n_2333)
);

XNOR2xp5_ASAP7_75t_L g2334 ( 
.A(n_2318),
.B(n_2302),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2320),
.Y(n_2335)
);

OR3x2_ASAP7_75t_L g2336 ( 
.A(n_2332),
.B(n_2333),
.C(n_2327),
.Y(n_2336)
);

NOR2x1_ASAP7_75t_L g2337 ( 
.A(n_2326),
.B(n_2306),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2319),
.B(n_2308),
.Y(n_2338)
);

AND3x4_ASAP7_75t_L g2339 ( 
.A(n_2330),
.B(n_2315),
.C(n_2312),
.Y(n_2339)
);

NOR3xp33_ASAP7_75t_L g2340 ( 
.A(n_2328),
.B(n_422),
.C(n_425),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2329),
.Y(n_2341)
);

OR3x1_ASAP7_75t_L g2342 ( 
.A(n_2322),
.B(n_426),
.C(n_427),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2323),
.Y(n_2343)
);

NAND2x1p5_ASAP7_75t_L g2344 ( 
.A(n_2324),
.B(n_1940),
.Y(n_2344)
);

AND4x1_ASAP7_75t_L g2345 ( 
.A(n_2325),
.B(n_428),
.C(n_429),
.D(n_433),
.Y(n_2345)
);

OR2x6_ASAP7_75t_L g2346 ( 
.A(n_2331),
.B(n_436),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2321),
.Y(n_2347)
);

INVxp67_ASAP7_75t_SL g2348 ( 
.A(n_2318),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2318),
.Y(n_2349)
);

AOI22xp5_ASAP7_75t_L g2350 ( 
.A1(n_2348),
.A2(n_1954),
.B1(n_441),
.B2(n_442),
.Y(n_2350)
);

OAI22x1_ASAP7_75t_L g2351 ( 
.A1(n_2334),
.A2(n_1954),
.B1(n_443),
.B2(n_445),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2349),
.A2(n_439),
.B1(n_447),
.B2(n_453),
.Y(n_2352)
);

XNOR2xp5_ASAP7_75t_L g2353 ( 
.A(n_2342),
.B(n_2337),
.Y(n_2353)
);

OAI22x1_ASAP7_75t_L g2354 ( 
.A1(n_2347),
.A2(n_454),
.B1(n_456),
.B2(n_459),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2341),
.Y(n_2355)
);

HB1xp67_ASAP7_75t_L g2356 ( 
.A(n_2335),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_2338),
.B(n_460),
.Y(n_2357)
);

INVxp67_ASAP7_75t_SL g2358 ( 
.A(n_2343),
.Y(n_2358)
);

AOI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2339),
.A2(n_461),
.B1(n_463),
.B2(n_464),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2356),
.Y(n_2360)
);

INVx2_ASAP7_75t_SL g2361 ( 
.A(n_2353),
.Y(n_2361)
);

AOI22xp33_ASAP7_75t_SL g2362 ( 
.A1(n_2358),
.A2(n_2355),
.B1(n_2346),
.B2(n_2344),
.Y(n_2362)
);

AOI22xp33_ASAP7_75t_L g2363 ( 
.A1(n_2351),
.A2(n_2336),
.B1(n_2340),
.B2(n_2346),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2357),
.Y(n_2364)
);

INVxp67_ASAP7_75t_L g2365 ( 
.A(n_2354),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2359),
.Y(n_2366)
);

AOI22xp33_ASAP7_75t_L g2367 ( 
.A1(n_2360),
.A2(n_2350),
.B1(n_2352),
.B2(n_2345),
.Y(n_2367)
);

AOI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2361),
.A2(n_465),
.B1(n_467),
.B2(n_469),
.Y(n_2368)
);

OAI22xp33_ASAP7_75t_SL g2369 ( 
.A1(n_2364),
.A2(n_470),
.B1(n_471),
.B2(n_473),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_L g2370 ( 
.A1(n_2365),
.A2(n_474),
.B1(n_475),
.B2(n_476),
.Y(n_2370)
);

AOI31xp33_ASAP7_75t_L g2371 ( 
.A1(n_2367),
.A2(n_2362),
.A3(n_2363),
.B(n_2366),
.Y(n_2371)
);

AOI22xp33_ASAP7_75t_L g2372 ( 
.A1(n_2368),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_2372)
);

AOI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_2369),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2371),
.A2(n_2370),
.B1(n_485),
.B2(n_486),
.Y(n_2374)
);

AOI22x1_ASAP7_75t_L g2375 ( 
.A1(n_2373),
.A2(n_483),
.B1(n_487),
.B2(n_488),
.Y(n_2375)
);

INVxp33_ASAP7_75t_L g2376 ( 
.A(n_2374),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2376),
.Y(n_2377)
);

XOR2xp5_ASAP7_75t_L g2378 ( 
.A(n_2377),
.B(n_2375),
.Y(n_2378)
);

OAI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2378),
.A2(n_2372),
.B(n_491),
.Y(n_2379)
);

OR2x6_ASAP7_75t_L g2380 ( 
.A(n_2378),
.B(n_490),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2379),
.A2(n_492),
.B(n_494),
.Y(n_2381)
);

OAI22xp33_ASAP7_75t_L g2382 ( 
.A1(n_2381),
.A2(n_2380),
.B1(n_495),
.B2(n_497),
.Y(n_2382)
);


endmodule