module fake_jpeg_2821_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_20),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_1),
.B(n_4),
.C(n_16),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_23),
.C(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_16),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_25),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_28),
.B1(n_22),
.B2(n_27),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_29),
.CI(n_31),
.CON(n_38),
.SN(n_38)
);

AOI221xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_33),
.B2(n_7),
.C(n_10),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_40),
.C(n_38),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_10),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_44),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_46),
.B(n_4),
.Y(n_47)
);


endmodule