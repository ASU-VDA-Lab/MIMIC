module fake_jpeg_2793_n_421 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_46),
.Y(n_125)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_49),
.Y(n_120)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_18),
.B(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_64),
.Y(n_97)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_1),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_72),
.Y(n_94)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_67),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_18),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_25),
.B(n_1),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_71),
.B(n_3),
.Y(n_126)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_2),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_74),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_31),
.B(n_3),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_80),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_21),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_35),
.B1(n_28),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_84),
.A2(n_114),
.B1(n_117),
.B2(n_12),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_35),
.B1(n_21),
.B2(n_42),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_89),
.A2(n_12),
.B1(n_14),
.B2(n_120),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_49),
.Y(n_146)
);

AND2x4_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_21),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_107),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_108),
.B(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_27),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_35),
.B1(n_39),
.B2(n_32),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_110),
.A2(n_113),
.B1(n_129),
.B2(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_39),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_124),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_60),
.A2(n_39),
.B1(n_32),
.B2(n_42),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_55),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_25),
.B(n_33),
.C(n_32),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_36),
.B(n_38),
.C(n_7),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_23),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_23),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_6),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_62),
.A2(n_66),
.B1(n_58),
.B2(n_78),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_49),
.B1(n_30),
.B2(n_36),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_59),
.A2(n_33),
.B1(n_36),
.B2(n_30),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_3),
.Y(n_135)
);

NAND2x1_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_10),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_43),
.B(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_36),
.B1(n_30),
.B2(n_38),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_81),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_138),
.B(n_160),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_139),
.Y(n_223)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_141),
.B(n_149),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_76),
.B1(n_75),
.B2(n_74),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_142),
.A2(n_145),
.B1(n_152),
.B2(n_140),
.Y(n_235)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_36),
.C(n_30),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_179),
.C(n_123),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_5),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_94),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_46),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_150),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_92),
.B1(n_132),
.B2(n_116),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_155),
.B(n_173),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_5),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_6),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_161),
.A2(n_167),
.B1(n_181),
.B2(n_86),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_14),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_162),
.B(n_158),
.Y(n_234)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_164),
.B(n_99),
.Y(n_217)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_118),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_123),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_84),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

BUFx8_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_183),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_8),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_175),
.A2(n_190),
.B1(n_132),
.B2(n_130),
.Y(n_194)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_176),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_101),
.B1(n_87),
.B2(n_122),
.Y(n_214)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_98),
.B(n_96),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_180),
.B(n_95),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_89),
.A2(n_12),
.B1(n_14),
.B2(n_107),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_187),
.B1(n_85),
.B2(n_90),
.Y(n_193)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_185),
.B(n_95),
.Y(n_232)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_112),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_107),
.A2(n_12),
.B1(n_115),
.B2(n_116),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_189),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_98),
.A2(n_85),
.B1(n_96),
.B2(n_90),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_193),
.A2(n_196),
.B1(n_216),
.B2(n_224),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_199),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_156),
.B1(n_174),
.B2(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_178),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_214),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_212),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_150),
.B(n_87),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_130),
.B1(n_86),
.B2(n_127),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_213),
.A2(n_235),
.B1(n_187),
.B2(n_146),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_217),
.B(n_232),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_150),
.B(n_153),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_225),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_146),
.B(n_173),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_157),
.A2(n_101),
.B1(n_119),
.B2(n_99),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_119),
.B1(n_122),
.B2(n_134),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_155),
.B(n_95),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_155),
.B(n_95),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_168),
.B(n_154),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_179),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_233),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_238),
.B(n_257),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_241),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

INVx6_ASAP7_75t_SL g302 ( 
.A(n_242),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_197),
.B(n_173),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_259),
.Y(n_279)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_151),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_253),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_228),
.C(n_200),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_268),
.C(n_271),
.Y(n_281)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_254),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_170),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_179),
.B(n_167),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_191),
.B(n_210),
.Y(n_297)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_207),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_196),
.A2(n_161),
.B(n_159),
.C(n_144),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_229),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_266),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_197),
.B(n_165),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_260),
.B(n_261),
.Y(n_298)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_252),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_205),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_183),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_171),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_270),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_186),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_188),
.C(n_189),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_208),
.B(n_139),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_221),
.C(n_226),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_198),
.B(n_143),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_274),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_209),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_193),
.B1(n_225),
.B2(n_232),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_277),
.B1(n_292),
.B2(n_295),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_248),
.B1(n_254),
.B2(n_243),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

CKINVDCx12_ASAP7_75t_R g287 ( 
.A(n_258),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_232),
.B1(n_206),
.B2(n_195),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_240),
.B(n_212),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_293),
.B(n_261),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_281),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_267),
.A2(n_224),
.B1(n_216),
.B2(n_231),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_243),
.A2(n_191),
.B1(n_192),
.B2(n_215),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_297),
.A2(n_241),
.B(n_262),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_236),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_259),
.B(n_191),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_305),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_192),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_255),
.A2(n_211),
.B1(n_223),
.B2(n_219),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_306),
.A2(n_264),
.B1(n_227),
.B2(n_219),
.Y(n_329)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_277),
.A2(n_239),
.B1(n_257),
.B2(n_263),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_309),
.A2(n_323),
.B1(n_324),
.B2(n_327),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_313),
.C(n_315),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_238),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_319),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_272),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_293),
.C(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_239),
.C(n_268),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_328),
.C(n_330),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_240),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_244),
.Y(n_320)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_320),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_321),
.A2(n_331),
.B(n_287),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_263),
.B1(n_262),
.B2(n_251),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_289),
.A2(n_263),
.B1(n_271),
.B2(n_250),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_326),
.B(n_280),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_256),
.B1(n_245),
.B2(n_249),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_265),
.C(n_227),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_329),
.A2(n_333),
.B1(n_290),
.B2(n_291),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_209),
.Y(n_330)
);

OAI32xp33_ASAP7_75t_L g331 ( 
.A1(n_279),
.A2(n_169),
.A3(n_176),
.B1(n_264),
.B2(n_303),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_288),
.Y(n_332)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_295),
.A2(n_278),
.B1(n_296),
.B2(n_306),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_288),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_334),
.B(n_282),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_283),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_337),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_278),
.Y(n_337)
);

FAx1_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_301),
.CI(n_297),
.CON(n_338),
.SN(n_338)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_342),
.Y(n_361)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_349),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_340),
.A2(n_347),
.B1(n_355),
.B2(n_331),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_311),
.A2(n_300),
.B(n_285),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_352),
.B(n_314),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_301),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_356),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_317),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_322),
.A2(n_282),
.B1(n_280),
.B2(n_275),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_326),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_319),
.B(n_307),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_307),
.B(n_275),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_333),
.A2(n_304),
.B1(n_325),
.B2(n_309),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_304),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_348),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_328),
.C(n_311),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_362),
.C(n_364),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_355),
.A2(n_323),
.B1(n_324),
.B2(n_332),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_360),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_351),
.B(n_321),
.C(n_330),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_352),
.B(n_338),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_314),
.C(n_320),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_317),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_367),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_327),
.C(n_329),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_354),
.C(n_356),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_337),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_341),
.Y(n_384)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_374),
.Y(n_387)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_378),
.Y(n_393)
);

XNOR2x1_ASAP7_75t_SL g378 ( 
.A(n_361),
.B(n_338),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_383),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_382),
.B(n_359),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_367),
.A2(n_340),
.B1(n_342),
.B2(n_347),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_390),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_341),
.C(n_304),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_392),
.A2(n_376),
.B(n_370),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_388),
.A2(n_361),
.B1(n_360),
.B2(n_375),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_394),
.Y(n_401)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_395),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_386),
.A2(n_361),
.B1(n_369),
.B2(n_358),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_399),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_368),
.C(n_362),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_398),
.A2(n_376),
.B(n_359),
.Y(n_402)
);

BUFx24_ASAP7_75t_SL g399 ( 
.A(n_381),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_400),
.A2(n_379),
.B1(n_387),
.B2(n_364),
.Y(n_405)
);

NAND3xp33_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_393),
.C(n_400),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_391),
.A2(n_387),
.B1(n_389),
.B2(n_380),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_403),
.A2(n_383),
.B1(n_378),
.B2(n_384),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_405),
.B(n_394),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_407),
.B(n_393),
.C(n_390),
.Y(n_410)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_404),
.A2(n_397),
.B(n_398),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_410),
.C(n_412),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_411),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_414),
.A2(n_406),
.B(n_401),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_416),
.A2(n_417),
.B(n_413),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_415),
.B(n_401),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_377),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_419),
.A2(n_357),
.B(n_304),
.Y(n_420)
);

BUFx24_ASAP7_75t_SL g421 ( 
.A(n_420),
.Y(n_421)
);


endmodule