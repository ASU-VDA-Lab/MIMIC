module fake_jpeg_14791_n_192 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_20),
.B1(n_16),
.B2(n_25),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_49),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_28),
.B1(n_24),
.B2(n_41),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_54),
.B1(n_53),
.B2(n_46),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_28),
.B1(n_33),
.B2(n_41),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_69),
.B1(n_45),
.B2(n_27),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_55),
.Y(n_92)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_58),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_15),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_38),
.B1(n_27),
.B2(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_92),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_87),
.B1(n_96),
.B2(n_100),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_90),
.C(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_21),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_46),
.B(n_55),
.C(n_43),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_51),
.B1(n_52),
.B2(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_51),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_16),
.B1(n_23),
.B2(n_38),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_37),
.C(n_32),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_35),
.C(n_32),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_31),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_110),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_66),
.B1(n_77),
.B2(n_74),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_119),
.B1(n_97),
.B2(n_89),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_51),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_71),
.B1(n_76),
.B2(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_89),
.B(n_88),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_101),
.C(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_128),
.C(n_129),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_90),
.B(n_118),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_111),
.B(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_84),
.C(n_90),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_96),
.C(n_82),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_116),
.C(n_119),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_30),
.B(n_3),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_110),
.B(n_118),
.C(n_104),
.D(n_120),
.Y(n_138)
);

AOI321xp33_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_144),
.A3(n_151),
.B1(n_134),
.B2(n_22),
.C(n_31),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_35),
.C(n_31),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_103),
.B1(n_104),
.B2(n_108),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_60),
.B(n_62),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_60),
.B(n_19),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_121),
.B1(n_123),
.B2(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_93),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_133),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_127),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_142),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_143),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_132),
.B1(n_134),
.B2(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_144),
.B1(n_146),
.B2(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.C(n_140),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_19),
.C(n_22),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_166),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_22),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_139),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_157),
.C(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_153),
.B1(n_158),
.B2(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_172),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_155),
.B1(n_159),
.B2(n_162),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_11),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_2),
.B(n_3),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_4),
.B(n_5),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_11),
.C(n_12),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_180),
.B1(n_5),
.B2(n_6),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_175),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_5),
.B(n_6),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_7),
.B(n_9),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_183),
.B(n_184),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.C(n_176),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_174),
.B(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_188),
.B(n_7),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_9),
.Y(n_192)
);


endmodule