module fake_jpeg_31557_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_16),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_50),
.Y(n_90)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_3),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_25),
.Y(n_64)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_62),
.B1(n_49),
.B2(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_67),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_68),
.B(n_74),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_39),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_51),
.B1(n_46),
.B2(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_98),
.B1(n_7),
.B2(n_13),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_100),
.Y(n_111)
);

OR2x4_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_6),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_85)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_92),
.B1(n_94),
.B2(n_4),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_38),
.B1(n_30),
.B2(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_23),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_101),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_27),
.B1(n_21),
.B2(n_17),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_39),
.B1(n_37),
.B2(n_32),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_37),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_5),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_32),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_43),
.B(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_43),
.B(n_8),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_11),
.Y(n_125)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx24_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_107),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_109),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_109),
.B1(n_135),
.B2(n_113),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_9),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_9),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_134),
.B1(n_86),
.B2(n_84),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_82),
.B(n_76),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_84),
.B(n_80),
.Y(n_142)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_130),
.Y(n_149)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_97),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_92),
.B1(n_86),
.B2(n_72),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_83),
.B(n_86),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_80),
.C(n_99),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_88),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_159),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_96),
.B1(n_70),
.B2(n_79),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_96),
.B1(n_70),
.B2(n_79),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_66),
.B1(n_135),
.B2(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_154),
.Y(n_169)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_110),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_157),
.B(n_118),
.Y(n_177)
);

AO22x2_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_110),
.B1(n_125),
.B2(n_129),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_143),
.B1(n_149),
.B2(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_107),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_118),
.B(n_107),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_170),
.B(n_145),
.Y(n_190)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_173),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_168),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_118),
.B(n_108),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_108),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_171),
.B(n_177),
.Y(n_204)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_185),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_148),
.A2(n_159),
.B1(n_136),
.B2(n_141),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_139),
.B1(n_156),
.B2(n_155),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_146),
.B(n_147),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_197),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_136),
.B(n_138),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_164),
.B(n_170),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_161),
.C(n_162),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_199),
.C(n_181),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_140),
.C(n_151),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_165),
.C(n_186),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_166),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_205),
.B1(n_179),
.B2(n_182),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_139),
.B1(n_165),
.B2(n_172),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_210),
.C(n_211),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_169),
.C(n_175),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_195),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_218),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_180),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_219),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_216),
.A2(n_203),
.B1(n_188),
.B2(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_184),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_194),
.B1(n_203),
.B2(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_215),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_201),
.B1(n_212),
.B2(n_190),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_209),
.C(n_211),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_187),
.C(n_202),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_191),
.B(n_193),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_228),
.A2(n_202),
.B(n_192),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_232),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_219),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_208),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_237),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_241),
.B(n_222),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_231),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_235),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_248),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_227),
.B1(n_221),
.B2(n_228),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_247),
.A2(n_242),
.B(n_192),
.C(n_198),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_221),
.B(n_176),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_244),
.B1(n_224),
.B2(n_176),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_251),
.A2(n_249),
.B(n_250),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_253),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_239),
.Y(n_256)
);


endmodule