module fake_jpeg_9823_n_274 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_26),
.B1(n_33),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_50),
.B1(n_54),
.B2(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_0),
.Y(n_95)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_23),
.B1(n_39),
.B2(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_25),
.B1(n_40),
.B2(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_26),
.B1(n_33),
.B2(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_37),
.B1(n_44),
.B2(n_22),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_67),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_65),
.B(n_69),
.Y(n_118)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2x1p5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_40),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_74),
.Y(n_113)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_42),
.B1(n_28),
.B2(n_29),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_18),
.B1(n_42),
.B2(n_31),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_24),
.B(n_22),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_87),
.B(n_90),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_82),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_18),
.B1(n_42),
.B2(n_31),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_37),
.C(n_35),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_37),
.B1(n_24),
.B2(n_34),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_35),
.B1(n_36),
.B2(n_45),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_22),
.B1(n_24),
.B2(n_34),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_95),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_56),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_35),
.B1(n_36),
.B2(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_2),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_116),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_34),
.C(n_45),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_90),
.C(n_86),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_127),
.B1(n_67),
.B2(n_71),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_84),
.A2(n_36),
.B1(n_34),
.B2(n_30),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_77),
.B(n_72),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_110),
.B(n_125),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_135),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_133),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_143),
.C(n_98),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_95),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_74),
.B1(n_63),
.B2(n_73),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_148),
.B1(n_156),
.B2(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_91),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_66),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_81),
.B(n_96),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_150),
.B(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_103),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_178),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_158),
.B(n_163),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_140),
.B1(n_152),
.B2(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_115),
.B1(n_70),
.B2(n_89),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_100),
.B(n_105),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_116),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_183),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_140),
.B1(n_148),
.B2(n_120),
.Y(n_185)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_121),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_156),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_175),
.B(n_36),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_182),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_101),
.B(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_147),
.C(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_195),
.B1(n_197),
.B2(n_200),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_193),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_133),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_205),
.C(n_159),
.Y(n_207)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_124),
.B1(n_120),
.B2(n_115),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_153),
.B1(n_124),
.B2(n_99),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_181),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_19),
.B1(n_10),
.B2(n_11),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_166),
.B1(n_167),
.B2(n_160),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_3),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_211),
.C(n_216),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_188),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_159),
.C(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_193),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_172),
.C(n_167),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_184),
.A2(n_166),
.B1(n_181),
.B2(n_165),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_200),
.B(n_201),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_161),
.C(n_176),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_SL g224 ( 
.A(n_206),
.B(n_202),
.C(n_205),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_227),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_230),
.Y(n_246)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_234),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_210),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_195),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_235),
.B(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_164),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_16),
.B(n_15),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_219),
.C(n_207),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_216),
.C(n_211),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_225),
.C(n_221),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_231),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_226),
.B1(n_230),
.B2(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_212),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_3),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_229),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_252),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_246),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_245),
.B(n_14),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_14),
.B(n_13),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_4),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_256),
.A2(n_238),
.B1(n_5),
.B2(n_6),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_254),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_246),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_253),
.B(n_238),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_241),
.C(n_240),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_262),
.C(n_259),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_266),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_260),
.C(n_261),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_4),
.C(n_5),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_5),
.B(n_6),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_7),
.C(n_8),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_9),
.B1(n_270),
.B2(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_9),
.Y(n_274)
);


endmodule