module fake_jpeg_16779_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx11_ASAP7_75t_SL g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_12),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_21),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_15),
.C(n_16),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_15),
.C(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_13),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_17),
.B(n_13),
.C(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_29),
.B1(n_18),
.B2(n_25),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_24),
.B1(n_34),
.B2(n_38),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_39),
.C(n_40),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_53),
.C(n_47),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_48),
.B1(n_14),
.B2(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_54),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_66),
.B(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_46),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_7),
.B(n_9),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_62),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_60),
.B(n_59),
.C(n_20),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_67),
.B(n_49),
.Y(n_72)
);

AOI221xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_71),
.B1(n_68),
.B2(n_43),
.C(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_74),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_28),
.C(n_38),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_37),
.B1(n_34),
.B2(n_28),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_77),
.C(n_7),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_9),
.Y(n_81)
);


endmodule