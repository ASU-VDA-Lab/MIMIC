module fake_jpeg_26827_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_28),
.B1(n_18),
.B2(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_28),
.B1(n_20),
.B2(n_19),
.Y(n_63)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_28),
.B1(n_19),
.B2(n_32),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_20),
.B1(n_32),
.B2(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_65),
.Y(n_103)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_68),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_39),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_74),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_41),
.B1(n_16),
.B2(n_17),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_24),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_81),
.B(n_87),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_40),
.B1(n_17),
.B2(n_24),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_67),
.B1(n_81),
.B2(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_78),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_88),
.B1(n_69),
.B2(n_81),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_25),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_85),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_83),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_22),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_21),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_4),
.C(n_5),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_30),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_21),
.B1(n_17),
.B2(n_26),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_43),
.B1(n_46),
.B2(n_55),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_90),
.A2(n_96),
.B1(n_97),
.B2(n_100),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_40),
.A3(n_26),
.B1(n_21),
.B2(n_17),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_72),
.C(n_77),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_93),
.B(n_98),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_20),
.B1(n_50),
.B2(n_30),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_34),
.B(n_40),
.C(n_57),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_0),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_107),
.C(n_76),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_62),
.B1(n_80),
.B2(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_77),
.Y(n_138)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_65),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_119),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_71),
.B(n_81),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_124),
.B(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_84),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_116),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_74),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_138),
.B(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_95),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_148),
.C(n_153),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_89),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_89),
.C(n_105),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_109),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_95),
.B1(n_105),
.B2(n_64),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_72),
.B1(n_5),
.B2(n_6),
.Y(n_182)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_159),
.B(n_75),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_98),
.C(n_102),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_129),
.C(n_137),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_90),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_139),
.C(n_133),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_124),
.C(n_102),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_174),
.C(n_179),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_178),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_130),
.B1(n_97),
.B2(n_91),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_159),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_113),
.C(n_114),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_67),
.B1(n_110),
.B2(n_72),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_70),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_70),
.C(n_72),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_166),
.C(n_167),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_188),
.C(n_195),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_163),
.C(n_144),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_150),
.B1(n_171),
.B2(n_186),
.Y(n_196)
);

BUFx12_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_150),
.B1(n_146),
.B2(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_140),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_151),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_163),
.C(n_141),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_200),
.B1(n_185),
.B2(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_152),
.B1(n_146),
.B2(n_176),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_180),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_184),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_154),
.B(n_142),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

OAI31xp33_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_141),
.A3(n_183),
.B(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_143),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_4),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_185),
.Y(n_209)
);

OAI31xp33_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_203),
.A3(n_200),
.B(n_191),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_204),
.B1(n_187),
.B2(n_143),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_216),
.B(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_5),
.Y(n_216)
);

AOI21x1_ASAP7_75t_SL g218 ( 
.A1(n_213),
.A2(n_210),
.B(n_206),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_219),
.B1(n_7),
.B2(n_10),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_222),
.A2(n_12),
.B(n_15),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_15),
.Y(n_224)
);


endmodule