module fake_ariane_930_n_188 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_188);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_188;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_159;
wire n_91;
wire n_107;
wire n_72;
wire n_128;
wire n_105;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_121;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

OR2x6_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_1),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

OR2x6_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_51),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_2),
.C(n_3),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_4),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_6),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_72),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_72),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_68),
.Y(n_76)
);

NAND2x1p5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_51),
.B1(n_50),
.B2(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_48),
.B(n_47),
.C(n_37),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_47),
.B1(n_43),
.B2(n_39),
.Y(n_88)
);

NOR2x1p5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_42),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_70),
.B(n_71),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_57),
.B(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_68),
.Y(n_94)
);

AO31x2_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_60),
.A3(n_65),
.B(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_76),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_65),
.B(n_60),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

OAI22x1_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_69),
.B1(n_66),
.B2(n_64),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_77),
.B(n_89),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_80),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_81),
.Y(n_106)
);

AOI21x1_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_87),
.B(n_88),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_83),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_98),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_119),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_103),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_103),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_101),
.B(n_112),
.Y(n_136)
);

OAI31xp33_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_111),
.A3(n_113),
.B(n_77),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_114),
.Y(n_140)
);

NAND3x1_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_131),
.C(n_127),
.Y(n_141)
);

NAND4xp25_ASAP7_75t_SL g142 ( 
.A(n_136),
.B(n_102),
.C(n_7),
.D(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

AOI222xp33_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_101),
.B1(n_64),
.B2(n_63),
.C1(n_114),
.C2(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_132),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_85),
.C(n_86),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_132),
.B(n_123),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_58),
.B1(n_124),
.B2(n_63),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_6),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_116),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_86),
.C(n_58),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_8),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_145),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_9),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_10),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_10),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_142),
.C(n_90),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_148),
.B(n_102),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_79),
.B(n_84),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_R g168 ( 
.A(n_158),
.B(n_11),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_159),
.A3(n_158),
.B1(n_153),
.B2(n_74),
.C1(n_73),
.C2(n_107),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_159),
.B1(n_74),
.B2(n_82),
.C(n_85),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_SL g171 ( 
.A(n_168),
.B(n_11),
.C(n_12),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_162),
.A2(n_82),
.A3(n_85),
.B1(n_99),
.B2(n_100),
.C1(n_105),
.C2(n_93),
.Y(n_172)
);

OAI211xp5_ASAP7_75t_SL g173 ( 
.A1(n_160),
.A2(n_91),
.B(n_93),
.C(n_105),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

OAI322xp33_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_85),
.A3(n_103),
.B1(n_95),
.B2(n_22),
.C1(n_23),
.C2(n_25),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g177 ( 
.A(n_175),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_162),
.B1(n_165),
.B2(n_168),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_103),
.B1(n_106),
.B2(n_85),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_14),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_106),
.C(n_95),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_177),
.B(n_181),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_176),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_173),
.B1(n_16),
.B2(n_26),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_15),
.B(n_27),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_182),
.B1(n_185),
.B2(n_184),
.C(n_186),
.Y(n_188)
);


endmodule