module fake_jpeg_16868_n_352 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_352);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_49),
.B1(n_47),
.B2(n_27),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_29),
.B1(n_21),
.B2(n_31),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_38),
.B1(n_26),
.B2(n_32),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_40),
.Y(n_79)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_29),
.B1(n_31),
.B2(n_17),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_17),
.B1(n_27),
.B2(n_22),
.Y(n_102)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_79),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_80),
.A2(n_84),
.B1(n_93),
.B2(n_94),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_51),
.B1(n_42),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_97),
.B1(n_100),
.B2(n_114),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_83),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_25),
.B1(n_49),
.B2(n_24),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_85),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_25),
.B1(n_49),
.B2(n_37),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_24),
.B1(n_37),
.B2(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_42),
.B1(n_44),
.B2(n_30),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_72),
.A2(n_32),
.B1(n_26),
.B2(n_45),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_112),
.B1(n_113),
.B2(n_41),
.Y(n_143)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_60),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_34),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_46),
.B1(n_45),
.B2(n_43),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_92),
.C(n_88),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_120),
.C(n_105),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_52),
.C(n_50),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_27),
.B1(n_17),
.B2(n_55),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_122),
.B(n_107),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_69),
.B1(n_36),
.B2(n_19),
.Y(n_122)
);

BUFx2_ASAP7_75t_SL g126 ( 
.A(n_76),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_54),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_108),
.B(n_106),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_89),
.A2(n_74),
.B1(n_53),
.B2(n_15),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_111),
.B1(n_87),
.B2(n_74),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_18),
.A3(n_41),
.B1(n_46),
.B2(n_43),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_89),
.B1(n_86),
.B2(n_98),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_111),
.B1(n_90),
.B2(n_110),
.Y(n_163)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_53),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_174),
.B(n_137),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_167),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_86),
.B1(n_101),
.B2(n_95),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_137),
.B1(n_129),
.B2(n_127),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_87),
.B1(n_90),
.B2(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_149),
.A2(n_151),
.B1(n_163),
.B2(n_173),
.Y(n_197)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_114),
.B1(n_99),
.B2(n_96),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_162),
.B1(n_169),
.B2(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_140),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_121),
.B(n_118),
.Y(n_179)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_157),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_120),
.C(n_130),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_111),
.B1(n_101),
.B2(n_87),
.Y(n_162)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_172),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_76),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_23),
.B(n_19),
.C(n_35),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_53),
.B1(n_68),
.B2(n_66),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_171),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_125),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_68),
.B1(n_66),
.B2(n_65),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_0),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_54),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_68),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_167),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_178),
.A2(n_186),
.B(n_190),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_179),
.A2(n_188),
.B(n_201),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_187),
.B1(n_204),
.B2(n_191),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_193),
.C(n_52),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_132),
.B(n_137),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_128),
.B1(n_134),
.B2(n_142),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_134),
.B(n_123),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_123),
.B(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_198),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_146),
.B1(n_172),
.B2(n_156),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_151),
.B(n_175),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_136),
.B1(n_144),
.B2(n_116),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_159),
.A2(n_54),
.B1(n_66),
.B2(n_65),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_205),
.A2(n_149),
.B1(n_160),
.B2(n_165),
.Y(n_211)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_50),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_SL g234 ( 
.A(n_206),
.B(n_35),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g207 ( 
.A(n_157),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_166),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_174),
.C(n_162),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_146),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_233),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_168),
.B(n_152),
.C(n_169),
.D(n_176),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_212),
.B(n_223),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_230),
.C(n_238),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_192),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_231),
.B1(n_235),
.B2(n_236),
.Y(n_241)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_161),
.A3(n_52),
.B1(n_65),
.B2(n_78),
.C1(n_116),
.C2(n_19),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_181),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_150),
.Y(n_226)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_161),
.B(n_36),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_234),
.B(n_190),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_199),
.B1(n_189),
.B2(n_208),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_161),
.C(n_78),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_36),
.B1(n_35),
.B2(n_23),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_184),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_191),
.A2(n_35),
.B1(n_23),
.B2(n_2),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_203),
.A2(n_35),
.B1(n_23),
.B2(n_2),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_23),
.C(n_16),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_15),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_16),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_15),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_179),
.C(n_205),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_248),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_252),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_177),
.B1(n_214),
.B2(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_249),
.B1(n_212),
.B2(n_239),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_178),
.C(n_184),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_255),
.C(n_257),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_200),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_185),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_197),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_197),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_180),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_261),
.C(n_227),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_226),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_0),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_180),
.C(n_198),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_177),
.B1(n_183),
.B2(n_209),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_262),
.A2(n_249),
.B1(n_240),
.B2(n_216),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_209),
.B(n_198),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_217),
.B(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_272),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_284),
.C(n_286),
.Y(n_288)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_270),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_263),
.A2(n_220),
.B1(n_232),
.B2(n_217),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_271),
.A2(n_278),
.B1(n_285),
.B2(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_233),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_279),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_211),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_280),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_241),
.B(n_252),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_210),
.B1(n_236),
.B2(n_13),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_264),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_13),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_0),
.C(n_1),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_250),
.A2(n_253),
.B1(n_259),
.B2(n_255),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_243),
.B(n_11),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_293),
.B(n_303),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_261),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_269),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_246),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_242),
.C(n_244),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_270),
.B1(n_281),
.B2(n_271),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_285),
.B(n_12),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_280),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_0),
.C(n_1),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_284),
.C(n_286),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_282),
.A2(n_2),
.B(n_3),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_12),
.Y(n_304)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_265),
.B1(n_274),
.B2(n_277),
.Y(n_306)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_317),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_309),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_289),
.A2(n_281),
.B1(n_11),
.B2(n_5),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_298),
.B(n_3),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_3),
.C(n_4),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_314),
.C(n_315),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_3),
.C(n_4),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_5),
.C(n_6),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_5),
.C(n_6),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_301),
.C(n_303),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_6),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_290),
.B(n_6),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_7),
.B(n_8),
.Y(n_330)
);

XOR2x1_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_292),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_289),
.B(n_295),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_300),
.B(n_297),
.Y(n_325)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_314),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_287),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_305),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_331),
.B(n_333),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_334),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_315),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_335),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_316),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_308),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_324),
.B1(n_326),
.B2(n_322),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_341),
.B(n_328),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_344),
.A2(n_345),
.B(n_342),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_335),
.Y(n_345)
);

AOI321xp33_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_346),
.A3(n_343),
.B1(n_336),
.B2(n_323),
.C(n_327),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_323),
.C(n_295),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_349),
.A2(n_9),
.B(n_10),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_9),
.C(n_10),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_10),
.Y(n_352)
);


endmodule