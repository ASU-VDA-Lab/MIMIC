module fake_jpeg_18386_n_144 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_77),
.A2(n_58),
.B1(n_64),
.B2(n_60),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_53),
.B1(n_52),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_65),
.B1(n_71),
.B2(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_56),
.B1(n_54),
.B2(n_46),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_62),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_70),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_70),
.B(n_55),
.C(n_54),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_94),
.B1(n_89),
.B2(n_85),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_96),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_69),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_99),
.B1(n_0),
.B2(n_2),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_63),
.B1(n_47),
.B2(n_26),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_3),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_116),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_23),
.B1(n_39),
.B2(n_38),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_107),
.B1(n_113),
.B2(n_115),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_21),
.B1(n_37),
.B2(n_35),
.Y(n_107)
);

NAND2x1_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_3),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_18),
.B1(n_33),
.B2(n_32),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_16),
.B1(n_31),
.B2(n_29),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_4),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_111),
.C(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_4),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_129),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_10),
.C(n_28),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_121),
.C(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_132),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_138),
.B(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_128),
.Y(n_140)
);

AOI21x1_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_130),
.B(n_6),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_22),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_40),
.C(n_6),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_5),
.Y(n_144)
);


endmodule