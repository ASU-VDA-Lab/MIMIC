module fake_netlist_1_2062_n_711 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_711);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_711;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_631;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_14), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_2), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_13), .Y(n_80) );
INVx1_ASAP7_75t_SL g81 ( .A(n_38), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_53), .Y(n_82) );
INVxp33_ASAP7_75t_L g83 ( .A(n_35), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_64), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_34), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_44), .Y(n_87) );
INVx1_ASAP7_75t_SL g88 ( .A(n_65), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_60), .Y(n_89) );
BUFx10_ASAP7_75t_L g90 ( .A(n_43), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_23), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
INVx3_ASAP7_75t_L g93 ( .A(n_59), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_21), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_33), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_0), .Y(n_97) );
CKINVDCx14_ASAP7_75t_R g98 ( .A(n_49), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_13), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_51), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_45), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_56), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_52), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_3), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_29), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_77), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_68), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_19), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_3), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_37), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_48), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_15), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_18), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_8), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_41), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_26), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_8), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_6), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_57), .Y(n_122) );
INVxp33_ASAP7_75t_L g123 ( .A(n_19), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_42), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_11), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_93), .B(n_1), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_123), .B(n_1), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_110), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
BUFx8_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_91), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_117), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_117), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_102), .B(n_4), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_87), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_108), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_111), .Y(n_151) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_124), .A2(n_39), .B(n_75), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_83), .B(n_5), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_82), .Y(n_155) );
INVx6_ASAP7_75t_L g156 ( .A(n_90), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_108), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_101), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_115), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_105), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_98), .B(n_78), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_107), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_115), .Y(n_165) );
BUFx2_ASAP7_75t_L g166 ( .A(n_104), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_112), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_78), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_131), .B(n_103), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_131), .B(n_103), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
NAND3x1_ASAP7_75t_L g176 ( .A(n_149), .B(n_84), .C(n_95), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
AND2x6_ASAP7_75t_L g180 ( .A(n_163), .B(n_84), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_156), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_126), .B(n_106), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_156), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_129), .A2(n_122), .B1(n_125), .B2(n_99), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_126), .B(n_118), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_149), .A2(n_121), .B1(n_119), .B2(n_95), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_126), .B(n_106), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_147), .Y(n_190) );
AND3x4_ASAP7_75t_L g191 ( .A(n_157), .B(n_10), .C(n_11), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_127), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_127), .Y(n_193) );
AO22x2_ASAP7_75t_L g194 ( .A1(n_163), .A2(n_121), .B1(n_119), .B2(n_116), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_142), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_143), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_166), .B(n_118), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_166), .B(n_113), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_157), .A2(n_114), .B1(n_109), .B2(n_97), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_153), .B(n_80), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_165), .B(n_79), .Y(n_205) );
BUFx10_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_136), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_132), .B(n_133), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_131), .B(n_96), .Y(n_212) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_153), .B(n_96), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
AO22x2_ASAP7_75t_L g215 ( .A1(n_132), .A2(n_86), .B1(n_88), .B2(n_81), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_131), .B(n_46), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_158), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_133), .B(n_47), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_162), .B(n_12), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_162), .B(n_40), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_162), .B(n_50), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_150), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_129), .B(n_12), .Y(n_224) );
OR2x2_ASAP7_75t_L g225 ( .A(n_162), .B(n_146), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_137), .B(n_14), .Y(n_226) );
NAND2xp33_ASAP7_75t_L g227 ( .A(n_155), .B(n_54), .Y(n_227) );
INVx6_ASAP7_75t_L g228 ( .A(n_158), .Y(n_228) );
AND2x6_ASAP7_75t_L g229 ( .A(n_137), .B(n_55), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_138), .B(n_15), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_158), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_212), .B(n_136), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_210), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_210), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_228), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_228), .Y(n_237) );
INVx5_ASAP7_75t_L g238 ( .A(n_229), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_212), .B(n_136), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_226), .A2(n_144), .B1(n_141), .B2(n_139), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_226), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_180), .A2(n_136), .B1(n_167), .B2(n_161), .Y(n_242) );
BUFx2_ASAP7_75t_SL g243 ( .A(n_206), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
BUFx4f_ASAP7_75t_L g245 ( .A(n_180), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_199), .B(n_155), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_173), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_172), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_230), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_230), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_170), .B(n_159), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_225), .B(n_144), .Y(n_254) );
INVx1_ASAP7_75t_SL g255 ( .A(n_177), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_172), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_209), .B(n_159), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_206), .B(n_161), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_220), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_213), .B(n_167), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_180), .B(n_140), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_182), .B(n_140), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_194), .B(n_141), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_194), .B(n_139), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_182), .B(n_145), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_187), .B(n_145), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_169), .B(n_138), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_178), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_187), .B(n_148), .Y(n_269) );
AND2x6_ASAP7_75t_L g270 ( .A(n_172), .B(n_148), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_184), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g272 ( .A1(n_188), .A2(n_168), .B(n_128), .C(n_150), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_174), .B(n_164), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_193), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_189), .B(n_164), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_215), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_189), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_171), .B(n_164), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_195), .Y(n_279) );
NAND2x1_ASAP7_75t_L g280 ( .A(n_229), .B(n_168), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_192), .Y(n_281) );
BUFx4f_ASAP7_75t_L g282 ( .A(n_202), .Y(n_282) );
BUFx12f_ASAP7_75t_L g283 ( .A(n_224), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_179), .Y(n_284) );
OR2x6_ASAP7_75t_L g285 ( .A(n_224), .B(n_168), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_202), .Y(n_286) );
AND2x6_ASAP7_75t_SL g287 ( .A(n_190), .B(n_16), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_185), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_202), .B(n_134), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_202), .B(n_186), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_218), .A2(n_134), .B(n_130), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_200), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_196), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_175), .B(n_134), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_181), .B(n_158), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_205), .B(n_130), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_185), .Y(n_297) );
AOI22xp5_ASAP7_75t_SL g298 ( .A1(n_201), .A2(n_135), .B1(n_17), .B2(n_18), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_186), .B(n_130), .Y(n_299) );
INVx3_ASAP7_75t_SL g300 ( .A(n_215), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_247), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_285), .B(n_183), .Y(n_302) );
AOI22xp5_ASAP7_75t_SL g303 ( .A1(n_288), .A2(n_201), .B1(n_191), .B2(n_229), .Y(n_303) );
BUFx12f_ASAP7_75t_L g304 ( .A(n_287), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_234), .A2(n_214), .B(n_197), .C(n_198), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_255), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_262), .A2(n_179), .B(n_218), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_292), .B(n_194), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_235), .B(n_215), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_272), .A2(n_223), .B(n_207), .C(n_204), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_251), .Y(n_312) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_245), .B(n_203), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_251), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_254), .B(n_188), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_240), .A2(n_176), .B1(n_179), .B2(n_222), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_285), .B(n_229), .Y(n_317) );
BUFx4f_ASAP7_75t_L g318 ( .A(n_285), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_265), .A2(n_269), .B(n_266), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_300), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_245), .Y(n_321) );
NOR2xp33_ASAP7_75t_SL g322 ( .A(n_300), .B(n_221), .Y(n_322) );
BUFx12f_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
INVx3_ASAP7_75t_SL g324 ( .A(n_270), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_248), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_270), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_243), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_248), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_268), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_272), .A2(n_222), .B(n_221), .C(n_135), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_246), .B(n_216), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_291), .A2(n_227), .B(n_208), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_276), .Y(n_334) );
AND2x4_ASAP7_75t_SL g335 ( .A(n_240), .B(n_135), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_270), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_260), .A2(n_219), .B(n_217), .C(n_232), .Y(n_337) );
NOR2xp33_ASAP7_75t_SL g338 ( .A(n_282), .B(n_135), .Y(n_338) );
INVx2_ASAP7_75t_SL g339 ( .A(n_253), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_275), .A2(n_231), .B(n_211), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_277), .A2(n_231), .B1(n_211), .B2(n_16), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_271), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_257), .B(n_17), .Y(n_343) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_296), .A2(n_231), .B(n_211), .C(n_24), .Y(n_344) );
CKINVDCx8_ASAP7_75t_R g345 ( .A(n_253), .Y(n_345) );
OAI221xp5_ASAP7_75t_L g346 ( .A1(n_296), .A2(n_20), .B1(n_22), .B2(n_27), .C(n_28), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_263), .B(n_30), .Y(n_347) );
BUFx12f_ASAP7_75t_L g348 ( .A(n_294), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_233), .A2(n_31), .B(n_32), .Y(n_349) );
NAND2x1_ASAP7_75t_SL g350 ( .A(n_242), .B(n_36), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_241), .A2(n_58), .B1(n_61), .B2(n_62), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_282), .Y(n_352) );
BUFx12f_ASAP7_75t_L g353 ( .A(n_294), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_329), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_331), .A2(n_291), .B(n_239), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_301), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_330), .A2(n_264), .B1(n_250), .B2(n_252), .Y(n_357) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_331), .A2(n_289), .B(n_261), .Y(n_358) );
BUFx3_ASAP7_75t_L g359 ( .A(n_324), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_324), .Y(n_360) );
CKINVDCx9p33_ASAP7_75t_R g361 ( .A(n_310), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_349), .A2(n_280), .B(n_295), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_342), .Y(n_363) );
AO21x1_ASAP7_75t_L g364 ( .A1(n_309), .A2(n_273), .B(n_279), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_267), .B1(n_259), .B2(n_273), .C(n_293), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_301), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_307), .A2(n_290), .B(n_299), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_330), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_326), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_350), .A2(n_274), .B(n_258), .Y(n_372) );
INVxp33_ASAP7_75t_L g373 ( .A(n_303), .Y(n_373) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_344), .B(n_298), .C(n_238), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_317), .B(n_238), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g376 ( .A1(n_311), .A2(n_267), .B(n_286), .C(n_249), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_319), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_340), .A2(n_278), .B(n_281), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g379 ( .A1(n_316), .A2(n_322), .B(n_343), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_286), .B1(n_249), .B2(n_281), .C(n_238), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_311), .A2(n_256), .B(n_248), .Y(n_381) );
NOR2x1p5_ASAP7_75t_L g382 ( .A(n_310), .B(n_238), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_325), .A2(n_284), .B(n_256), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_305), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_328), .A2(n_284), .B(n_256), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_308), .B(n_270), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_373), .A2(n_348), .B1(n_353), .B2(n_343), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_370), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_370), .A2(n_318), .B1(n_306), .B2(n_348), .Y(n_389) );
OAI22xp33_ASAP7_75t_SL g390 ( .A1(n_354), .A2(n_318), .B1(n_334), .B2(n_327), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_354), .B(n_323), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_359), .A2(n_327), .B1(n_320), .B2(n_339), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_365), .A2(n_332), .B1(n_317), .B2(n_302), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_363), .Y(n_394) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_379), .A2(n_335), .B(n_332), .C(n_305), .Y(n_395) );
INVxp33_ASAP7_75t_SL g396 ( .A(n_361), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_382), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_357), .A2(n_335), .B1(n_302), .B2(n_347), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
OA21x2_ASAP7_75t_L g401 ( .A1(n_381), .A2(n_344), .B(n_328), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_382), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_356), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_366), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_379), .A2(n_341), .B(n_346), .C(n_312), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_365), .A2(n_314), .B1(n_313), .B2(n_351), .C(n_337), .Y(n_408) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_375), .B(n_338), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_366), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_384), .A2(n_352), .B1(n_321), .B2(n_333), .C(n_313), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_384), .A2(n_304), .B1(n_321), .B2(n_333), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_381), .A2(n_248), .B(n_284), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_336), .B(n_244), .C(n_237), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_388), .B(n_364), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_394), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_400), .B(n_377), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_400), .B(n_377), .Y(n_418) );
NOR2x1p5_ASAP7_75t_L g419 ( .A(n_396), .B(n_374), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_388), .B(n_364), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_403), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_409), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_405), .B(n_358), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_405), .B(n_358), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_407), .B(n_375), .Y(n_425) );
OR2x6_ASAP7_75t_L g426 ( .A(n_399), .B(n_359), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_394), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_403), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_407), .B(n_358), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_410), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_398), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_410), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_398), .B(n_364), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_404), .B(n_393), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_396), .A2(n_359), .B1(n_375), .B2(n_360), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_412), .B(n_358), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
NOR2xp67_ASAP7_75t_L g440 ( .A(n_402), .B(n_360), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_389), .B(n_358), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_387), .B(n_355), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_401), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_391), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_390), .B(n_386), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_395), .B(n_355), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_402), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_392), .B(n_355), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_406), .B(n_386), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_423), .B(n_355), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_417), .B(n_411), .Y(n_452) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_438), .A2(n_413), .B(n_385), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_417), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_438), .Y(n_455) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_419), .B(n_414), .Y(n_456) );
NAND2x1_ASAP7_75t_L g457 ( .A(n_426), .B(n_367), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_438), .Y(n_458) );
AOI21xp33_ASAP7_75t_L g459 ( .A1(n_442), .A2(n_408), .B(n_376), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_416), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_423), .B(n_368), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_436), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_421), .A2(n_383), .B(n_385), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_424), .B(n_372), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_424), .B(n_368), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_436), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_418), .B(n_386), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
BUFx3_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_439), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_450), .A2(n_397), .B1(n_375), .B2(n_380), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_439), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_429), .B(n_368), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_443), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_422), .A2(n_375), .B1(n_360), .B2(n_372), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_429), .B(n_372), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_443), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_434), .A2(n_376), .B1(n_380), .B2(n_371), .C(n_361), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_418), .B(n_369), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_431), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_446), .B(n_385), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_434), .A2(n_371), .B1(n_367), .B2(n_236), .C(n_336), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_421), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_421), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_428), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_435), .B(n_367), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_442), .B(n_369), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_433), .Y(n_493) );
AOI33xp33_ASAP7_75t_L g494 ( .A1(n_450), .A2(n_63), .A3(n_66), .B1(n_69), .B2(n_70), .B3(n_71), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_446), .B(n_432), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_428), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_430), .B(n_369), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_433), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_430), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_432), .B(n_378), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_425), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_460), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_451), .B(n_437), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_454), .B(n_415), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_477), .Y(n_505) );
INVx4_ASAP7_75t_L g506 ( .A(n_487), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_487), .B(n_449), .Y(n_507) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_494), .A2(n_419), .B(n_440), .C(n_447), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_454), .B(n_415), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_461), .B(n_425), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_490), .B(n_420), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_493), .A2(n_445), .B1(n_448), .B2(n_449), .C(n_444), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_490), .B(n_420), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_464), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_472), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_464), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_467), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_467), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_471), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_461), .B(n_425), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_461), .B(n_447), .Y(n_522) );
INVx6_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_471), .Y(n_524) );
NAND4xp25_ASAP7_75t_L g525 ( .A(n_481), .B(n_441), .C(n_440), .D(n_437), .Y(n_525) );
OAI211xp5_ASAP7_75t_L g526 ( .A1(n_481), .A2(n_441), .B(n_448), .C(n_444), .Y(n_526) );
BUFx2_ASAP7_75t_L g527 ( .A(n_472), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_466), .B(n_448), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_483), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_483), .B(n_448), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_451), .B(n_426), .Y(n_531) );
OAI31xp33_ASAP7_75t_L g532 ( .A1(n_491), .A2(n_371), .A3(n_426), .B(n_448), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_451), .B(n_426), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_466), .B(n_367), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_466), .B(n_367), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_488), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_488), .Y(n_537) );
NAND5xp2_ASAP7_75t_SL g538 ( .A(n_474), .B(n_72), .C(n_73), .D(n_74), .E(n_76), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
NOR2xp33_ASAP7_75t_R g540 ( .A(n_487), .B(n_367), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_493), .B(n_378), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_476), .B(n_367), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_452), .B(n_378), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_487), .B(n_383), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_498), .B(n_362), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_498), .B(n_362), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_476), .B(n_383), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_452), .B(n_362), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_487), .B(n_256), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_477), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_482), .B(n_284), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_480), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_482), .B(n_270), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_476), .B(n_469), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_501), .B(n_469), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_501), .B(n_482), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_480), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_495), .B(n_479), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_554), .B(n_486), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_502), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_509), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_559), .B(n_495), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_557), .B(n_486), .Y(n_566) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_540), .B(n_491), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_559), .B(n_495), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_532), .B(n_478), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_503), .B(n_479), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_510), .B(n_470), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_504), .B(n_479), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_527), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_503), .B(n_497), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_515), .B(n_497), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_531), .B(n_465), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_531), .B(n_465), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_506), .B(n_457), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_505), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_505), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_519), .B(n_497), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_512), .B(n_486), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_539), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_520), .B(n_470), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_540), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_514), .B(n_486), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_511), .B(n_486), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_524), .B(n_459), .Y(n_590) );
AOI211xp5_ASAP7_75t_SL g591 ( .A1(n_526), .A2(n_459), .B(n_492), .C(n_485), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_533), .B(n_465), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_506), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_529), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_536), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_533), .B(n_465), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_526), .B(n_478), .Y(n_597) );
OAI22xp33_ASAP7_75t_SL g598 ( .A1(n_506), .A2(n_457), .B1(n_501), .B2(n_456), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_537), .B(n_492), .Y(n_599) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_508), .B(n_456), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_521), .B(n_492), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_528), .B(n_465), .Y(n_602) );
NOR2x1p5_ASAP7_75t_L g603 ( .A(n_525), .B(n_455), .Y(n_603) );
NOR2x1p5_ASAP7_75t_L g604 ( .A(n_507), .B(n_455), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_516), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_555), .B(n_499), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_507), .B(n_516), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_539), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_543), .B(n_455), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_550), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_552), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_556), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_522), .B(n_489), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_543), .B(n_455), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_563), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_593), .A2(n_523), .B1(n_507), .B2(n_544), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_573), .B(n_508), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_SL g618 ( .A1(n_569), .A2(n_597), .B(n_587), .C(n_591), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_590), .B(n_548), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_564), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_569), .A2(n_523), .B1(n_474), .B2(n_513), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_565), .B(n_523), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_578), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_568), .B(n_548), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_568), .B(n_558), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_582), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_594), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_595), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_570), .B(n_561), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_570), .B(n_560), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_571), .B(n_530), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g632 ( .A1(n_597), .A2(n_544), .A3(n_553), .B(n_484), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_610), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_576), .B(n_542), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_611), .Y(n_635) );
AOI211x1_ASAP7_75t_SL g636 ( .A1(n_586), .A2(n_546), .B(n_545), .C(n_541), .Y(n_636) );
OAI22x1_ASAP7_75t_L g637 ( .A1(n_603), .A2(n_544), .B1(n_549), .B2(n_484), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_593), .A2(n_535), .B1(n_534), .B2(n_458), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_593), .A2(n_549), .B(n_485), .C(n_553), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_612), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_571), .B(n_547), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_572), .B(n_455), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_600), .A2(n_484), .B1(n_551), .B2(n_458), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_567), .A2(n_614), .B1(n_609), .B2(n_607), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_574), .B(n_489), .Y(n_645) );
OAI22xp33_ASAP7_75t_SL g646 ( .A1(n_605), .A2(n_549), .B1(n_458), .B2(n_489), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_613), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_599), .B(n_458), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_606), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g650 ( .A1(n_567), .A2(n_463), .B(n_551), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_598), .A2(n_463), .B(n_538), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_618), .A2(n_576), .B(n_596), .C(n_592), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_621), .A2(n_579), .B1(n_607), .B2(n_604), .Y(n_653) );
XNOR2xp5_ASAP7_75t_L g654 ( .A(n_641), .B(n_602), .Y(n_654) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_617), .B(n_579), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_633), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
NAND2xp33_ASAP7_75t_L g658 ( .A(n_637), .B(n_562), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_635), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_625), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_640), .Y(n_661) );
AOI221x1_ASAP7_75t_SL g662 ( .A1(n_619), .A2(n_607), .B1(n_579), .B2(n_583), .C(n_575), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_646), .A2(n_585), .B(n_584), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_624), .B(n_592), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_SL g665 ( .A1(n_639), .A2(n_566), .B(n_601), .C(n_589), .Y(n_665) );
AOI211xp5_ASAP7_75t_SL g666 ( .A1(n_638), .A2(n_596), .B(n_577), .C(n_588), .Y(n_666) );
XNOR2x1_ASAP7_75t_L g667 ( .A(n_644), .B(n_577), .Y(n_667) );
INVx1_ASAP7_75t_SL g668 ( .A(n_647), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_632), .A2(n_608), .B(n_581), .C(n_580), .Y(n_669) );
XNOR2xp5_ASAP7_75t_L g670 ( .A(n_649), .B(n_602), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_651), .B(n_608), .C(n_581), .Y(n_671) );
XNOR2xp5_ASAP7_75t_L g672 ( .A(n_631), .B(n_580), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_615), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_620), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_668), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_660), .Y(n_676) );
OA211x2_ASAP7_75t_L g677 ( .A1(n_653), .A2(n_650), .B(n_622), .C(n_616), .Y(n_677) );
OAI211xp5_ASAP7_75t_L g678 ( .A1(n_653), .A2(n_616), .B(n_643), .C(n_651), .Y(n_678) );
AOI31xp33_ASAP7_75t_L g679 ( .A1(n_652), .A2(n_638), .A3(n_630), .B(n_629), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_656), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_666), .A2(n_645), .B1(n_628), .B2(n_627), .Y(n_681) );
A2O1A1Ixp33_ASAP7_75t_L g682 ( .A1(n_662), .A2(n_634), .B(n_623), .C(n_626), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_657), .B(n_642), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_665), .A2(n_648), .B(n_499), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_655), .B(n_484), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_657), .A2(n_484), .B1(n_458), .B2(n_500), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_671), .A2(n_636), .B1(n_499), .B2(n_496), .Y(n_687) );
NAND2xp33_ASAP7_75t_SL g688 ( .A(n_667), .B(n_462), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_681), .B(n_671), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_677), .A2(n_658), .B1(n_672), .B2(n_663), .Y(n_690) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_678), .A2(n_669), .B1(n_674), .B2(n_661), .C(n_673), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_676), .B(n_659), .Y(n_692) );
AOI211xp5_ASAP7_75t_L g693 ( .A1(n_681), .A2(n_654), .B(n_670), .C(n_664), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_679), .A2(n_500), .B1(n_462), .B2(n_468), .C(n_473), .Y(n_694) );
NAND5xp2_ASAP7_75t_L g695 ( .A(n_687), .B(n_500), .C(n_453), .D(n_468), .E(n_473), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_675), .B(n_462), .Y(n_696) );
NOR2xp67_ASAP7_75t_L g697 ( .A(n_690), .B(n_684), .Y(n_697) );
NAND3xp33_ASAP7_75t_SL g698 ( .A(n_693), .B(n_688), .C(n_687), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_691), .A2(n_682), .B1(n_683), .B2(n_685), .Y(n_699) );
AND3x4_ASAP7_75t_L g700 ( .A(n_689), .B(n_686), .C(n_680), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_699), .A2(n_692), .B1(n_696), .B2(n_694), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_697), .B(n_695), .Y(n_702) );
INVx2_ASAP7_75t_SL g703 ( .A(n_700), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_703), .Y(n_704) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_702), .A2(n_698), .B(n_453), .Y(n_705) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_704), .B(n_701), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_705), .A2(n_468), .B1(n_473), .B2(n_475), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_706), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_707), .B(n_453), .Y(n_709) );
XNOR2xp5_ASAP7_75t_L g710 ( .A(n_709), .B(n_453), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_710), .A2(n_453), .B1(n_475), .B2(n_708), .Y(n_711) );
endmodule