module fake_jpeg_31374_n_507 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_507);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_507;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_70),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_22),
.B(n_3),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_36),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_3),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_92),
.Y(n_142)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_93),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_22),
.B(n_3),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_33),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_47),
.B1(n_51),
.B2(n_29),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_27),
.B1(n_50),
.B2(n_41),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_106),
.A2(n_129),
.B1(n_148),
.B2(n_165),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_112),
.B(n_43),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_27),
.B1(n_50),
.B2(n_41),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_31),
.B(n_49),
.C(n_48),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_128),
.B(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_50),
.Y(n_131)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_54),
.B(n_33),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_R g210 ( 
.A(n_132),
.B(n_36),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_41),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_51),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_96),
.A2(n_47),
.B1(n_49),
.B2(n_48),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_75),
.B(n_51),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_159),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_75),
.B(n_20),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_52),
.A2(n_20),
.B1(n_48),
.B2(n_45),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_168),
.B(n_181),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_119),
.A2(n_93),
.B1(n_45),
.B2(n_38),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_170),
.Y(n_248)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_178),
.Y(n_225)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_113),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_125),
.A2(n_61),
.B1(n_103),
.B2(n_74),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_179),
.A2(n_193),
.B1(n_194),
.B2(n_206),
.Y(n_243)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_31),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_183),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_184),
.B(n_189),
.Y(n_223)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_185),
.Y(n_264)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_119),
.Y(n_189)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_130),
.A2(n_88),
.B1(n_101),
.B2(n_100),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_111),
.A2(n_71),
.B1(n_98),
.B2(n_95),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

BUFx4f_ASAP7_75t_SL g261 ( 
.A(n_196),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_105),
.C(n_78),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_221),
.C(n_20),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_121),
.B(n_38),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_214),
.Y(n_231)
);

INVx13_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_109),
.Y(n_200)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_122),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_210),
.Y(n_232)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_68),
.B1(n_65),
.B2(n_64),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_207),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_136),
.A2(n_49),
.B1(n_45),
.B2(n_44),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_208),
.A2(n_218),
.B1(n_25),
.B2(n_142),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_215),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_120),
.A2(n_44),
.B1(n_43),
.B2(n_38),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_135),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_124),
.B(n_44),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_30),
.B(n_25),
.Y(n_251)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_217),
.A2(n_219),
.B1(n_220),
.B2(n_203),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_136),
.A2(n_43),
.B1(n_29),
.B2(n_31),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_141),
.B(n_30),
.C(n_29),
.Y(n_221)
);

OAI22x1_ASAP7_75t_SL g235 ( 
.A1(n_171),
.A2(n_148),
.B1(n_129),
.B2(n_147),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_235),
.A2(n_206),
.B1(n_197),
.B2(n_190),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_108),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_252),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

OAI22x1_ASAP7_75t_R g249 ( 
.A1(n_184),
.A2(n_142),
.B1(n_147),
.B2(n_120),
.Y(n_249)
);

AO22x1_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_176),
.B1(n_156),
.B2(n_186),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_21),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_168),
.B(n_25),
.C(n_30),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_172),
.C(n_175),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_263),
.B1(n_166),
.B2(n_110),
.Y(n_287)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_198),
.A2(n_36),
.B(n_5),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_4),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_108),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_260),
.B(n_183),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_195),
.A2(n_118),
.B1(n_160),
.B2(n_166),
.Y(n_263)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_223),
.A2(n_192),
.B(n_221),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_266),
.A2(n_271),
.B(n_272),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_202),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_274),
.C(n_254),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_268),
.A2(n_276),
.B(n_283),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_298),
.B1(n_232),
.B2(n_263),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_167),
.B(n_174),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_222),
.A2(n_205),
.B(n_220),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_185),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_222),
.A2(n_177),
.B(n_212),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_282),
.B(n_284),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_235),
.A2(n_182),
.B(n_180),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_286),
.Y(n_333)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_287),
.A2(n_290),
.B1(n_296),
.B2(n_236),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_252),
.Y(n_304)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_291),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_249),
.B1(n_239),
.B2(n_257),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_233),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_300),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_246),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_295),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_243),
.A2(n_160),
.B1(n_118),
.B2(n_204),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_199),
.C(n_196),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_288),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_239),
.A2(n_140),
.B1(n_143),
.B2(n_164),
.Y(n_298)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_241),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_231),
.B(n_191),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_304),
.B(n_309),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_321),
.B1(n_265),
.B2(n_275),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_295),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_310),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_240),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_312),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_232),
.C(n_260),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g339 ( 
.A1(n_313),
.A2(n_287),
.B1(n_296),
.B2(n_276),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_269),
.A2(n_253),
.B1(n_224),
.B2(n_143),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_314),
.A2(n_316),
.B1(n_324),
.B2(n_305),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_256),
.B1(n_259),
.B2(n_209),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_317),
.B(n_323),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_325),
.B1(n_298),
.B2(n_272),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_299),
.A2(n_245),
.B1(n_230),
.B2(n_228),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_297),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_293),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_299),
.A2(n_259),
.B1(n_238),
.B2(n_262),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_290),
.A2(n_156),
.B1(n_262),
.B2(n_244),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_244),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_332),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_281),
.A2(n_245),
.B1(n_230),
.B2(n_228),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_330),
.A2(n_248),
.B(n_234),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_238),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_285),
.B(n_266),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g372 ( 
.A1(n_334),
.A2(n_338),
.B(n_340),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_318),
.A2(n_270),
.B1(n_325),
.B2(n_313),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_336),
.A2(n_337),
.B1(n_358),
.B2(n_330),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_320),
.A2(n_313),
.B(n_333),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g382 ( 
.A1(n_339),
.A2(n_348),
.B(n_356),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_333),
.B(n_319),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_248),
.C(n_201),
.Y(n_381)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_344),
.A2(n_351),
.B1(n_307),
.B2(n_328),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_346),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_268),
.B(n_277),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_355),
.Y(n_369)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_302),
.B(n_267),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_352),
.Y(n_374)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_354),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_294),
.Y(n_355)
);

AO32x1_ASAP7_75t_L g356 ( 
.A1(n_306),
.A2(n_297),
.A3(n_292),
.B1(n_279),
.B2(n_280),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_316),
.B1(n_302),
.B2(n_324),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_306),
.B(n_286),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_359),
.Y(n_390)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_361),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_301),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_311),
.A2(n_291),
.B1(n_289),
.B2(n_265),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_362),
.A2(n_363),
.B1(n_327),
.B2(n_312),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_322),
.A2(n_250),
.B1(n_234),
.B2(n_227),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_331),
.A2(n_326),
.B(n_315),
.Y(n_364)
);

AO22x1_ASAP7_75t_SL g365 ( 
.A1(n_364),
.A2(n_315),
.B1(n_310),
.B2(n_304),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_365),
.B(n_340),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_367),
.A2(n_373),
.B1(n_380),
.B2(n_384),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_304),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_391),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_301),
.B1(n_328),
.B2(n_332),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_362),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_327),
.Y(n_378)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g396 ( 
.A(n_379),
.B(n_348),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_343),
.A2(n_309),
.B1(n_250),
.B2(n_227),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_386),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_357),
.B1(n_339),
.B2(n_356),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_336),
.A2(n_188),
.B1(n_170),
.B2(n_261),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_385),
.A2(n_393),
.B1(n_353),
.B2(n_354),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_261),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_4),
.Y(n_387)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_387),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_36),
.C(n_21),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_388),
.B(n_392),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_36),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_21),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_36),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_21),
.C(n_7),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_339),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_393)
);

OA22x2_ASAP7_75t_L g394 ( 
.A1(n_384),
.A2(n_337),
.B1(n_364),
.B2(n_339),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_394),
.A2(n_365),
.B1(n_392),
.B2(n_370),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_396),
.A2(n_411),
.B1(n_413),
.B2(n_385),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_374),
.B(n_335),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_408),
.Y(n_425)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_368),
.B(n_338),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_419),
.Y(n_420)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_335),
.C(n_334),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_412),
.Y(n_433)
);

XOR2x1_ASAP7_75t_SL g411 ( 
.A(n_382),
.B(n_347),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_369),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_345),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_414),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_393),
.A2(n_360),
.B1(n_8),
.B2(n_9),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_415),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_6),
.Y(n_416)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_417),
.B(n_418),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_369),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_397),
.C(n_386),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_428),
.C(n_430),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_372),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_429),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_381),
.C(n_380),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_389),
.C(n_377),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_403),
.A2(n_372),
.B(n_367),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_431),
.A2(n_394),
.B(n_395),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_391),
.C(n_373),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_435),
.B(n_410),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_388),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_419),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_439),
.A2(n_383),
.B1(n_9),
.B2(n_10),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_401),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_442),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_402),
.Y(n_441)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_441),
.Y(n_460)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_433),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_444),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_423),
.A2(n_416),
.B(n_400),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_408),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_445),
.B(n_447),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_432),
.A2(n_417),
.B1(n_394),
.B2(n_396),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_436),
.A2(n_394),
.B1(n_413),
.B2(n_371),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_448),
.A2(n_431),
.B1(n_432),
.B2(n_424),
.Y(n_462)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_438),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_449),
.B(n_450),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_410),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_451),
.B(n_453),
.Y(n_457)
);

NOR2x1_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_437),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_454),
.A2(n_420),
.B1(n_429),
.B2(n_430),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_455),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_465)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_456),
.B(n_11),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_462),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_455),
.A2(n_434),
.B1(n_435),
.B2(n_428),
.Y(n_463)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_463),
.Y(n_476)
);

OAI321xp33_ASAP7_75t_L g464 ( 
.A1(n_441),
.A2(n_434),
.A3(n_420),
.B1(n_421),
.B2(n_11),
.C(n_12),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_12),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_466),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_21),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_469),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_445),
.B(n_12),
.Y(n_469)
);

INVx11_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_446),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_471),
.A2(n_452),
.B(n_454),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_481),
.B(n_467),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_459),
.Y(n_490)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_478),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_446),
.C(n_453),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_483),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_460),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_482),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_461),
.A2(n_13),
.B(n_14),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_13),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_21),
.C(n_14),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_487),
.B(n_489),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_458),
.Y(n_488)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_488),
.Y(n_495)
);

AO21x1_ASAP7_75t_L g498 ( 
.A1(n_490),
.A2(n_465),
.B(n_14),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_470),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_491),
.B(n_468),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_473),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_492),
.A2(n_479),
.B1(n_476),
.B2(n_483),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_494),
.Y(n_499)
);

NOR3xp33_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_477),
.C(n_474),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_497),
.Y(n_500)
);

O2A1O1Ixp33_ASAP7_75t_SL g501 ( 
.A1(n_498),
.A2(n_484),
.B(n_485),
.C(n_15),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_495),
.B(n_496),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_503),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_499),
.A2(n_500),
.B(n_490),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g505 ( 
.A1(n_504),
.A2(n_497),
.B(n_14),
.C(n_16),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_505),
.B(n_13),
.C(n_16),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_16),
.Y(n_507)
);


endmodule