module fake_jpeg_13697_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_59),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_70),
.Y(n_78)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_1),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_56),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_54),
.B1(n_57),
.B2(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_57),
.B1(n_52),
.B2(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_52),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_100),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_47),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_92),
.Y(n_106)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_44),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_48),
.B1(n_58),
.B2(n_53),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_102),
.B(n_6),
.Y(n_114)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_5),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_53),
.B1(n_46),
.B2(n_45),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_98),
.A2(n_74),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_118),
.B1(n_32),
.B2(n_33),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_108),
.B1(n_114),
.B2(n_18),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_112),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_26),
.B(n_40),
.C(n_39),
.D(n_11),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_31),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_14),
.C(n_15),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_124),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

AND2x4_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_28),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_106),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_108),
.B1(n_104),
.B2(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_138),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_128),
.C(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_121),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_141),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_122),
.B(n_137),
.C(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_128),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_136),
.B(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_138),
.B1(n_126),
.B2(n_142),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_34),
.B(n_37),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_42),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_38),
.Y(n_150)
);


endmodule