module fake_jpeg_31976_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_9),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_13),
.B1(n_18),
.B2(n_16),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_14),
.B1(n_22),
.B2(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_9),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_21),
.C(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_38),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_26),
.B(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_33),
.B1(n_34),
.B2(n_15),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_12),
.B1(n_11),
.B2(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_14),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_36),
.C(n_34),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.C(n_52),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_51),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_39),
.C(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_45),
.C(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_46),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_54),
.C(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_11),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_7),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.C(n_7),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_8),
.Y(n_62)
);


endmodule