module fake_ibex_1650_n_4738 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4738);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4738;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_4688;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_4615;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4687;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_4632;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_3838;
wire n_957;
wire n_4514;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_4668;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_4731;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_4648;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_4601;
wire n_3340;
wire n_4142;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_3458;
wire n_2955;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4708;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_875;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_4652;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_4673;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_4690;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_4578;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_4447;
wire n_4491;
wire n_4672;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_4723;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4510;
wire n_4389;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_4312;
wire n_4567;
wire n_917;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_4214;
wire n_1313;
wire n_3973;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_4724;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_4721;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_4517;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_4735;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_4667;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_4711;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_4671;
wire n_971;
wire n_1326;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_4676;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_4714;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4732;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_3217;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_2401;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_4252;
wire n_1332;
wire n_2660;
wire n_4505;
wire n_3971;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_4692;
wire n_4713;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2646;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3963;
wire n_3887;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4126;
wire n_3583;
wire n_2019;
wire n_4103;
wire n_4710;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_4680;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_4693;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4549;
wire n_1441;
wire n_4105;
wire n_4090;
wire n_4573;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3320;
wire n_3117;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_4700;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4411;
wire n_1964;
wire n_4523;
wire n_4156;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_4712;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3634;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_4571;
wire n_959;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_4725;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4681;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_4374;
wire n_4501;
wire n_1985;
wire n_1140;
wire n_4375;
wire n_3815;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_4403;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4485;
wire n_4608;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1890;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_907;
wire n_1990;
wire n_1179;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_2999;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_4706;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2991;
wire n_2234;
wire n_2699;
wire n_847;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4674;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4679;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4456;
wire n_4215;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_3578;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_4734;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_4559;
wire n_1395;
wire n_998;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4660;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_4664;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_4709;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_4552;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1539;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_4683;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3718;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4291;
wire n_2781;
wire n_4035;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_4694;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_4717;
wire n_2507;
wire n_2759;
wire n_3682;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3434;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_4719;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_1967;
wire n_903;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4256;
wire n_1185;
wire n_1683;
wire n_4176;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_4685;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_4716;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_3284;
wire n_2524;
wire n_2875;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_4185;
wire n_2422;
wire n_3902;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_991;
wire n_1223;
wire n_961;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_4704;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4388;
wire n_4071;
wire n_4593;
wire n_996;
wire n_4247;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3673;
wire n_3476;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4123;
wire n_3154;
wire n_4000;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3696;
wire n_3113;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_4007;
wire n_3960;
wire n_3769;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_4707;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1962;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_4638;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_4319;
wire n_4637;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1923;
wire n_1224;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_4736;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_2194;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_4320;
wire n_2736;
wire n_4019;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_4697;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_4730;
wire n_1415;
wire n_1238;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_4720;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_4282;
wire n_4715;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3619;
wire n_3928;
wire n_3349;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_4698;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1989;
wire n_1740;
wire n_3649;
wire n_1838;
wire n_3540;
wire n_3604;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2576;
wire n_2675;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_4666;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_4663;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_4618;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4611;
wire n_897;
wire n_1622;
wire n_2757;
wire n_4148;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2816;
wire n_2803;
wire n_2433;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_4670;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2667;
wire n_2218;
wire n_4524;
wire n_3062;
wire n_4265;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2864;
wire n_2406;
wire n_1632;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1542;
wire n_1586;
wire n_1547;
wire n_946;
wire n_1362;
wire n_3497;
wire n_4696;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_3561;
wire n_956;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_4659;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2593;
wire n_3899;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_4729;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_4562;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_4345;
wire n_4281;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_4675;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_4737;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1572;
wire n_1635;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_3163;
wire n_2701;
wire n_2929;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1297;
wire n_1912;
wire n_1369;
wire n_3143;
wire n_1734;
wire n_3655;
wire n_3543;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_4686;
wire n_1529;
wire n_1824;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4682;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_4147;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_4218;
wire n_3898;
wire n_3366;
wire n_4705;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_4733;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_4684;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_2005;
wire n_1284;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_980;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3067;
wire n_1074;
wire n_3557;
wire n_3225;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_4657;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4718;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1904;
wire n_1262;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_4412;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3286;
wire n_999;
wire n_2634;
wire n_2982;
wire n_3124;
wire n_1092;
wire n_4038;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3398;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1516;
wire n_1027;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_2104;
wire n_2357;
wire n_2855;
wire n_2653;
wire n_2618;
wire n_3938;
wire n_4354;
wire n_924;
wire n_4448;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4532;
wire n_4401;
wire n_4727;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_4701;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_4726;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_4544;
wire n_4728;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_2066;
wire n_1158;
wire n_2988;
wire n_4275;
wire n_1882;
wire n_4046;
wire n_3945;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_2168;
wire n_1948;
wire n_3247;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_4689;
wire n_3613;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_4702;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_4506;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_856;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_4606;
wire n_1287;
wire n_2769;
wire n_3865;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3911;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_4703;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_4691;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_4662;
wire n_2658;

INVx2_ASAP7_75t_SL g845 ( 
.A(n_771),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_516),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_793),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_617),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_232),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_94),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_97),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_820),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_595),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_646),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_753),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_340),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_508),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_219),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_796),
.Y(n_859)
);

BUFx10_ASAP7_75t_L g860 ( 
.A(n_323),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_494),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_677),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_436),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_523),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_788),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_590),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_464),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_174),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_162),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_816),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_771),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_253),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_532),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_583),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_294),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_87),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_63),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_750),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_450),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_248),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_67),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_187),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_115),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_572),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_675),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_832),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_693),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_761),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_752),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_612),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_267),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_744),
.Y(n_892)
);

INVxp33_ASAP7_75t_L g893 ( 
.A(n_575),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_654),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_763),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_23),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_446),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_489),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_803),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_107),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_385),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_444),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_833),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_41),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_73),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_810),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_219),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_99),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_614),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_660),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_797),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_770),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_181),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_633),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_388),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_322),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_260),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_821),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_478),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_802),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_361),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_831),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_366),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_780),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_216),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_754),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_259),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_619),
.Y(n_928)
);

BUFx10_ASAP7_75t_L g929 ( 
.A(n_225),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_176),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_707),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_98),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_467),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_393),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_518),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_388),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_538),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_343),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_13),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_821),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_672),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_340),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_825),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_207),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_186),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_839),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_352),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_173),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_633),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_71),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_128),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_725),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_380),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_815),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_715),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_243),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_801),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_765),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_711),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_147),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_359),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_575),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_271),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_685),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_195),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_518),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_496),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_34),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_566),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_312),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_156),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_551),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_258),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_257),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_816),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_529),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_447),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_442),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_413),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_101),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_412),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_199),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_777),
.Y(n_983)
);

CKINVDCx14_ASAP7_75t_R g984 ( 
.A(n_126),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_576),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_183),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_178),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_210),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_35),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_393),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_496),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_783),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_593),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_702),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_664),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_824),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_823),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_337),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_776),
.Y(n_999)
);

BUFx2_ASAP7_75t_SL g1000 ( 
.A(n_762),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_479),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_438),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_448),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_231),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_329),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_585),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_687),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_552),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_213),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_783),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_392),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_682),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_732),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_745),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_499),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_416),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_212),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_174),
.Y(n_1018)
);

CKINVDCx14_ASAP7_75t_R g1019 ( 
.A(n_545),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_798),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_205),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_154),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_623),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_103),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_200),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_462),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_699),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_10),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_362),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_477),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_777),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_268),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_439),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_445),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_141),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_639),
.Y(n_1036)
);

CKINVDCx16_ASAP7_75t_R g1037 ( 
.A(n_283),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_540),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_642),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_192),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_792),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_385),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_20),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_335),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_350),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_672),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_789),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_179),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_789),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_192),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_640),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_769),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_634),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_730),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_45),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_12),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_132),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_711),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_774),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_749),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_565),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_146),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_521),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_449),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_360),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_828),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_786),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_706),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_309),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_143),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_194),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_392),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_37),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_729),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_91),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_321),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_656),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_602),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_230),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_176),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_839),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_586),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_627),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_641),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_801),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_457),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_645),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_763),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_786),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_809),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_500),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_61),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_600),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_618),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_726),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_744),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_493),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_617),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_81),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_790),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_508),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_697),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_594),
.Y(n_1103)
);

CKINVDCx16_ASAP7_75t_R g1104 ( 
.A(n_131),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_56),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_301),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_34),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_619),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_58),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_810),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_818),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_288),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_811),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_813),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_772),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_35),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_755),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_817),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_206),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_297),
.Y(n_1120)
);

BUFx2_ASAP7_75t_SL g1121 ( 
.A(n_545),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_685),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_807),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_85),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_192),
.Y(n_1125)
);

CKINVDCx16_ASAP7_75t_R g1126 ( 
.A(n_599),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_494),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_0),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_768),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_668),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_177),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_799),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_745),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_781),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_211),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_766),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_353),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_665),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_719),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_784),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_59),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_806),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_203),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_600),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_173),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_91),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_245),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_616),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_357),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_372),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_661),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_272),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_782),
.Y(n_1153)
);

CKINVDCx6p67_ASAP7_75t_R g1154 ( 
.A(n_145),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_653),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_111),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_645),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_235),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_207),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_62),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_77),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_215),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_830),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_794),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_88),
.Y(n_1165)
);

CKINVDCx16_ASAP7_75t_R g1166 ( 
.A(n_373),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_484),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_694),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_332),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_661),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_130),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_774),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_803),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_313),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_264),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_727),
.Y(n_1176)
);

BUFx8_ASAP7_75t_SL g1177 ( 
.A(n_693),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_125),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_383),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_246),
.Y(n_1180)
);

BUFx2_ASAP7_75t_SL g1181 ( 
.A(n_730),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_245),
.Y(n_1182)
);

CKINVDCx14_ASAP7_75t_R g1183 ( 
.A(n_181),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_606),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_210),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_488),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_674),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_161),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_787),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_663),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_581),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_45),
.Y(n_1192)
);

BUFx2_ASAP7_75t_SL g1193 ( 
.A(n_128),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_236),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_75),
.Y(n_1195)
);

CKINVDCx14_ASAP7_75t_R g1196 ( 
.A(n_607),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_228),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_499),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_107),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_800),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_421),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_696),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_464),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_111),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_280),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_361),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_713),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_417),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_62),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_197),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_787),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_43),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_332),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_775),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_234),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_131),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_764),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_307),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_369),
.Y(n_1219)
);

INVxp33_ASAP7_75t_SL g1220 ( 
.A(n_701),
.Y(n_1220)
);

BUFx5_ASAP7_75t_L g1221 ( 
.A(n_469),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_581),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_370),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_28),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_321),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_374),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_805),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_570),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_460),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_565),
.Y(n_1230)
);

BUFx5_ASAP7_75t_L g1231 ( 
.A(n_808),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_220),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_211),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_156),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_330),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_750),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_237),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_832),
.Y(n_1238)
);

CKINVDCx16_ASAP7_75t_R g1239 ( 
.A(n_467),
.Y(n_1239)
);

BUFx5_ASAP7_75t_L g1240 ( 
.A(n_282),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_691),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_224),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_236),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_530),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_354),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_631),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_428),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_552),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_520),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_221),
.Y(n_1250)
);

CKINVDCx16_ASAP7_75t_R g1251 ( 
.A(n_574),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_778),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_132),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_110),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_624),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_708),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_770),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_121),
.Y(n_1258)
);

CKINVDCx14_ASAP7_75t_R g1259 ( 
.A(n_656),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_430),
.Y(n_1260)
);

BUFx5_ASAP7_75t_L g1261 ( 
.A(n_30),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_471),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_799),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_829),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_260),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_716),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_428),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_127),
.Y(n_1268)
);

CKINVDCx14_ASAP7_75t_R g1269 ( 
.A(n_549),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_757),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_764),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_317),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_815),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_747),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_68),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_785),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_694),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_122),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_773),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_776),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_714),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_292),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_316),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_812),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_254),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_257),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_188),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_58),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_618),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_827),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_791),
.Y(n_1291)
);

CKINVDCx14_ASAP7_75t_R g1292 ( 
.A(n_311),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_779),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_31),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_736),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_715),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_301),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_682),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_439),
.Y(n_1299)
);

BUFx10_ASAP7_75t_L g1300 ( 
.A(n_521),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_28),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_403),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_369),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_215),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_731),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_394),
.Y(n_1306)
);

BUFx10_ASAP7_75t_L g1307 ( 
.A(n_104),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_187),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_62),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_729),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_698),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_606),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_804),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_163),
.Y(n_1314)
);

CKINVDCx14_ASAP7_75t_R g1315 ( 
.A(n_32),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_419),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_607),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_826),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_628),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_597),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_19),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_455),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_580),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_490),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_354),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_822),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_43),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_408),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_252),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_649),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_70),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_814),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_252),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_38),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_602),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_670),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_709),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_418),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_577),
.Y(n_1339)
);

CKINVDCx14_ASAP7_75t_R g1340 ( 
.A(n_323),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_403),
.Y(n_1341)
);

BUFx8_ASAP7_75t_SL g1342 ( 
.A(n_96),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_844),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_242),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_402),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_781),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_182),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_328),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_41),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_819),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_266),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_239),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_775),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_320),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_497),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_27),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_207),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_446),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_326),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_611),
.Y(n_1360)
);

BUFx10_ASAP7_75t_L g1361 ( 
.A(n_180),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_622),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_835),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_364),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_114),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_512),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_767),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_515),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_758),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_795),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_328),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_313),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_188),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_60),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_216),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_279),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_469),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_800),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_167),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_465),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_700),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1232),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1232),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_984),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1232),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1175),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1342),
.Y(n_1387)
);

INVxp67_ASAP7_75t_SL g1388 ( 
.A(n_1032),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1185),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1183),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1242),
.Y(n_1391)
);

INVxp33_ASAP7_75t_SL g1392 ( 
.A(n_904),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1342),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1315),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_929),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1265),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1352),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1301),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1160),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1160),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1216),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1216),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1294),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_875),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1294),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1154),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_845),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_845),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1154),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1177),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1177),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_970),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_970),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_990),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_917),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_893),
.B(n_0),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_896),
.Y(n_1417)
);

CKINVDCx16_ASAP7_75t_R g1418 ( 
.A(n_1028),
.Y(n_1418)
);

INVxp33_ASAP7_75t_SL g1419 ( 
.A(n_1031),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1032),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_875),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_896),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_877),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_990),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_905),
.Y(n_1425)
);

INVxp33_ASAP7_75t_SL g1426 ( 
.A(n_905),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_907),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_877),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1050),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1098),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_882),
.Y(n_1431)
);

NOR2xp67_ASAP7_75t_L g1432 ( 
.A(n_1098),
.B(n_0),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1311),
.Y(n_1433)
);

INVxp67_ASAP7_75t_SL g1434 ( 
.A(n_1050),
.Y(n_1434)
);

XNOR2x1_ASAP7_75t_L g1435 ( 
.A(n_907),
.B(n_1),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_955),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1311),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_882),
.Y(n_1438)
);

NAND2xp33_ASAP7_75t_R g1439 ( 
.A(n_977),
.B(n_1),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1081),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1037),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1176),
.B(n_1),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1104),
.B(n_2),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1105),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1312),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1312),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_908),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1245),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1313),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_908),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1329),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_850),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1329),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1334),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_858),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_869),
.Y(n_1456)
);

CKINVDCx16_ASAP7_75t_R g1457 ( 
.A(n_929),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_876),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1316),
.B(n_2),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1366),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1334),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_913),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1019),
.Y(n_1463)
);

INVxp33_ASAP7_75t_SL g1464 ( 
.A(n_851),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_913),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_883),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_927),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1196),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_1105),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_932),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_963),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_927),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1259),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1269),
.Y(n_1474)
);

NOR2xp67_ASAP7_75t_L g1475 ( 
.A(n_1322),
.B(n_2),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_965),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_1292),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1240),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_973),
.B(n_3),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_974),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_982),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_986),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_900),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1340),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_987),
.Y(n_1485)
);

CKINVDCx16_ASAP7_75t_R g1486 ( 
.A(n_929),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_900),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_988),
.Y(n_1488)
);

CKINVDCx16_ASAP7_75t_R g1489 ( 
.A(n_989),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_868),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_872),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1009),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1021),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1024),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1240),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1025),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_968),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_880),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_881),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_891),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1073),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_925),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1109),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_968),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1240),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_930),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1112),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1079),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1120),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1420),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1399),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1426),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1457),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1486),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1386),
.B(n_1091),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1398),
.B(n_989),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1400),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1401),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1451),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1420),
.Y(n_1520)
);

INVxp33_ASAP7_75t_L g1521 ( 
.A(n_1450),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1382),
.Y(n_1522)
);

BUFx2_ASAP7_75t_L g1523 ( 
.A(n_1422),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_SL g1524 ( 
.A(n_1389),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_1467),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1383),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1489),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1425),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1427),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1395),
.Y(n_1530)
);

INVx6_ASAP7_75t_L g1531 ( 
.A(n_1418),
.Y(n_1531)
);

AND2x6_ASAP7_75t_L g1532 ( 
.A(n_1395),
.B(n_1091),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1402),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1467),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1403),
.Y(n_1535)
);

AND2x6_ASAP7_75t_L g1536 ( 
.A(n_1417),
.B(n_1093),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1478),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1508),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1405),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1388),
.B(n_944),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1429),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1447),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1434),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1453),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1391),
.B(n_1093),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1468),
.B(n_1220),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1454),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1461),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1444),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1393),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1469),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1464),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1407),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1408),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1478),
.A2(n_1161),
.B(n_939),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1412),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1415),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1508),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1385),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1404),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1413),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1421),
.A2(n_1428),
.B1(n_1431),
.B2(n_1423),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1415),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1414),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1490),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1441),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1392),
.B(n_945),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1441),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1424),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1406),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1438),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1430),
.Y(n_1572)
);

CKINVDCx16_ASAP7_75t_R g1573 ( 
.A(n_1384),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1409),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1433),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1387),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1437),
.B(n_1220),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1491),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1396),
.B(n_1095),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1495),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1495),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1505),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1445),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1446),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_L g1585 ( 
.A(n_1452),
.B(n_1240),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1462),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1449),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1505),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1397),
.B(n_1095),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1483),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1487),
.Y(n_1591)
);

CKINVDCx16_ASAP7_75t_R g1592 ( 
.A(n_1384),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1455),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1456),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1498),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1436),
.B(n_948),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1458),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1466),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1440),
.B(n_950),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1470),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1471),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1465),
.Y(n_1602)
);

NOR2xp33_ASAP7_75t_R g1603 ( 
.A(n_1390),
.B(n_1126),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1476),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1480),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1472),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1499),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1481),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1482),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1459),
.Y(n_1610)
);

AND2x2_ASAP7_75t_SL g1611 ( 
.A(n_1416),
.B(n_1166),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1500),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1502),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1506),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1448),
.B(n_1460),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1485),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1488),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1492),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1463),
.B(n_1239),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1497),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1493),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1494),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1473),
.B(n_1240),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1410),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1496),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1501),
.Y(n_1626)
);

CKINVDCx6p67_ASAP7_75t_R g1627 ( 
.A(n_1390),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1503),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1507),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1509),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1411),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1416),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1394),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1419),
.B(n_951),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1435),
.Y(n_1635)
);

CKINVDCx16_ASAP7_75t_R g1636 ( 
.A(n_1394),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1475),
.B(n_853),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1432),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1442),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1479),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1442),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1443),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1474),
.B(n_1477),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1504),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1435),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1484),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1439),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1439),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1426),
.Y(n_1649)
);

INVx4_ASAP7_75t_L g1650 ( 
.A(n_1395),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1451),
.B(n_1000),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1399),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1420),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1426),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1426),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1399),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1426),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1399),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1386),
.B(n_853),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1426),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1420),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1395),
.B(n_956),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1467),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1426),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1426),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1420),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1420),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1467),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1426),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1420),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1426),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1399),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1386),
.B(n_861),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1399),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1426),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1420),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1395),
.B(n_1251),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1422),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1420),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1420),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1399),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1422),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1426),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1395),
.B(n_960),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1399),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1426),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1439),
.A2(n_1119),
.B1(n_1125),
.B2(n_1079),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1422),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1382),
.A2(n_1161),
.B(n_939),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1420),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1399),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_1426),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1426),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1426),
.Y(n_1694)
);

XNOR2x2_ASAP7_75t_R g1695 ( 
.A(n_1387),
.B(n_3),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1426),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1395),
.B(n_971),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1399),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_1467),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1399),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_SL g1701 ( 
.A(n_1457),
.B(n_989),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1426),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1426),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1420),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1399),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1426),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1467),
.A2(n_1125),
.B1(n_1178),
.B2(n_1119),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1399),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1399),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1395),
.B(n_980),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1420),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1426),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1399),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1426),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1399),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1451),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1420),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1420),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1451),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1399),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1426),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1426),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1516),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1519),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1621),
.B(n_1070),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1554),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1689),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1555),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1520),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1615),
.B(n_895),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1521),
.B(n_1070),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1642),
.A2(n_1375),
.B1(n_1373),
.B2(n_1018),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1554),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1556),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1555),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1650),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1520),
.Y(n_1737)
);

AND2x6_ASAP7_75t_L g1738 ( 
.A(n_1648),
.B(n_1288),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1513),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1530),
.B(n_1004),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1641),
.A2(n_1128),
.B1(n_1147),
.B2(n_1145),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1520),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1556),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1632),
.B(n_1070),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1531),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1610),
.B(n_1240),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1625),
.Y(n_1747)
);

CKINVDCx20_ASAP7_75t_R g1748 ( 
.A(n_1560),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1530),
.B(n_1017),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1632),
.B(n_1307),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1639),
.A2(n_1156),
.B1(n_1159),
.B2(n_1152),
.Y(n_1751)
);

NAND2xp33_ASAP7_75t_SL g1752 ( 
.A(n_1647),
.B(n_1022),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1625),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1651),
.B(n_848),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1651),
.B(n_852),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1651),
.B(n_854),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1540),
.B(n_1240),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1650),
.B(n_1035),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

BUFx4_ASAP7_75t_L g1760 ( 
.A(n_1695),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1531),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1716),
.B(n_897),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1523),
.B(n_1121),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1511),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1639),
.A2(n_1180),
.B1(n_1194),
.B2(n_1171),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1515),
.B(n_855),
.Y(n_1766)
);

NAND2x1p5_ASAP7_75t_L g1767 ( 
.A(n_1529),
.B(n_849),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1661),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1541),
.B(n_1261),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1543),
.B(n_1261),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1639),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1517),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1632),
.B(n_1307),
.Y(n_1773)
);

AND2x6_ASAP7_75t_L g1774 ( 
.A(n_1549),
.B(n_1288),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1661),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1719),
.B(n_1307),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1567),
.B(n_897),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1701),
.B(n_1361),
.Y(n_1778)
);

NOR2x1p5_ASAP7_75t_L g1779 ( 
.A(n_1514),
.B(n_898),
.Y(n_1779)
);

BUFx10_ASAP7_75t_L g1780 ( 
.A(n_1524),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1611),
.A2(n_1043),
.B1(n_1048),
.B2(n_1040),
.Y(n_1781)
);

BUFx2_ASAP7_75t_L g1782 ( 
.A(n_1678),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1682),
.B(n_1361),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1532),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1661),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1527),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1518),
.Y(n_1787)
);

BUFx10_ASAP7_75t_L g1788 ( 
.A(n_1524),
.Y(n_1788)
);

INVx5_ASAP7_75t_L g1789 ( 
.A(n_1532),
.Y(n_1789)
);

AND2x6_ASAP7_75t_L g1790 ( 
.A(n_1551),
.B(n_1116),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1667),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1532),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1667),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1688),
.B(n_1634),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1578),
.B(n_1614),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1667),
.Y(n_1796)
);

INVx5_ASAP7_75t_L g1797 ( 
.A(n_1532),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1680),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1659),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1565),
.B(n_1361),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1533),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1680),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1659),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1535),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1662),
.B(n_1055),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1590),
.B(n_1261),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1673),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1539),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1680),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1684),
.B(n_1056),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1515),
.B(n_865),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1652),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1656),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1591),
.B(n_1261),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1697),
.B(n_1057),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1711),
.Y(n_1816)
);

BUFx10_ASAP7_75t_L g1817 ( 
.A(n_1552),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1711),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1710),
.B(n_1062),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1658),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1711),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_SL g1822 ( 
.A1(n_1707),
.A2(n_1254),
.B1(n_1275),
.B2(n_1178),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1594),
.B(n_1261),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1672),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1674),
.Y(n_1825)
);

CKINVDCx20_ASAP7_75t_R g1826 ( 
.A(n_1571),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1681),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1545),
.B(n_871),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1685),
.Y(n_1829)
);

BUFx10_ASAP7_75t_L g1830 ( 
.A(n_1512),
.Y(n_1830)
);

INVx4_ASAP7_75t_L g1831 ( 
.A(n_1718),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1691),
.Y(n_1832)
);

INVx4_ASAP7_75t_L g1833 ( 
.A(n_1718),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1586),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1718),
.Y(n_1835)
);

AND2x6_ASAP7_75t_L g1836 ( 
.A(n_1638),
.B(n_1116),
.Y(n_1836)
);

AND2x6_ASAP7_75t_L g1837 ( 
.A(n_1640),
.B(n_1116),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_SL g1838 ( 
.A(n_1595),
.B(n_1254),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1510),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1597),
.B(n_1071),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1598),
.B(n_1261),
.Y(n_1841)
);

AND2x6_ASAP7_75t_L g1842 ( 
.A(n_1643),
.B(n_1116),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1653),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1649),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1596),
.B(n_1075),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1545),
.B(n_878),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1698),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1599),
.B(n_1080),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1666),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1677),
.A2(n_1099),
.B1(n_1106),
.B2(n_1092),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1700),
.Y(n_1851)
);

CKINVDCx20_ASAP7_75t_R g1852 ( 
.A(n_1602),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_1536),
.Y(n_1853)
);

BUFx10_ASAP7_75t_L g1854 ( 
.A(n_1654),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1670),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1601),
.B(n_1604),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1655),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1676),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1579),
.B(n_886),
.Y(n_1859)
);

AND2x6_ASAP7_75t_L g1860 ( 
.A(n_1646),
.B(n_1124),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1536),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1605),
.B(n_1107),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1679),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1609),
.B(n_1261),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1690),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1546),
.B(n_1131),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1577),
.A2(n_1141),
.B1(n_1143),
.B2(n_1135),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1705),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1657),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1708),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1660),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1537),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1616),
.B(n_1146),
.Y(n_1873)
);

INVx5_ASAP7_75t_L g1874 ( 
.A(n_1537),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1622),
.B(n_1626),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1606),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_SL g1877 ( 
.A(n_1607),
.B(n_1275),
.Y(n_1877)
);

INVx5_ASAP7_75t_L g1878 ( 
.A(n_1537),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1709),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1717),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1579),
.B(n_889),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1582),
.Y(n_1882)
);

AND2x6_ASAP7_75t_L g1883 ( 
.A(n_1628),
.B(n_1124),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1713),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1687),
.B(n_898),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1522),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1715),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1620),
.Y(n_1888)
);

AO21x2_ASAP7_75t_L g1889 ( 
.A1(n_1585),
.A2(n_1199),
.B(n_1195),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1664),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1548),
.A2(n_1162),
.B1(n_1165),
.B2(n_1158),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1665),
.Y(n_1892)
);

INVx4_ASAP7_75t_L g1893 ( 
.A(n_1536),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1644),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1629),
.B(n_1182),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1720),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1630),
.B(n_1188),
.Y(n_1897)
);

BUFx10_ASAP7_75t_L g1898 ( 
.A(n_1669),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1553),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1561),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1564),
.Y(n_1901)
);

INVx6_ASAP7_75t_L g1902 ( 
.A(n_1673),
.Y(n_1902)
);

AND2x6_ASAP7_75t_L g1903 ( 
.A(n_1569),
.B(n_1124),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1593),
.B(n_1197),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1526),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_SL g1906 ( 
.A(n_1612),
.B(n_1331),
.Y(n_1906)
);

INVx4_ASAP7_75t_L g1907 ( 
.A(n_1536),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1559),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1589),
.B(n_890),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1572),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1582),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1575),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1671),
.Y(n_1913)
);

INVx2_ASAP7_75t_SL g1914 ( 
.A(n_1675),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1687),
.B(n_901),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1683),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1583),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1600),
.B(n_1205),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1686),
.B(n_901),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1692),
.B(n_860),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1589),
.B(n_1209),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1584),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1608),
.B(n_1210),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1693),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1637),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1637),
.B(n_892),
.Y(n_1926)
);

OR2x6_ASAP7_75t_L g1927 ( 
.A(n_1562),
.B(n_1181),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1694),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1617),
.B(n_1212),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1587),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1557),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1582),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1696),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1623),
.B(n_1233),
.Y(n_1934)
);

HB1xp67_ASAP7_75t_L g1935 ( 
.A(n_1702),
.Y(n_1935)
);

INVx5_ASAP7_75t_L g1936 ( 
.A(n_1588),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1618),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1588),
.B(n_1234),
.Y(n_1938)
);

BUFx3_ASAP7_75t_L g1939 ( 
.A(n_1703),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1580),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1581),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1528),
.A2(n_1258),
.B1(n_1268),
.B2(n_1243),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1706),
.Y(n_1943)
);

BUFx3_ASAP7_75t_L g1944 ( 
.A(n_1712),
.Y(n_1944)
);

OAI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1714),
.A2(n_1722),
.B1(n_1721),
.B2(n_1645),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1542),
.B(n_1547),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1544),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1613),
.Y(n_1948)
);

INVx2_ASAP7_75t_SL g1949 ( 
.A(n_1603),
.Y(n_1949)
);

INVx4_ASAP7_75t_L g1950 ( 
.A(n_1570),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1619),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1574),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1635),
.B(n_860),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_L g1954 ( 
.A(n_1550),
.B(n_1221),
.Y(n_1954)
);

INVx5_ASAP7_75t_L g1955 ( 
.A(n_1573),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1624),
.Y(n_1956)
);

BUFx6f_ASAP7_75t_L g1957 ( 
.A(n_1631),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1627),
.B(n_860),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1563),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1592),
.B(n_1282),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1566),
.B(n_1287),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1568),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1633),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1636),
.B(n_1001),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1525),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1576),
.Y(n_1966)
);

INVx5_ASAP7_75t_L g1967 ( 
.A(n_1534),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1538),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1558),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1699),
.B(n_1001),
.Y(n_1970)
);

INVx4_ASAP7_75t_SL g1971 ( 
.A(n_1663),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1668),
.B(n_902),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1689),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1554),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1516),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1610),
.B(n_1304),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_SL g1977 ( 
.A1(n_1525),
.A2(n_1365),
.B1(n_1331),
.B2(n_857),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1521),
.B(n_1001),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1610),
.B(n_1314),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1641),
.A2(n_1204),
.B1(n_1237),
.B2(n_1215),
.Y(n_1980)
);

NAND2xp33_ASAP7_75t_L g1981 ( 
.A(n_1532),
.B(n_1221),
.Y(n_1981)
);

AO21x2_ASAP7_75t_L g1982 ( 
.A1(n_1689),
.A2(n_1253),
.B(n_1250),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1530),
.B(n_1321),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1531),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1554),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1554),
.Y(n_1986)
);

NAND2xp33_ASAP7_75t_L g1987 ( 
.A(n_1532),
.B(n_1221),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1621),
.B(n_1344),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1615),
.B(n_902),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1689),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_1531),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1516),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1610),
.B(n_1347),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1554),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1610),
.B(n_1349),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1621),
.B(n_1351),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1554),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1554),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1554),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1554),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1521),
.B(n_1163),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1555),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1689),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1554),
.Y(n_2004)
);

INVx4_ASAP7_75t_L g2005 ( 
.A(n_1532),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1554),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1689),
.Y(n_2007)
);

INVx1_ASAP7_75t_SL g2008 ( 
.A(n_1519),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1689),
.Y(n_2009)
);

BUFx6f_ASAP7_75t_L g2010 ( 
.A(n_1555),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1555),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1689),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1736),
.Y(n_2013)
);

NAND3xp33_ASAP7_75t_SL g2014 ( 
.A(n_1871),
.B(n_1371),
.C(n_857),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1723),
.B(n_894),
.Y(n_2015)
);

NAND2x1p5_ASAP7_75t_L g2016 ( 
.A(n_1724),
.B(n_1224),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1764),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1784),
.B(n_1356),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1976),
.B(n_1357),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1979),
.B(n_1278),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1937),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1993),
.B(n_909),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1995),
.B(n_909),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1784),
.B(n_912),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1772),
.Y(n_2025)
);

NOR3xp33_ASAP7_75t_SL g2026 ( 
.A(n_1739),
.B(n_1786),
.C(n_1931),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1767),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1845),
.B(n_912),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1792),
.B(n_2005),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1782),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1848),
.B(n_914),
.Y(n_2031)
);

O2A1O1Ixp33_ASAP7_75t_L g2032 ( 
.A1(n_1730),
.A2(n_1286),
.B(n_1297),
.C(n_1285),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1787),
.Y(n_2033)
);

O2A1O1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1989),
.A2(n_1885),
.B(n_1915),
.C(n_1961),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1745),
.Y(n_2035)
);

NAND2x1_ASAP7_75t_L g2036 ( 
.A(n_1792),
.B(n_1124),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1805),
.B(n_1328),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_1774),
.A2(n_1308),
.B1(n_1327),
.B2(n_1309),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1810),
.B(n_1328),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1819),
.B(n_1332),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1774),
.B(n_1332),
.Y(n_2041)
);

NOR3xp33_ASAP7_75t_L g2042 ( 
.A(n_1945),
.B(n_1082),
.C(n_1045),
.Y(n_2042)
);

NOR2xp33_ASAP7_75t_L g2043 ( 
.A(n_1951),
.B(n_1335),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1774),
.B(n_1335),
.Y(n_2044)
);

INVxp67_ASAP7_75t_L g2045 ( 
.A(n_2008),
.Y(n_2045)
);

A2O1A1Ixp33_ASAP7_75t_L g2046 ( 
.A1(n_1801),
.A2(n_1374),
.B(n_1379),
.C(n_1333),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1731),
.B(n_1336),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1758),
.B(n_1336),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_2005),
.B(n_1337),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1804),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1875),
.B(n_1337),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1895),
.B(n_1338),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1728),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1897),
.B(n_1338),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1732),
.B(n_1341),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1808),
.B(n_1341),
.Y(n_2056)
);

AND2x6_ASAP7_75t_SL g2057 ( 
.A(n_1927),
.B(n_1371),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1975),
.B(n_856),
.Y(n_2058)
);

NAND2xp33_ASAP7_75t_L g2059 ( 
.A(n_1789),
.B(n_1231),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1937),
.Y(n_2060)
);

AOI22xp33_ASAP7_75t_L g2061 ( 
.A1(n_1738),
.A2(n_1193),
.B1(n_1376),
.B2(n_1192),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1812),
.B(n_846),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1789),
.B(n_847),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1771),
.A2(n_863),
.B1(n_918),
.B2(n_856),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1789),
.B(n_859),
.Y(n_2065)
);

A2O1A1Ixp33_ASAP7_75t_L g2066 ( 
.A1(n_1813),
.A2(n_906),
.B(n_910),
.C(n_899),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1782),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1820),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1937),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1728),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1824),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_1831),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1825),
.B(n_864),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1827),
.B(n_867),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1834),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1829),
.B(n_870),
.Y(n_2076)
);

INVx5_ASAP7_75t_L g2077 ( 
.A(n_1790),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1992),
.B(n_863),
.Y(n_2078)
);

AOI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1738),
.A2(n_947),
.B1(n_953),
.B2(n_918),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1832),
.B(n_873),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1847),
.Y(n_2081)
);

INVx2_ASAP7_75t_SL g2082 ( 
.A(n_1984),
.Y(n_2082)
);

A2O1A1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_1851),
.A2(n_915),
.B(n_916),
.C(n_911),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1794),
.B(n_947),
.Y(n_2084)
);

INVx2_ASAP7_75t_SL g2085 ( 
.A(n_1991),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1797),
.B(n_874),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1738),
.A2(n_964),
.B1(n_972),
.B2(n_953),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1776),
.B(n_964),
.Y(n_2088)
);

AND2x6_ASAP7_75t_SL g2089 ( 
.A(n_1927),
.B(n_972),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1940),
.Y(n_2090)
);

INVxp67_ASAP7_75t_L g2091 ( 
.A(n_1838),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1868),
.B(n_879),
.Y(n_2092)
);

A2O1A1Ixp33_ASAP7_75t_L g2093 ( 
.A1(n_1870),
.A2(n_926),
.B(n_934),
.C(n_921),
.Y(n_2093)
);

OAI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_1751),
.A2(n_1011),
.B1(n_1046),
.B2(n_976),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1940),
.Y(n_2095)
);

NAND2x1_ASAP7_75t_L g2096 ( 
.A(n_1790),
.B(n_1192),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1879),
.B(n_1884),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1940),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1887),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1777),
.B(n_1919),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1797),
.B(n_884),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1896),
.B(n_885),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_1740),
.A2(n_1376),
.B1(n_1192),
.B2(n_1011),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1899),
.B(n_887),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1726),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1900),
.B(n_888),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_1762),
.B(n_976),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1901),
.B(n_1910),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1797),
.B(n_919),
.Y(n_2109)
);

INVx2_ASAP7_75t_SL g2110 ( 
.A(n_1780),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_1727),
.A2(n_946),
.B(n_938),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1795),
.B(n_920),
.Y(n_2112)
);

AOI22xp33_ASAP7_75t_L g2113 ( 
.A1(n_1866),
.A2(n_1765),
.B1(n_1754),
.B2(n_1756),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1912),
.B(n_923),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1783),
.B(n_1046),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1733),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1917),
.B(n_924),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1922),
.B(n_928),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1930),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1850),
.B(n_931),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1800),
.B(n_1087),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1734),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1953),
.B(n_1087),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_SL g2124 ( 
.A1(n_1822),
.A2(n_1172),
.B1(n_1186),
.B2(n_1090),
.Y(n_2124)
);

O2A1O1Ixp5_ASAP7_75t_L g2125 ( 
.A1(n_1744),
.A2(n_1750),
.B(n_1773),
.C(n_1815),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1743),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1749),
.B(n_933),
.Y(n_2127)
);

AO22x1_ASAP7_75t_L g2128 ( 
.A1(n_1967),
.A2(n_1172),
.B1(n_1186),
.B2(n_1090),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_1978),
.B(n_1214),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_1972),
.B(n_1208),
.Y(n_2130)
);

AND2x2_ASAP7_75t_SL g2131 ( 
.A(n_1877),
.B(n_1214),
.Y(n_2131)
);

INVx2_ASAP7_75t_SL g2132 ( 
.A(n_1780),
.Y(n_2132)
);

AOI22xp33_ASAP7_75t_SL g2133 ( 
.A1(n_1906),
.A2(n_1226),
.B1(n_1238),
.B2(n_1228),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_1844),
.B(n_1213),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1886),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1983),
.B(n_935),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1754),
.B(n_937),
.Y(n_2137)
);

NAND2x1_ASAP7_75t_L g2138 ( 
.A(n_1790),
.B(n_1192),
.Y(n_2138)
);

AO22x1_ASAP7_75t_L g2139 ( 
.A1(n_1967),
.A2(n_1228),
.B1(n_1238),
.B2(n_1226),
.Y(n_2139)
);

A2O1A1Ixp33_ASAP7_75t_L g2140 ( 
.A1(n_1757),
.A2(n_959),
.B(n_978),
.C(n_958),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1905),
.Y(n_2141)
);

OAI221xp5_ASAP7_75t_L g2142 ( 
.A1(n_1781),
.A2(n_1350),
.B1(n_942),
.B2(n_949),
.C(n_941),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1904),
.B(n_940),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2001),
.B(n_1263),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1856),
.A2(n_1296),
.B1(n_1310),
.B2(n_1263),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1755),
.B(n_952),
.Y(n_2146)
);

INVx8_ASAP7_75t_L g2147 ( 
.A(n_1842),
.Y(n_2147)
);

BUFx3_ASAP7_75t_L g2148 ( 
.A(n_1761),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1755),
.B(n_954),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1908),
.Y(n_2150)
);

NAND2x1p5_ASAP7_75t_L g2151 ( 
.A(n_1950),
.B(n_1376),
.Y(n_2151)
);

BUFx2_ASAP7_75t_L g2152 ( 
.A(n_1844),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1974),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1756),
.B(n_957),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1985),
.Y(n_2155)
);

NOR3xp33_ASAP7_75t_L g2156 ( 
.A(n_1960),
.B(n_966),
.C(n_962),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_SL g2157 ( 
.A(n_1950),
.B(n_1296),
.Y(n_2157)
);

NAND3xp33_ASAP7_75t_L g2158 ( 
.A(n_1942),
.B(n_969),
.C(n_967),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1918),
.B(n_979),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1923),
.B(n_981),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1861),
.B(n_983),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1929),
.B(n_985),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1861),
.B(n_993),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1725),
.B(n_991),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1746),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1986),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1741),
.B(n_994),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_L g2168 ( 
.A(n_2002),
.B(n_1221),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_1766),
.A2(n_1376),
.B1(n_1339),
.B2(n_1362),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1857),
.B(n_1310),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1806),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_1766),
.A2(n_1362),
.B1(n_1339),
.B2(n_999),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_L g2173 ( 
.A(n_1920),
.B(n_995),
.Y(n_2173)
);

AND2x2_ASAP7_75t_SL g2174 ( 
.A(n_1857),
.B(n_861),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1814),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1769),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1994),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1980),
.B(n_996),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1893),
.B(n_1907),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1770),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1921),
.B(n_997),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1867),
.B(n_1811),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1811),
.B(n_998),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1925),
.Y(n_2184)
);

AND2x6_ASAP7_75t_L g2185 ( 
.A(n_1853),
.B(n_862),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1893),
.B(n_1002),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_1907),
.B(n_1003),
.Y(n_2187)
);

BUFx8_ASAP7_75t_L g2188 ( 
.A(n_1924),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1828),
.B(n_1006),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_1988),
.B(n_992),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1747),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1828),
.B(n_1007),
.Y(n_2192)
);

AOI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_1891),
.A2(n_1010),
.B1(n_1015),
.B2(n_1012),
.C(n_1005),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1997),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1928),
.B(n_1892),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1846),
.B(n_1859),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1998),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1943),
.B(n_1008),
.Y(n_2198)
);

AOI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_1753),
.A2(n_1231),
.B1(n_1221),
.B2(n_1042),
.Y(n_2199)
);

INVx4_ASAP7_75t_L g2200 ( 
.A(n_1788),
.Y(n_2200)
);

OAI22xp33_ASAP7_75t_L g2201 ( 
.A1(n_1928),
.A2(n_1369),
.B1(n_1378),
.B2(n_1368),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1902),
.B(n_1013),
.Y(n_2202)
);

AND3x1_ASAP7_75t_L g2203 ( 
.A(n_1760),
.B(n_1049),
.C(n_1020),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1876),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_SL g2205 ( 
.A(n_1853),
.B(n_1014),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1902),
.B(n_1016),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1799),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_2002),
.Y(n_2208)
);

BUFx5_ASAP7_75t_L g2209 ( 
.A(n_1883),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_1936),
.B(n_1934),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1803),
.Y(n_2211)
);

AOI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1999),
.A2(n_1231),
.B1(n_1221),
.B2(n_1052),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_1962),
.B(n_1023),
.Y(n_2213)
);

AOI22xp33_ASAP7_75t_L g2214 ( 
.A1(n_1846),
.A2(n_1053),
.B1(n_1058),
.B2(n_1051),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_2010),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_1936),
.B(n_1752),
.Y(n_2216)
);

INVx2_ASAP7_75t_SL g2217 ( 
.A(n_1788),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1807),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_1955),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2000),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1859),
.B(n_1026),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_1913),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2004),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1881),
.B(n_1027),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1881),
.B(n_1029),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2006),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_1947),
.B(n_1030),
.Y(n_2227)
);

NAND2x1p5_ASAP7_75t_L g2228 ( 
.A(n_1916),
.B(n_1059),
.Y(n_2228)
);

OAI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_2010),
.A2(n_1069),
.B1(n_1108),
.B2(n_1066),
.Y(n_2229)
);

AND2x2_ASAP7_75t_SL g2230 ( 
.A(n_1935),
.B(n_862),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1909),
.B(n_1033),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1936),
.B(n_1034),
.Y(n_2232)
);

OR2x6_ASAP7_75t_L g2233 ( 
.A(n_1763),
.B(n_903),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1909),
.B(n_1038),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1982),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1938),
.B(n_1041),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1926),
.B(n_1044),
.Y(n_2237)
);

INVx2_ASAP7_75t_SL g2238 ( 
.A(n_1955),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_1977),
.B(n_1047),
.Y(n_2239)
);

AND2x2_ASAP7_75t_SL g2240 ( 
.A(n_1760),
.B(n_903),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_1941),
.A2(n_1231),
.B1(n_1221),
.B2(n_1115),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1926),
.B(n_1054),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1735),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_1973),
.A2(n_1117),
.B(n_1110),
.Y(n_2244)
);

INVxp67_ASAP7_75t_L g2245 ( 
.A(n_1939),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1840),
.B(n_1862),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1873),
.B(n_1060),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1996),
.B(n_1061),
.Y(n_2248)
);

OR2x6_ASAP7_75t_L g2249 ( 
.A(n_1763),
.B(n_922),
.Y(n_2249)
);

BUFx2_ASAP7_75t_L g2250 ( 
.A(n_1944),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1778),
.B(n_1063),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1759),
.B(n_1064),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1823),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1841),
.B(n_1065),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1864),
.B(n_1067),
.Y(n_2255)
);

INVxp67_ASAP7_75t_SL g2256 ( 
.A(n_2011),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_1964),
.B(n_1068),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_1842),
.B(n_1074),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2011),
.B(n_1076),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1735),
.Y(n_2260)
);

O2A1O1Ixp33_ASAP7_75t_L g2261 ( 
.A1(n_1946),
.A2(n_1130),
.B(n_1133),
.C(n_1127),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1842),
.B(n_1077),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1869),
.B(n_1163),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1839),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1735),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1889),
.B(n_1078),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1952),
.B(n_1083),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1843),
.B(n_1084),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1849),
.B(n_1085),
.Y(n_2269)
);

INVx2_ASAP7_75t_SL g2270 ( 
.A(n_1955),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1855),
.B(n_1086),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1990),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_1830),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1858),
.B(n_1088),
.Y(n_2274)
);

OR2x2_ASAP7_75t_L g2275 ( 
.A(n_1890),
.B(n_1089),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1863),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1865),
.B(n_1094),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_1948),
.B(n_1096),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_1981),
.A2(n_1231),
.B1(n_1140),
.B2(n_1144),
.Y(n_2279)
);

AND3x1_ASAP7_75t_L g2280 ( 
.A(n_1970),
.B(n_1149),
.C(n_1137),
.Y(n_2280)
);

AOI22xp33_ASAP7_75t_L g2281 ( 
.A1(n_1880),
.A2(n_1153),
.B1(n_1155),
.B2(n_1151),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_1914),
.B(n_1097),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2003),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2007),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_1933),
.B(n_1300),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2009),
.B(n_1100),
.Y(n_2286)
);

NAND2xp33_ASAP7_75t_L g2287 ( 
.A(n_1883),
.B(n_1231),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_1949),
.B(n_1102),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2012),
.B(n_1103),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_1956),
.B(n_1111),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1837),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_L g2292 ( 
.A(n_1958),
.B(n_1114),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1837),
.Y(n_2293)
);

OAI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_1779),
.A2(n_1187),
.B1(n_1190),
.B2(n_1157),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1954),
.B(n_1118),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_1833),
.B(n_1122),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_1959),
.B(n_1123),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1737),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1987),
.B(n_1129),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_1968),
.B(n_1132),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1833),
.B(n_1134),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1837),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_1957),
.B(n_1136),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_1969),
.B(n_1138),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_1957),
.B(n_1139),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_1966),
.B(n_1142),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_1791),
.A2(n_1211),
.B1(n_1217),
.B2(n_1207),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1874),
.B(n_1148),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1874),
.B(n_1150),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_1965),
.B(n_1167),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1737),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1874),
.B(n_1168),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_1737),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_1836),
.A2(n_1231),
.B1(n_1229),
.B2(n_1223),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_1965),
.B(n_1169),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_1888),
.B(n_1170),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_SL g2317 ( 
.A(n_1957),
.B(n_1173),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1836),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1878),
.B(n_1174),
.Y(n_2319)
);

OAI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_1802),
.A2(n_1249),
.B1(n_1255),
.B2(n_1247),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_1963),
.B(n_1271),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_SL g2322 ( 
.A(n_1817),
.B(n_1300),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_1742),
.Y(n_2323)
);

INVx4_ASAP7_75t_L g2324 ( 
.A(n_1830),
.Y(n_2324)
);

NAND3xp33_ASAP7_75t_L g2325 ( 
.A(n_1963),
.B(n_1184),
.C(n_1179),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1878),
.B(n_1189),
.Y(n_2326)
);

OAI22xp33_ASAP7_75t_L g2327 ( 
.A1(n_1967),
.A2(n_1200),
.B1(n_1201),
.B2(n_1191),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_L g2328 ( 
.A(n_1854),
.B(n_1203),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_1878),
.B(n_1202),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_1854),
.B(n_1218),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_1742),
.B(n_1206),
.Y(n_2331)
);

NOR2xp33_ASAP7_75t_L g2332 ( 
.A(n_1898),
.B(n_1222),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1860),
.B(n_1809),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_1742),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_1898),
.B(n_1225),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1816),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_1836),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_1860),
.B(n_1219),
.Y(n_2338)
);

OAI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_1911),
.A2(n_1274),
.B(n_1273),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1860),
.B(n_1227),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_1963),
.B(n_1230),
.Y(n_2341)
);

INVx4_ASAP7_75t_L g2342 ( 
.A(n_1817),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1835),
.B(n_1235),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_1729),
.B(n_1236),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1768),
.B(n_1241),
.Y(n_2345)
);

AOI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_1903),
.A2(n_1279),
.B1(n_1280),
.B2(n_1276),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1775),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1785),
.B(n_1244),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_1816),
.B(n_1246),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_1793),
.A2(n_1291),
.B(n_1281),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_2045),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2188),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2017),
.B(n_1796),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2016),
.B(n_1971),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_R g2355 ( 
.A(n_2157),
.B(n_1748),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2284),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2272),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2283),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2131),
.B(n_2100),
.Y(n_2359)
);

BUFx4f_ASAP7_75t_L g2360 ( 
.A(n_2240),
.Y(n_2360)
);

BUFx3_ASAP7_75t_L g2361 ( 
.A(n_2188),
.Y(n_2361)
);

CKINVDCx6p67_ASAP7_75t_R g2362 ( 
.A(n_2324),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2035),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2025),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2088),
.B(n_1894),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2033),
.B(n_1798),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2050),
.B(n_1818),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2068),
.Y(n_2368)
);

AND2x6_ASAP7_75t_L g2369 ( 
.A(n_2053),
.B(n_1816),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2071),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_2053),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2084),
.B(n_1300),
.Y(n_2372)
);

BUFx3_ASAP7_75t_L g2373 ( 
.A(n_2222),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_2053),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_2067),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2081),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2099),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2119),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2097),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2030),
.B(n_1971),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2108),
.Y(n_2381)
);

BUFx3_ASAP7_75t_L g2382 ( 
.A(n_2250),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_R g2383 ( 
.A(n_2322),
.B(n_1826),
.Y(n_2383)
);

INVx4_ASAP7_75t_L g2384 ( 
.A(n_2324),
.Y(n_2384)
);

NAND2x1p5_ASAP7_75t_L g2385 ( 
.A(n_2342),
.B(n_1872),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2165),
.B(n_1821),
.Y(n_2386)
);

NOR3xp33_ASAP7_75t_SL g2387 ( 
.A(n_2014),
.B(n_1252),
.C(n_1248),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2135),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2105),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2171),
.B(n_1299),
.Y(n_2390)
);

BUFx3_ASAP7_75t_L g2391 ( 
.A(n_2152),
.Y(n_2391)
);

BUFx6f_ASAP7_75t_L g2392 ( 
.A(n_2070),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_R g2393 ( 
.A(n_2075),
.B(n_1852),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_R g2394 ( 
.A(n_2204),
.B(n_1256),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2195),
.B(n_2174),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_2038),
.B(n_1872),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2064),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2170),
.B(n_1257),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2175),
.B(n_1302),
.Y(n_2399)
);

BUFx3_ASAP7_75t_L g2400 ( 
.A(n_2342),
.Y(n_2400)
);

AND3x1_ASAP7_75t_SL g2401 ( 
.A(n_2142),
.B(n_1318),
.C(n_1305),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_2070),
.Y(n_2402)
);

INVx5_ASAP7_75t_L g2403 ( 
.A(n_2147),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_SL g2404 ( 
.A(n_2147),
.B(n_1883),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2141),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2150),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2176),
.B(n_1319),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_L g2408 ( 
.A(n_2228),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2191),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_2026),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2226),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2116),
.Y(n_2412)
);

BUFx12f_ASAP7_75t_L g2413 ( 
.A(n_2200),
.Y(n_2413)
);

NOR3xp33_ASAP7_75t_SL g2414 ( 
.A(n_2124),
.B(n_2294),
.C(n_2107),
.Y(n_2414)
);

BUFx3_ASAP7_75t_L g2415 ( 
.A(n_2200),
.Y(n_2415)
);

INVx4_ASAP7_75t_L g2416 ( 
.A(n_2147),
.Y(n_2416)
);

HB1xp67_ASAP7_75t_L g2417 ( 
.A(n_2027),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_R g2418 ( 
.A(n_2273),
.B(n_1260),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_2057),
.Y(n_2419)
);

INVx5_ASAP7_75t_L g2420 ( 
.A(n_2185),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2072),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2122),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_SL g2423 ( 
.A(n_2034),
.B(n_1266),
.C(n_1264),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2264),
.Y(n_2424)
);

AOI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2123),
.A2(n_2094),
.B1(n_2121),
.B2(n_2058),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_2070),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_2110),
.B(n_1326),
.Y(n_2427)
);

NOR2xp33_ASAP7_75t_L g2428 ( 
.A(n_2129),
.B(n_1267),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_2057),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2144),
.B(n_1270),
.Y(n_2430)
);

CKINVDCx20_ASAP7_75t_R g2431 ( 
.A(n_2124),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2276),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_2089),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_2115),
.B(n_1277),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2196),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2180),
.B(n_1330),
.Y(n_2436)
);

INVx4_ASAP7_75t_SL g2437 ( 
.A(n_2185),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2148),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2126),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2182),
.B(n_1353),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_2089),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2032),
.B(n_1354),
.Y(n_2442)
);

AOI22xp33_ASAP7_75t_L g2443 ( 
.A1(n_2230),
.A2(n_1289),
.B1(n_1290),
.B2(n_1283),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2082),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2153),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2155),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2038),
.B(n_1872),
.Y(n_2447)
);

CKINVDCx20_ASAP7_75t_R g2448 ( 
.A(n_2245),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2253),
.B(n_1358),
.Y(n_2449)
);

AND2x4_ASAP7_75t_L g2450 ( 
.A(n_2132),
.B(n_1359),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2113),
.B(n_1364),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2217),
.B(n_1367),
.Y(n_2452)
);

INVx4_ASAP7_75t_L g2453 ( 
.A(n_2233),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2046),
.B(n_1381),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2145),
.B(n_1293),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2020),
.B(n_1882),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2166),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2177),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2201),
.B(n_1882),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2194),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2327),
.B(n_1882),
.Y(n_2461)
);

AND3x2_ASAP7_75t_SL g2462 ( 
.A(n_2128),
.B(n_1372),
.C(n_1363),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2197),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2091),
.B(n_1932),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_2085),
.Y(n_2465)
);

NOR2xp33_ASAP7_75t_R g2466 ( 
.A(n_2134),
.B(n_1295),
.Y(n_2466)
);

BUFx3_ASAP7_75t_L g2467 ( 
.A(n_2219),
.Y(n_2467)
);

CKINVDCx20_ASAP7_75t_R g2468 ( 
.A(n_2233),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2140),
.B(n_1932),
.Y(n_2469)
);

BUFx12f_ASAP7_75t_L g2470 ( 
.A(n_2233),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2220),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2208),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_2078),
.B(n_1298),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2208),
.Y(n_2474)
);

CKINVDCx20_ASAP7_75t_R g2475 ( 
.A(n_2249),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2223),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2275),
.B(n_2282),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2145),
.B(n_1303),
.Y(n_2478)
);

INVx4_ASAP7_75t_L g2479 ( 
.A(n_2249),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2151),
.B(n_1932),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_L g2481 ( 
.A1(n_2042),
.A2(n_1317),
.B1(n_1320),
.B2(n_1306),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2015),
.Y(n_2482)
);

NOR3xp33_ASAP7_75t_SL g2483 ( 
.A(n_2158),
.B(n_1324),
.C(n_1323),
.Y(n_2483)
);

NOR3xp33_ASAP7_75t_SL g2484 ( 
.A(n_2328),
.B(n_1343),
.C(n_1325),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2015),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2280),
.B(n_1345),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_SL g2487 ( 
.A(n_2041),
.B(n_1346),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_2139),
.Y(n_2488)
);

INVxp67_ASAP7_75t_SL g2489 ( 
.A(n_2208),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2244),
.B(n_922),
.Y(n_2490)
);

INVx4_ASAP7_75t_L g2491 ( 
.A(n_2249),
.Y(n_2491)
);

O2A1O1Ixp33_ASAP7_75t_L g2492 ( 
.A1(n_2066),
.A2(n_2093),
.B(n_2083),
.C(n_2229),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2133),
.Y(n_2493)
);

BUFx2_ASAP7_75t_L g2494 ( 
.A(n_2079),
.Y(n_2494)
);

AND2x4_ASAP7_75t_L g2495 ( 
.A(n_2164),
.B(n_936),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2207),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2211),
.Y(n_2497)
);

HB1xp67_ASAP7_75t_L g2498 ( 
.A(n_2077),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2218),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2019),
.B(n_936),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2184),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2235),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_2072),
.Y(n_2503)
);

NOR3xp33_ASAP7_75t_SL g2504 ( 
.A(n_2330),
.B(n_1355),
.C(n_1348),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2051),
.B(n_975),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2056),
.B(n_975),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2257),
.B(n_1360),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2022),
.B(n_1039),
.Y(n_2508)
);

BUFx3_ASAP7_75t_L g2509 ( 
.A(n_2238),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2347),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2023),
.B(n_1039),
.Y(n_2511)
);

BUFx12f_ASAP7_75t_L g2512 ( 
.A(n_2270),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2060),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2060),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2321),
.Y(n_2515)
);

AND2x6_ASAP7_75t_L g2516 ( 
.A(n_2215),
.B(n_1072),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2321),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2079),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_2215),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2215),
.Y(n_2520)
);

INVx4_ASAP7_75t_L g2521 ( 
.A(n_2077),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2239),
.A2(n_1380),
.B1(n_943),
.B2(n_961),
.Y(n_2522)
);

NOR3xp33_ASAP7_75t_SL g2523 ( 
.A(n_2332),
.B(n_3),
.C(n_4),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2087),
.B(n_1072),
.Y(n_2524)
);

INVx1_ASAP7_75t_SL g2525 ( 
.A(n_2341),
.Y(n_2525)
);

AND2x4_ASAP7_75t_L g2526 ( 
.A(n_2164),
.B(n_1164),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2137),
.B(n_1164),
.Y(n_2527)
);

XNOR2xp5_ASAP7_75t_L g2528 ( 
.A(n_2087),
.B(n_4),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2169),
.Y(n_2529)
);

INVx3_ASAP7_75t_L g2530 ( 
.A(n_2013),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2021),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2077),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2214),
.B(n_1198),
.Y(n_2533)
);

BUFx3_ASAP7_75t_L g2534 ( 
.A(n_2185),
.Y(n_2534)
);

AOI22xp33_ASAP7_75t_SL g2535 ( 
.A1(n_2130),
.A2(n_943),
.B1(n_961),
.B2(n_866),
.Y(n_2535)
);

AND2x4_ASAP7_75t_L g2536 ( 
.A(n_2246),
.B(n_1198),
.Y(n_2536)
);

INVx5_ASAP7_75t_L g2537 ( 
.A(n_2185),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2044),
.B(n_866),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2043),
.B(n_1262),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_2316),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2103),
.B(n_1262),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2069),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2190),
.Y(n_2543)
);

BUFx2_ASAP7_75t_L g2544 ( 
.A(n_2203),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2190),
.Y(n_2545)
);

BUFx3_ASAP7_75t_L g2546 ( 
.A(n_2263),
.Y(n_2546)
);

AOI211xp5_ASAP7_75t_L g2547 ( 
.A1(n_2173),
.A2(n_1363),
.B(n_1372),
.C(n_1284),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2298),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2311),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2062),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2052),
.B(n_1284),
.Y(n_2551)
);

NOR3xp33_ASAP7_75t_SL g2552 ( 
.A(n_2335),
.B(n_4),
.C(n_5),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2054),
.B(n_2111),
.Y(n_2553)
);

AND2x4_ASAP7_75t_L g2554 ( 
.A(n_2303),
.B(n_1903),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2013),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_R g2556 ( 
.A(n_2172),
.B(n_5),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2285),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2073),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2074),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2076),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2080),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2313),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_2305),
.B(n_1903),
.Y(n_2563)
);

NAND2x1p5_ASAP7_75t_L g2564 ( 
.A(n_2216),
.B(n_2018),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2310),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2047),
.B(n_5),
.Y(n_2566)
);

INVx1_ASAP7_75t_SL g2567 ( 
.A(n_2301),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2286),
.B(n_6),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2289),
.B(n_2092),
.Y(n_2569)
);

BUFx12f_ASAP7_75t_L g2570 ( 
.A(n_2317),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2292),
.B(n_6),
.Y(n_2571)
);

AOI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2315),
.A2(n_2156),
.B1(n_2181),
.B2(n_2297),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2102),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2146),
.B(n_2149),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2104),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2106),
.B(n_6),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2323),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2114),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2117),
.Y(n_2579)
);

INVx3_ASAP7_75t_L g2580 ( 
.A(n_2036),
.Y(n_2580)
);

NOR3xp33_ASAP7_75t_SL g2581 ( 
.A(n_2325),
.B(n_7),
.C(n_8),
.Y(n_2581)
);

INVx2_ASAP7_75t_SL g2582 ( 
.A(n_2296),
.Y(n_2582)
);

NOR3xp33_ASAP7_75t_SL g2583 ( 
.A(n_2154),
.B(n_2112),
.C(n_2031),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2346),
.B(n_866),
.Y(n_2584)
);

CKINVDCx20_ASAP7_75t_R g2585 ( 
.A(n_2346),
.Y(n_2585)
);

INVx5_ASAP7_75t_L g2586 ( 
.A(n_2243),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2118),
.Y(n_2587)
);

BUFx2_ASAP7_75t_L g2588 ( 
.A(n_2308),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2232),
.B(n_2278),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2199),
.B(n_7),
.Y(n_2590)
);

BUFx3_ASAP7_75t_L g2591 ( 
.A(n_2309),
.Y(n_2591)
);

A2O1A1Ixp33_ASAP7_75t_L g2592 ( 
.A1(n_2199),
.A2(n_961),
.B(n_1036),
.C(n_943),
.Y(n_2592)
);

HB1xp67_ASAP7_75t_L g2593 ( 
.A(n_2320),
.Y(n_2593)
);

BUFx3_ASAP7_75t_L g2594 ( 
.A(n_2312),
.Y(n_2594)
);

OAI21xp33_ASAP7_75t_L g2595 ( 
.A1(n_2028),
.A2(n_961),
.B(n_943),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2300),
.Y(n_2596)
);

AND2x6_ASAP7_75t_L g2597 ( 
.A(n_2260),
.B(n_1036),
.Y(n_2597)
);

AND2x6_ASAP7_75t_SL g2598 ( 
.A(n_2304),
.B(n_7),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2334),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_2090),
.Y(n_2600)
);

OAI22xp5_ASAP7_75t_SL g2601 ( 
.A1(n_2198),
.A2(n_1101),
.B1(n_1113),
.B2(n_1036),
.Y(n_2601)
);

BUFx3_ASAP7_75t_L g2602 ( 
.A(n_2319),
.Y(n_2602)
);

BUFx4f_ASAP7_75t_L g2603 ( 
.A(n_2291),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2212),
.B(n_8),
.Y(n_2604)
);

BUFx2_ASAP7_75t_L g2605 ( 
.A(n_2329),
.Y(n_2605)
);

BUFx2_ASAP7_75t_L g2606 ( 
.A(n_2343),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2212),
.B(n_8),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2344),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2095),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2345),
.Y(n_2610)
);

INVx3_ASAP7_75t_L g2611 ( 
.A(n_2098),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2336),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2339),
.B(n_9),
.Y(n_2613)
);

A2O1A1Ixp33_ASAP7_75t_L g2614 ( 
.A1(n_2261),
.A2(n_1101),
.B(n_1113),
.C(n_1036),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_L g2615 ( 
.A(n_2055),
.B(n_9),
.Y(n_2615)
);

BUFx3_ASAP7_75t_L g2616 ( 
.A(n_2252),
.Y(n_2616)
);

NAND2x1p5_ASAP7_75t_L g2617 ( 
.A(n_2331),
.B(n_1101),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2024),
.B(n_9),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2193),
.B(n_10),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2265),
.Y(n_2620)
);

CKINVDCx5p33_ASAP7_75t_R g2621 ( 
.A(n_2213),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2096),
.Y(n_2622)
);

OR2x6_ASAP7_75t_L g2623 ( 
.A(n_2326),
.B(n_2205),
.Y(n_2623)
);

NAND3xp33_ASAP7_75t_SL g2624 ( 
.A(n_2241),
.B(n_1113),
.C(n_1101),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2183),
.B(n_10),
.Y(n_2625)
);

NOR3xp33_ASAP7_75t_SL g2626 ( 
.A(n_2037),
.B(n_11),
.C(n_12),
.Y(n_2626)
);

AND2x4_ASAP7_75t_SL g2627 ( 
.A(n_2307),
.B(n_1113),
.Y(n_2627)
);

NOR3xp33_ASAP7_75t_SL g2628 ( 
.A(n_2039),
.B(n_11),
.C(n_12),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2348),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2138),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2189),
.B(n_1272),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_R g2632 ( 
.A(n_2209),
.B(n_11),
.Y(n_2632)
);

BUFx6f_ASAP7_75t_L g2633 ( 
.A(n_2333),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2040),
.B(n_13),
.Y(n_2634)
);

INVx1_ASAP7_75t_SL g2635 ( 
.A(n_2258),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2029),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2268),
.Y(n_2637)
);

BUFx3_ASAP7_75t_L g2638 ( 
.A(n_2192),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2209),
.Y(n_2639)
);

INVx4_ASAP7_75t_L g2640 ( 
.A(n_2209),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2048),
.B(n_13),
.Y(n_2641)
);

AOI22xp33_ASAP7_75t_L g2642 ( 
.A1(n_2120),
.A2(n_1370),
.B1(n_1377),
.B2(n_1272),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2269),
.Y(n_2643)
);

INVxp67_ASAP7_75t_SL g2644 ( 
.A(n_2256),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2271),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2221),
.Y(n_2646)
);

OR2x2_ASAP7_75t_L g2647 ( 
.A(n_2224),
.B(n_14),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2209),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2266),
.B(n_14),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2274),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2227),
.Y(n_2651)
);

AND2x4_ASAP7_75t_SL g2652 ( 
.A(n_2202),
.B(n_2206),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_2267),
.Y(n_2653)
);

OR2x2_ASAP7_75t_L g2654 ( 
.A(n_2225),
.B(n_14),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2277),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2167),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2209),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2178),
.Y(n_2658)
);

AOI21xp5_ASAP7_75t_L g2659 ( 
.A1(n_2168),
.A2(n_1370),
.B(n_1272),
.Y(n_2659)
);

INVx5_ASAP7_75t_L g2660 ( 
.A(n_2287),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2236),
.Y(n_2661)
);

AOI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_2290),
.A2(n_1370),
.B1(n_1377),
.B2(n_1272),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_L g2663 ( 
.A(n_2231),
.B(n_15),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2143),
.Y(n_2664)
);

INVx2_ASAP7_75t_SL g2665 ( 
.A(n_2349),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2241),
.B(n_15),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2159),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2160),
.B(n_15),
.Y(n_2668)
);

BUFx2_ASAP7_75t_L g2669 ( 
.A(n_2262),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_R g2670 ( 
.A(n_2234),
.B(n_16),
.Y(n_2670)
);

BUFx2_ASAP7_75t_L g2671 ( 
.A(n_2338),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2179),
.Y(n_2672)
);

AND2x4_ASAP7_75t_L g2673 ( 
.A(n_2049),
.B(n_16),
.Y(n_2673)
);

NOR3xp33_ASAP7_75t_SL g2674 ( 
.A(n_2288),
.B(n_16),
.C(n_17),
.Y(n_2674)
);

NOR3xp33_ASAP7_75t_SL g2675 ( 
.A(n_2127),
.B(n_17),
.C(n_18),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2237),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2162),
.Y(n_2677)
);

OR2x2_ASAP7_75t_L g2678 ( 
.A(n_2242),
.B(n_17),
.Y(n_2678)
);

OR2x6_ASAP7_75t_L g2679 ( 
.A(n_2210),
.B(n_1370),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2293),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2281),
.B(n_18),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2125),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2302),
.Y(n_2683)
);

NAND2xp33_ASAP7_75t_SL g2684 ( 
.A(n_2136),
.B(n_1377),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2340),
.B(n_1377),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2318),
.Y(n_2686)
);

INVx4_ASAP7_75t_L g2687 ( 
.A(n_2337),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2350),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2248),
.Y(n_2689)
);

INVx4_ASAP7_75t_L g2690 ( 
.A(n_2063),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2306),
.B(n_18),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2259),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2247),
.B(n_19),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2254),
.B(n_19),
.Y(n_2694)
);

BUFx6f_ASAP7_75t_L g2695 ( 
.A(n_2065),
.Y(n_2695)
);

INVx3_ASAP7_75t_L g2696 ( 
.A(n_2299),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2255),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2086),
.Y(n_2698)
);

BUFx6f_ASAP7_75t_L g2699 ( 
.A(n_2101),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_SL g2700 ( 
.A(n_2251),
.B(n_21),
.Y(n_2700)
);

BUFx4f_ASAP7_75t_L g2701 ( 
.A(n_2161),
.Y(n_2701)
);

BUFx3_ASAP7_75t_L g2702 ( 
.A(n_2314),
.Y(n_2702)
);

BUFx3_ASAP7_75t_L g2703 ( 
.A(n_2314),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2279),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2109),
.Y(n_2705)
);

NOR2xp33_ASAP7_75t_R g2706 ( 
.A(n_2059),
.B(n_20),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_2163),
.B(n_20),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2279),
.B(n_21),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2186),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2187),
.Y(n_2710)
);

BUFx2_ASAP7_75t_L g2711 ( 
.A(n_2295),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2061),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2324),
.B(n_21),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2017),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2284),
.Y(n_2715)
);

INVxp67_ASAP7_75t_L g2716 ( 
.A(n_2067),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2017),
.B(n_22),
.Y(n_2717)
);

BUFx2_ASAP7_75t_L g2718 ( 
.A(n_2045),
.Y(n_2718)
);

BUFx6f_ASAP7_75t_L g2719 ( 
.A(n_2053),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2016),
.B(n_23),
.Y(n_2720)
);

NAND2x1p5_ASAP7_75t_L g2721 ( 
.A(n_2324),
.B(n_22),
.Y(n_2721)
);

AND2x2_ASAP7_75t_SL g2722 ( 
.A(n_2131),
.B(n_22),
.Y(n_2722)
);

AND2x4_ASAP7_75t_L g2723 ( 
.A(n_2324),
.B(n_23),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2284),
.Y(n_2724)
);

NOR2xp33_ASAP7_75t_R g2725 ( 
.A(n_2157),
.B(n_24),
.Y(n_2725)
);

CKINVDCx20_ASAP7_75t_R g2726 ( 
.A(n_2188),
.Y(n_2726)
);

BUFx8_ASAP7_75t_L g2727 ( 
.A(n_2222),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2284),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2284),
.Y(n_2729)
);

BUFx2_ASAP7_75t_L g2730 ( 
.A(n_2045),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2017),
.Y(n_2731)
);

NOR3xp33_ASAP7_75t_SL g2732 ( 
.A(n_2014),
.B(n_24),
.C(n_25),
.Y(n_2732)
);

INVx3_ASAP7_75t_L g2733 ( 
.A(n_2072),
.Y(n_2733)
);

BUFx2_ASAP7_75t_L g2734 ( 
.A(n_2045),
.Y(n_2734)
);

BUFx6f_ASAP7_75t_L g2735 ( 
.A(n_2053),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2017),
.Y(n_2736)
);

NOR3xp33_ASAP7_75t_SL g2737 ( 
.A(n_2014),
.B(n_24),
.C(n_25),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2017),
.B(n_25),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2284),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2017),
.B(n_26),
.Y(n_2740)
);

NOR2xp33_ASAP7_75t_SL g2741 ( 
.A(n_2147),
.B(n_26),
.Y(n_2741)
);

INVx3_ASAP7_75t_L g2742 ( 
.A(n_2072),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2017),
.B(n_26),
.Y(n_2743)
);

CKINVDCx5p33_ASAP7_75t_R g2744 ( 
.A(n_2188),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2017),
.B(n_27),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2017),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2284),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2017),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2017),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2017),
.B(n_27),
.Y(n_2750)
);

INVx5_ASAP7_75t_L g2751 ( 
.A(n_2147),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_R g2752 ( 
.A(n_2157),
.B(n_28),
.Y(n_2752)
);

INVx3_ASAP7_75t_L g2753 ( 
.A(n_2072),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2017),
.B(n_29),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2016),
.B(n_29),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2235),
.A2(n_29),
.B(n_30),
.Y(n_2756)
);

AND3x1_ASAP7_75t_SL g2757 ( 
.A(n_2142),
.B(n_30),
.C(n_31),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2017),
.B(n_31),
.Y(n_2758)
);

BUFx3_ASAP7_75t_L g2759 ( 
.A(n_2188),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2045),
.Y(n_2760)
);

INVx4_ASAP7_75t_L g2761 ( 
.A(n_2324),
.Y(n_2761)
);

HB1xp67_ASAP7_75t_L g2762 ( 
.A(n_2045),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2017),
.Y(n_2763)
);

INVx5_ASAP7_75t_L g2764 ( 
.A(n_2147),
.Y(n_2764)
);

OR2x2_ASAP7_75t_L g2765 ( 
.A(n_2045),
.B(n_32),
.Y(n_2765)
);

HB1xp67_ASAP7_75t_L g2766 ( 
.A(n_2045),
.Y(n_2766)
);

BUFx2_ASAP7_75t_L g2767 ( 
.A(n_2045),
.Y(n_2767)
);

BUFx2_ASAP7_75t_L g2768 ( 
.A(n_2045),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2017),
.B(n_32),
.Y(n_2769)
);

AND2x4_ASAP7_75t_L g2770 ( 
.A(n_2324),
.B(n_33),
.Y(n_2770)
);

NOR2x1p5_ASAP7_75t_L g2771 ( 
.A(n_2014),
.B(n_33),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2284),
.Y(n_2772)
);

INVx1_ASAP7_75t_SL g2773 ( 
.A(n_2016),
.Y(n_2773)
);

INVx4_ASAP7_75t_L g2774 ( 
.A(n_2324),
.Y(n_2774)
);

NOR3xp33_ASAP7_75t_SL g2775 ( 
.A(n_2014),
.B(n_33),
.C(n_34),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2017),
.Y(n_2776)
);

OR2x6_ASAP7_75t_SL g2777 ( 
.A(n_2064),
.B(n_36),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2017),
.B(n_35),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2017),
.B(n_36),
.Y(n_2779)
);

INVx4_ASAP7_75t_L g2780 ( 
.A(n_2324),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2284),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2017),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2284),
.Y(n_2783)
);

BUFx10_ASAP7_75t_L g2784 ( 
.A(n_2273),
.Y(n_2784)
);

INVx2_ASAP7_75t_SL g2785 ( 
.A(n_2188),
.Y(n_2785)
);

OR2x2_ASAP7_75t_L g2786 ( 
.A(n_2045),
.B(n_36),
.Y(n_2786)
);

AO22x1_ASAP7_75t_L g2787 ( 
.A1(n_2188),
.A2(n_39),
.B1(n_40),
.B2(n_38),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2017),
.B(n_37),
.Y(n_2788)
);

INVx3_ASAP7_75t_L g2789 ( 
.A(n_2072),
.Y(n_2789)
);

AOI22xp33_ASAP7_75t_L g2790 ( 
.A1(n_2131),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2284),
.Y(n_2791)
);

OAI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2038),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_2792)
);

NOR3xp33_ASAP7_75t_SL g2793 ( 
.A(n_2014),
.B(n_40),
.C(n_42),
.Y(n_2793)
);

INVxp67_ASAP7_75t_SL g2794 ( 
.A(n_2053),
.Y(n_2794)
);

BUFx6f_ASAP7_75t_L g2795 ( 
.A(n_2053),
.Y(n_2795)
);

HB1xp67_ASAP7_75t_L g2796 ( 
.A(n_2045),
.Y(n_2796)
);

BUFx3_ASAP7_75t_L g2797 ( 
.A(n_2188),
.Y(n_2797)
);

HB1xp67_ASAP7_75t_L g2798 ( 
.A(n_2045),
.Y(n_2798)
);

BUFx2_ASAP7_75t_L g2799 ( 
.A(n_2045),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2284),
.Y(n_2800)
);

BUFx3_ASAP7_75t_L g2801 ( 
.A(n_2188),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_2188),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2284),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2017),
.Y(n_2804)
);

BUFx3_ASAP7_75t_L g2805 ( 
.A(n_2188),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2017),
.B(n_42),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2017),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2284),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2045),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2017),
.B(n_42),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2016),
.B(n_44),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2284),
.Y(n_2812)
);

INVx4_ASAP7_75t_L g2813 ( 
.A(n_2324),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2017),
.Y(n_2814)
);

AND3x1_ASAP7_75t_SL g2815 ( 
.A(n_2142),
.B(n_51),
.C(n_43),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2017),
.Y(n_2816)
);

INVx5_ASAP7_75t_L g2817 ( 
.A(n_2147),
.Y(n_2817)
);

NAND2x1p5_ASAP7_75t_L g2818 ( 
.A(n_2324),
.B(n_44),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2017),
.B(n_44),
.Y(n_2819)
);

INVx5_ASAP7_75t_L g2820 ( 
.A(n_2147),
.Y(n_2820)
);

AOI22xp33_ASAP7_75t_L g2821 ( 
.A1(n_2131),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2017),
.B(n_46),
.Y(n_2822)
);

INVx4_ASAP7_75t_L g2823 ( 
.A(n_2324),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2284),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2017),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2017),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_R g2827 ( 
.A(n_2157),
.B(n_46),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2284),
.Y(n_2828)
);

INVx2_ASAP7_75t_SL g2829 ( 
.A(n_2188),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_R g2830 ( 
.A(n_2157),
.B(n_47),
.Y(n_2830)
);

AND2x4_ASAP7_75t_L g2831 ( 
.A(n_2324),
.B(n_47),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2016),
.B(n_49),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2324),
.B(n_48),
.Y(n_2833)
);

NOR2xp67_ASAP7_75t_L g2834 ( 
.A(n_2045),
.B(n_48),
.Y(n_2834)
);

BUFx2_ASAP7_75t_L g2835 ( 
.A(n_2045),
.Y(n_2835)
);

NOR2xp67_ASAP7_75t_L g2836 ( 
.A(n_2045),
.B(n_48),
.Y(n_2836)
);

INVx3_ASAP7_75t_L g2837 ( 
.A(n_2072),
.Y(n_2837)
);

CKINVDCx8_ASAP7_75t_R g2838 ( 
.A(n_2057),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2017),
.B(n_49),
.Y(n_2839)
);

NOR2xp33_ASAP7_75t_L g2840 ( 
.A(n_2088),
.B(n_49),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2284),
.Y(n_2841)
);

BUFx2_ASAP7_75t_L g2842 ( 
.A(n_2045),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2017),
.B(n_50),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2084),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2017),
.B(n_50),
.Y(n_2845)
);

AND2x4_ASAP7_75t_L g2846 ( 
.A(n_2324),
.B(n_51),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2045),
.Y(n_2847)
);

INVx3_ASAP7_75t_SL g2848 ( 
.A(n_2324),
.Y(n_2848)
);

OAI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2235),
.A2(n_52),
.B(n_53),
.Y(n_2849)
);

CKINVDCx20_ASAP7_75t_R g2850 ( 
.A(n_2188),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2017),
.Y(n_2851)
);

CKINVDCx8_ASAP7_75t_R g2852 ( 
.A(n_2057),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2017),
.Y(n_2853)
);

AOI22xp33_ASAP7_75t_L g2854 ( 
.A1(n_2131),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2854)
);

HB1xp67_ASAP7_75t_L g2855 ( 
.A(n_2045),
.Y(n_2855)
);

INVxp67_ASAP7_75t_L g2856 ( 
.A(n_2067),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2017),
.B(n_53),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2284),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2188),
.Y(n_2859)
);

AND2x6_ASAP7_75t_L g2860 ( 
.A(n_2053),
.B(n_55),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2017),
.B(n_54),
.Y(n_2861)
);

NOR2xp33_ASAP7_75t_R g2862 ( 
.A(n_2157),
.B(n_54),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2017),
.B(n_55),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2017),
.Y(n_2864)
);

INVx3_ASAP7_75t_L g2865 ( 
.A(n_2072),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2017),
.Y(n_2866)
);

INVx5_ASAP7_75t_L g2867 ( 
.A(n_2147),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2017),
.B(n_55),
.Y(n_2868)
);

BUFx6f_ASAP7_75t_L g2869 ( 
.A(n_2053),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2017),
.B(n_56),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2053),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2053),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2016),
.B(n_56),
.Y(n_2873)
);

AOI21x1_ASAP7_75t_L g2874 ( 
.A1(n_2396),
.A2(n_57),
.B(n_58),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2379),
.B(n_57),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2381),
.B(n_57),
.Y(n_2876)
);

OAI21x1_ASAP7_75t_L g2877 ( 
.A1(n_2502),
.A2(n_59),
.B(n_60),
.Y(n_2877)
);

OAI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2593),
.A2(n_2585),
.B1(n_2792),
.B2(n_2535),
.Y(n_2878)
);

OAI21xp33_ASAP7_75t_L g2879 ( 
.A1(n_2556),
.A2(n_59),
.B(n_60),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2593),
.B(n_2435),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2397),
.B(n_61),
.Y(n_2881)
);

OA21x2_ASAP7_75t_L g2882 ( 
.A1(n_2682),
.A2(n_61),
.B(n_63),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2397),
.B(n_63),
.Y(n_2883)
);

OAI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2792),
.A2(n_2535),
.B1(n_2613),
.B2(n_2702),
.Y(n_2884)
);

AOI21xp33_ASAP7_75t_L g2885 ( 
.A1(n_2569),
.A2(n_64),
.B(n_65),
.Y(n_2885)
);

INVx2_ASAP7_75t_SL g2886 ( 
.A(n_2413),
.Y(n_2886)
);

AO21x2_ASAP7_75t_L g2887 ( 
.A1(n_2624),
.A2(n_64),
.B(n_65),
.Y(n_2887)
);

INVx2_ASAP7_75t_SL g2888 ( 
.A(n_2727),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2619),
.B(n_2550),
.Y(n_2889)
);

OAI21x1_ASAP7_75t_L g2890 ( 
.A1(n_2489),
.A2(n_64),
.B(n_65),
.Y(n_2890)
);

AND2x4_ASAP7_75t_L g2891 ( 
.A(n_2384),
.B(n_2761),
.Y(n_2891)
);

BUFx3_ASAP7_75t_L g2892 ( 
.A(n_2848),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2370),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2558),
.B(n_66),
.Y(n_2894)
);

AOI21xp5_ASAP7_75t_L g2895 ( 
.A1(n_2553),
.A2(n_66),
.B(n_67),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2376),
.Y(n_2896)
);

AND2x4_ASAP7_75t_L g2897 ( 
.A(n_2384),
.B(n_68),
.Y(n_2897)
);

OAI21x1_ASAP7_75t_L g2898 ( 
.A1(n_2794),
.A2(n_68),
.B(n_69),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2848),
.Y(n_2899)
);

AOI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_2553),
.A2(n_69),
.B(n_70),
.Y(n_2900)
);

OAI21x1_ASAP7_75t_L g2901 ( 
.A1(n_2794),
.A2(n_2659),
.B(n_2648),
.Y(n_2901)
);

OAI21x1_ASAP7_75t_L g2902 ( 
.A1(n_2659),
.A2(n_69),
.B(n_70),
.Y(n_2902)
);

OAI21x1_ASAP7_75t_L g2903 ( 
.A1(n_2639),
.A2(n_71),
.B(n_72),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2364),
.Y(n_2904)
);

BUFx3_ASAP7_75t_L g2905 ( 
.A(n_2362),
.Y(n_2905)
);

OAI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2569),
.A2(n_71),
.B(n_72),
.Y(n_2906)
);

OAI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2704),
.A2(n_72),
.B(n_73),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_2494),
.B(n_73),
.Y(n_2908)
);

OAI21xp33_ASAP7_75t_SL g2909 ( 
.A1(n_2849),
.A2(n_2722),
.B(n_2613),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2395),
.B(n_74),
.Y(n_2910)
);

AOI221x1_ASAP7_75t_L g2911 ( 
.A1(n_2756),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.C(n_77),
.Y(n_2911)
);

OAI21x1_ASAP7_75t_L g2912 ( 
.A1(n_2657),
.A2(n_74),
.B(n_75),
.Y(n_2912)
);

OAI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2649),
.A2(n_76),
.B(n_77),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2703),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2368),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_SL g2916 ( 
.A(n_2773),
.B(n_305),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2356),
.Y(n_2917)
);

OAI21x1_ASAP7_75t_L g2918 ( 
.A1(n_2469),
.A2(n_78),
.B(n_79),
.Y(n_2918)
);

NAND2x1p5_ASAP7_75t_L g2919 ( 
.A(n_2761),
.B(n_80),
.Y(n_2919)
);

CKINVDCx20_ASAP7_75t_R g2920 ( 
.A(n_2726),
.Y(n_2920)
);

OAI21x1_ASAP7_75t_SL g2921 ( 
.A1(n_2849),
.A2(n_80),
.B(n_81),
.Y(n_2921)
);

INVx2_ASAP7_75t_SL g2922 ( 
.A(n_2727),
.Y(n_2922)
);

OAI21xp33_ASAP7_75t_L g2923 ( 
.A1(n_2425),
.A2(n_80),
.B(n_81),
.Y(n_2923)
);

OAI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2649),
.A2(n_82),
.B(n_83),
.Y(n_2924)
);

AOI21xp33_ASAP7_75t_L g2925 ( 
.A1(n_2492),
.A2(n_2634),
.B(n_2641),
.Y(n_2925)
);

AND2x2_ASAP7_75t_L g2926 ( 
.A(n_2359),
.B(n_2518),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2559),
.B(n_2560),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2774),
.B(n_2780),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2561),
.B(n_82),
.Y(n_2929)
);

AO31x2_ASAP7_75t_L g2930 ( 
.A1(n_2592),
.A2(n_84),
.A3(n_82),
.B(n_83),
.Y(n_2930)
);

O2A1O1Ixp33_ASAP7_75t_L g2931 ( 
.A1(n_2423),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2573),
.B(n_84),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2666),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_2933)
);

OA21x2_ASAP7_75t_L g2934 ( 
.A1(n_2595),
.A2(n_86),
.B(n_87),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2575),
.B(n_86),
.Y(n_2935)
);

NAND3xp33_ASAP7_75t_L g2936 ( 
.A(n_2523),
.B(n_88),
.C(n_89),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2377),
.Y(n_2937)
);

OAI21x1_ASAP7_75t_L g2938 ( 
.A1(n_2480),
.A2(n_88),
.B(n_89),
.Y(n_2938)
);

HB1xp67_ASAP7_75t_L g2939 ( 
.A(n_2760),
.Y(n_2939)
);

INVx8_ASAP7_75t_L g2940 ( 
.A(n_2860),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2500),
.A2(n_89),
.B(n_90),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_2850),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_2773),
.B(n_305),
.Y(n_2943)
);

OAI21x1_ASAP7_75t_L g2944 ( 
.A1(n_2357),
.A2(n_90),
.B(n_91),
.Y(n_2944)
);

AO21x1_ASAP7_75t_L g2945 ( 
.A1(n_2741),
.A2(n_307),
.B(n_306),
.Y(n_2945)
);

OAI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2360),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_2946)
);

A2O1A1Ixp33_ASAP7_75t_L g2947 ( 
.A1(n_2691),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2360),
.B(n_306),
.Y(n_2948)
);

AO31x2_ASAP7_75t_L g2949 ( 
.A1(n_2756),
.A2(n_94),
.A3(n_92),
.B(n_93),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2500),
.A2(n_95),
.B(n_96),
.Y(n_2950)
);

OAI21x1_ASAP7_75t_L g2951 ( 
.A1(n_2358),
.A2(n_95),
.B(n_96),
.Y(n_2951)
);

OAI22x1_ASAP7_75t_L g2952 ( 
.A1(n_2528),
.A2(n_98),
.B1(n_95),
.B2(n_97),
.Y(n_2952)
);

OAI21x1_ASAP7_75t_L g2953 ( 
.A1(n_2680),
.A2(n_97),
.B(n_98),
.Y(n_2953)
);

OAI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2666),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2578),
.B(n_99),
.Y(n_2955)
);

HB1xp67_ASAP7_75t_L g2956 ( 
.A(n_2760),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2715),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2708),
.A2(n_100),
.B(n_101),
.Y(n_2958)
);

OAI22x1_ASAP7_75t_L g2959 ( 
.A1(n_2721),
.A2(n_2818),
.B1(n_2771),
.B2(n_2488),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2579),
.B(n_100),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2762),
.B(n_102),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2355),
.B(n_308),
.Y(n_2962)
);

NAND3xp33_ASAP7_75t_L g2963 ( 
.A(n_2523),
.B(n_102),
.C(n_103),
.Y(n_2963)
);

OR2x6_ASAP7_75t_L g2964 ( 
.A(n_2470),
.B(n_102),
.Y(n_2964)
);

OAI21x1_ASAP7_75t_L g2965 ( 
.A1(n_2683),
.A2(n_103),
.B(n_104),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2378),
.Y(n_2966)
);

AOI211x1_ASAP7_75t_L g2967 ( 
.A1(n_2787),
.A2(n_2423),
.B(n_2668),
.C(n_2634),
.Y(n_2967)
);

OAI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2708),
.A2(n_104),
.B(n_105),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2714),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2418),
.B(n_308),
.Y(n_2970)
);

OAI21x1_ASAP7_75t_L g2971 ( 
.A1(n_2686),
.A2(n_105),
.B(n_106),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2724),
.Y(n_2972)
);

AOI21xp5_ASAP7_75t_L g2973 ( 
.A1(n_2456),
.A2(n_105),
.B(n_106),
.Y(n_2973)
);

O2A1O1Ixp33_ASAP7_75t_L g2974 ( 
.A1(n_2720),
.A2(n_108),
.B(n_106),
.C(n_107),
.Y(n_2974)
);

AND2x4_ASAP7_75t_L g2975 ( 
.A(n_2774),
.B(n_108),
.Y(n_2975)
);

OAI21x1_ASAP7_75t_L g2976 ( 
.A1(n_2456),
.A2(n_108),
.B(n_109),
.Y(n_2976)
);

AOI21xp5_ASAP7_75t_L g2977 ( 
.A1(n_2508),
.A2(n_109),
.B(n_110),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2587),
.B(n_2664),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2371),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2667),
.B(n_111),
.Y(n_2980)
);

OAI21x1_ASAP7_75t_L g2981 ( 
.A1(n_2600),
.A2(n_112),
.B(n_113),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2728),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2677),
.B(n_112),
.Y(n_2983)
);

AO31x2_ASAP7_75t_L g2984 ( 
.A1(n_2614),
.A2(n_114),
.A3(n_112),
.B(n_113),
.Y(n_2984)
);

INVx1_ASAP7_75t_SL g2985 ( 
.A(n_2375),
.Y(n_2985)
);

O2A1O1Ixp5_ASAP7_75t_L g2986 ( 
.A1(n_2461),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2729),
.Y(n_2987)
);

NOR2xp67_ASAP7_75t_L g2988 ( 
.A(n_2403),
.B(n_116),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2725),
.B(n_309),
.Y(n_2989)
);

BUFx12f_ASAP7_75t_L g2990 ( 
.A(n_2744),
.Y(n_2990)
);

BUFx2_ASAP7_75t_L g2991 ( 
.A(n_2448),
.Y(n_2991)
);

OAI21x1_ASAP7_75t_L g2992 ( 
.A1(n_2609),
.A2(n_115),
.B(n_116),
.Y(n_2992)
);

NAND2x1_ASAP7_75t_L g2993 ( 
.A(n_2860),
.B(n_116),
.Y(n_2993)
);

AOI21xp33_ASAP7_75t_L g2994 ( 
.A1(n_2492),
.A2(n_117),
.B(n_118),
.Y(n_2994)
);

OAI21xp5_ASAP7_75t_L g2995 ( 
.A1(n_2590),
.A2(n_117),
.B(n_118),
.Y(n_2995)
);

NOR2xp67_ASAP7_75t_SL g2996 ( 
.A(n_2802),
.B(n_117),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2661),
.B(n_118),
.Y(n_2997)
);

AOI21x1_ASAP7_75t_L g2998 ( 
.A1(n_2447),
.A2(n_119),
.B(n_120),
.Y(n_2998)
);

OAI21xp5_ASAP7_75t_SL g2999 ( 
.A1(n_2790),
.A2(n_119),
.B(n_120),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2731),
.Y(n_3000)
);

OAI21xp5_ASAP7_75t_L g3001 ( 
.A1(n_2590),
.A2(n_119),
.B(n_120),
.Y(n_3001)
);

OAI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_2604),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_3002)
);

INVx2_ASAP7_75t_SL g3003 ( 
.A(n_2784),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2752),
.B(n_310),
.Y(n_3004)
);

OR2x2_ASAP7_75t_L g3005 ( 
.A(n_2762),
.B(n_2766),
.Y(n_3005)
);

OAI21x1_ASAP7_75t_L g3006 ( 
.A1(n_2611),
.A2(n_123),
.B(n_124),
.Y(n_3006)
);

AO31x2_ASAP7_75t_L g3007 ( 
.A1(n_2688),
.A2(n_125),
.A3(n_123),
.B(n_124),
.Y(n_3007)
);

OAI21x1_ASAP7_75t_L g3008 ( 
.A1(n_2611),
.A2(n_124),
.B(n_125),
.Y(n_3008)
);

OAI21x1_ASAP7_75t_SL g3009 ( 
.A1(n_2640),
.A2(n_126),
.B(n_127),
.Y(n_3009)
);

OAI21x1_ASAP7_75t_L g3010 ( 
.A1(n_2464),
.A2(n_126),
.B(n_127),
.Y(n_3010)
);

OAI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2580),
.A2(n_128),
.B(n_129),
.Y(n_3011)
);

AOI21xp5_ASAP7_75t_L g3012 ( 
.A1(n_2508),
.A2(n_129),
.B(n_130),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2766),
.B(n_129),
.Y(n_3013)
);

OAI21x1_ASAP7_75t_L g3014 ( 
.A1(n_2580),
.A2(n_130),
.B(n_131),
.Y(n_3014)
);

INVxp67_ASAP7_75t_SL g3015 ( 
.A(n_2796),
.Y(n_3015)
);

INVx4_ASAP7_75t_L g3016 ( 
.A(n_2403),
.Y(n_3016)
);

OAI21x1_ASAP7_75t_L g3017 ( 
.A1(n_2385),
.A2(n_2685),
.B(n_2739),
.Y(n_3017)
);

OAI21x1_ASAP7_75t_L g3018 ( 
.A1(n_2385),
.A2(n_132),
.B(n_133),
.Y(n_3018)
);

CKINVDCx14_ASAP7_75t_R g3019 ( 
.A(n_2383),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2697),
.B(n_133),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2736),
.B(n_133),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2746),
.Y(n_3022)
);

OAI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2604),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_3023)
);

OAI21x1_ASAP7_75t_L g3024 ( 
.A1(n_2747),
.A2(n_134),
.B(n_135),
.Y(n_3024)
);

OA21x2_ASAP7_75t_L g3025 ( 
.A1(n_2490),
.A2(n_134),
.B(n_135),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2748),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2827),
.B(n_310),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2796),
.B(n_136),
.Y(n_3028)
);

NOR2xp67_ASAP7_75t_SL g3029 ( 
.A(n_2859),
.B(n_136),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2798),
.B(n_137),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2749),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2763),
.B(n_2776),
.Y(n_3032)
);

AO31x2_ASAP7_75t_L g3033 ( 
.A1(n_2607),
.A2(n_139),
.A3(n_137),
.B(n_138),
.Y(n_3033)
);

OAI21x1_ASAP7_75t_L g3034 ( 
.A1(n_2772),
.A2(n_137),
.B(n_138),
.Y(n_3034)
);

O2A1O1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2811),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2781),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2782),
.Y(n_3037)
);

BUFx3_ASAP7_75t_L g3038 ( 
.A(n_2415),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2804),
.B(n_140),
.Y(n_3039)
);

O2A1O1Ixp5_ASAP7_75t_L g3040 ( 
.A1(n_2459),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_3040)
);

HB1xp67_ASAP7_75t_L g3041 ( 
.A(n_2798),
.Y(n_3041)
);

BUFx3_ASAP7_75t_L g3042 ( 
.A(n_2352),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2511),
.A2(n_141),
.B(n_142),
.Y(n_3043)
);

OAI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2607),
.A2(n_142),
.B(n_143),
.Y(n_3044)
);

OAI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2641),
.A2(n_143),
.B(n_144),
.Y(n_3045)
);

NAND2xp33_ASAP7_75t_SL g3046 ( 
.A(n_2632),
.B(n_144),
.Y(n_3046)
);

AO31x2_ASAP7_75t_L g3047 ( 
.A1(n_2490),
.A2(n_146),
.A3(n_144),
.B(n_145),
.Y(n_3047)
);

A2O1A1Ixp33_ASAP7_75t_L g3048 ( 
.A1(n_2615),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_3048)
);

NOR2xp67_ASAP7_75t_L g3049 ( 
.A(n_2403),
.B(n_2751),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2807),
.B(n_147),
.Y(n_3050)
);

INVx2_ASAP7_75t_SL g3051 ( 
.A(n_2784),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2511),
.A2(n_148),
.B(n_149),
.Y(n_3052)
);

AOI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2551),
.A2(n_148),
.B(n_149),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2551),
.A2(n_148),
.B(n_149),
.Y(n_3054)
);

NOR3xp33_ASAP7_75t_L g3055 ( 
.A(n_2477),
.B(n_150),
.C(n_151),
.Y(n_3055)
);

A2O1A1Ixp33_ASAP7_75t_L g3056 ( 
.A1(n_2663),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_3056)
);

INVx3_ASAP7_75t_L g3057 ( 
.A(n_2403),
.Y(n_3057)
);

CKINVDCx5p33_ASAP7_75t_R g3058 ( 
.A(n_2393),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2814),
.B(n_2816),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2361),
.Y(n_3060)
);

AO31x2_ASAP7_75t_L g3061 ( 
.A1(n_2568),
.A2(n_152),
.A3(n_150),
.B(n_151),
.Y(n_3061)
);

OAI21xp33_ASAP7_75t_L g3062 ( 
.A1(n_2840),
.A2(n_152),
.B(n_153),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2825),
.B(n_153),
.Y(n_3063)
);

AOI21xp5_ASAP7_75t_L g3064 ( 
.A1(n_2505),
.A2(n_153),
.B(n_154),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2826),
.Y(n_3065)
);

OA21x2_ASAP7_75t_L g3066 ( 
.A1(n_2568),
.A2(n_154),
.B(n_155),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2505),
.A2(n_155),
.B(n_156),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2529),
.B(n_155),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2506),
.A2(n_157),
.B(n_158),
.Y(n_3069)
);

OR2x2_ASAP7_75t_L g3070 ( 
.A(n_2855),
.B(n_157),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2855),
.B(n_157),
.Y(n_3071)
);

NOR2xp67_ASAP7_75t_SL g3072 ( 
.A(n_2759),
.B(n_2797),
.Y(n_3072)
);

OAI21x1_ASAP7_75t_L g3073 ( 
.A1(n_2783),
.A2(n_158),
.B(n_159),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2851),
.B(n_158),
.Y(n_3074)
);

OAI21x1_ASAP7_75t_L g3075 ( 
.A1(n_2791),
.A2(n_159),
.B(n_160),
.Y(n_3075)
);

AO31x2_ASAP7_75t_L g3076 ( 
.A1(n_2717),
.A2(n_161),
.A3(n_159),
.B(n_160),
.Y(n_3076)
);

CKINVDCx20_ASAP7_75t_R g3077 ( 
.A(n_2801),
.Y(n_3077)
);

OAI22xp5_ASAP7_75t_L g3078 ( 
.A1(n_2440),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_3078)
);

BUFx12f_ASAP7_75t_L g3079 ( 
.A(n_2785),
.Y(n_3079)
);

OAI22xp5_ASAP7_75t_SL g3080 ( 
.A1(n_2431),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2853),
.B(n_163),
.Y(n_3081)
);

OAI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2668),
.A2(n_2576),
.B(n_2656),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2800),
.Y(n_3083)
);

OAI21x1_ASAP7_75t_L g3084 ( 
.A1(n_2803),
.A2(n_164),
.B(n_165),
.Y(n_3084)
);

OAI21x1_ASAP7_75t_L g3085 ( 
.A1(n_2808),
.A2(n_166),
.B(n_167),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2864),
.B(n_2866),
.Y(n_3086)
);

AND2x2_ASAP7_75t_L g3087 ( 
.A(n_2408),
.B(n_166),
.Y(n_3087)
);

OAI21x1_ASAP7_75t_L g3088 ( 
.A1(n_2812),
.A2(n_167),
.B(n_168),
.Y(n_3088)
);

OAI21x1_ASAP7_75t_L g3089 ( 
.A1(n_2824),
.A2(n_168),
.B(n_169),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_2408),
.B(n_168),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2506),
.A2(n_169),
.B(n_170),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2828),
.Y(n_3092)
);

AO31x2_ASAP7_75t_L g3093 ( 
.A1(n_2717),
.A2(n_171),
.A3(n_169),
.B(n_170),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2751),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2375),
.B(n_170),
.Y(n_3095)
);

INVx5_ASAP7_75t_L g3096 ( 
.A(n_2860),
.Y(n_3096)
);

INVx4_ASAP7_75t_L g3097 ( 
.A(n_2751),
.Y(n_3097)
);

OAI21x1_ASAP7_75t_L g3098 ( 
.A1(n_2841),
.A2(n_171),
.B(n_172),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2858),
.Y(n_3099)
);

OAI21x1_ASAP7_75t_L g3100 ( 
.A1(n_2538),
.A2(n_171),
.B(n_172),
.Y(n_3100)
);

OAI21x1_ASAP7_75t_L g3101 ( 
.A1(n_2617),
.A2(n_172),
.B(n_173),
.Y(n_3101)
);

AOI21xp5_ASAP7_75t_L g3102 ( 
.A1(n_2684),
.A2(n_174),
.B(n_175),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2414),
.B(n_175),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2543),
.B(n_175),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2539),
.A2(n_176),
.B(n_177),
.Y(n_3105)
);

AND3x1_ASAP7_75t_SL g3106 ( 
.A(n_2838),
.B(n_177),
.C(n_178),
.Y(n_3106)
);

AOI21x1_ASAP7_75t_SL g3107 ( 
.A1(n_2576),
.A2(n_178),
.B(n_179),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_SL g3108 ( 
.A(n_2830),
.B(n_311),
.Y(n_3108)
);

AOI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2539),
.A2(n_179),
.B(n_180),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2738),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2545),
.B(n_180),
.Y(n_3111)
);

NOR3xp33_ASAP7_75t_L g3112 ( 
.A(n_2832),
.B(n_181),
.C(n_182),
.Y(n_3112)
);

INVx4_ASAP7_75t_L g3113 ( 
.A(n_2751),
.Y(n_3113)
);

OAI21x1_ASAP7_75t_SL g3114 ( 
.A1(n_2640),
.A2(n_182),
.B(n_183),
.Y(n_3114)
);

AOI21x1_ASAP7_75t_L g3115 ( 
.A1(n_2631),
.A2(n_184),
.B(n_185),
.Y(n_3115)
);

OAI21x1_ASAP7_75t_L g3116 ( 
.A1(n_2617),
.A2(n_2549),
.B(n_2548),
.Y(n_3116)
);

AO31x2_ASAP7_75t_L g3117 ( 
.A1(n_2738),
.A2(n_186),
.A3(n_184),
.B(n_185),
.Y(n_3117)
);

NOR2x1_ASAP7_75t_L g3118 ( 
.A(n_2780),
.B(n_185),
.Y(n_3118)
);

OAI21x1_ASAP7_75t_L g3119 ( 
.A1(n_2562),
.A2(n_186),
.B(n_187),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2637),
.B(n_188),
.Y(n_3120)
);

INVx3_ASAP7_75t_L g3121 ( 
.A(n_2764),
.Y(n_3121)
);

AO31x2_ASAP7_75t_L g3122 ( 
.A1(n_2740),
.A2(n_191),
.A3(n_189),
.B(n_190),
.Y(n_3122)
);

BUFx3_ASAP7_75t_L g3123 ( 
.A(n_2805),
.Y(n_3123)
);

AOI21x1_ASAP7_75t_L g3124 ( 
.A1(n_2440),
.A2(n_189),
.B(n_190),
.Y(n_3124)
);

OAI21x1_ASAP7_75t_L g3125 ( 
.A1(n_2577),
.A2(n_189),
.B(n_190),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2643),
.B(n_191),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_2414),
.B(n_191),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_2755),
.B(n_2873),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2386),
.A2(n_193),
.B(n_194),
.Y(n_3129)
);

OAI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_2740),
.A2(n_2745),
.B1(n_2750),
.B2(n_2743),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2386),
.A2(n_193),
.B(n_194),
.Y(n_3131)
);

CKINVDCx16_ASAP7_75t_R g3132 ( 
.A(n_2862),
.Y(n_3132)
);

OAI21xp5_ASAP7_75t_L g3133 ( 
.A1(n_2658),
.A2(n_193),
.B(n_195),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2645),
.B(n_195),
.Y(n_3134)
);

OAI21x1_ASAP7_75t_L g3135 ( 
.A1(n_2599),
.A2(n_196),
.B(n_197),
.Y(n_3135)
);

OA21x2_ASAP7_75t_L g3136 ( 
.A1(n_2754),
.A2(n_196),
.B(n_197),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2650),
.B(n_2655),
.Y(n_3137)
);

OAI21x1_ASAP7_75t_L g3138 ( 
.A1(n_2612),
.A2(n_196),
.B(n_198),
.Y(n_3138)
);

NOR2xp67_ASAP7_75t_L g3139 ( 
.A(n_2764),
.B(n_199),
.Y(n_3139)
);

AOI21xp5_ASAP7_75t_SL g3140 ( 
.A1(n_2624),
.A2(n_198),
.B(n_199),
.Y(n_3140)
);

OAI21x1_ASAP7_75t_L g3141 ( 
.A1(n_2353),
.A2(n_198),
.B(n_200),
.Y(n_3141)
);

BUFx6f_ASAP7_75t_L g3142 ( 
.A(n_2371),
.Y(n_3142)
);

OAI21x1_ASAP7_75t_SL g3143 ( 
.A1(n_2754),
.A2(n_200),
.B(n_201),
.Y(n_3143)
);

O2A1O1Ixp5_ASAP7_75t_L g3144 ( 
.A1(n_2380),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_3144)
);

OAI22x1_ASAP7_75t_L g3145 ( 
.A1(n_2721),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_3145)
);

AOI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_2390),
.A2(n_202),
.B(n_204),
.Y(n_3146)
);

AOI21xp5_ASAP7_75t_L g3147 ( 
.A1(n_2390),
.A2(n_204),
.B(n_205),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2758),
.Y(n_3148)
);

OA22x2_ASAP7_75t_L g3149 ( 
.A1(n_2544),
.A2(n_2429),
.B1(n_2433),
.B2(n_2419),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2758),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_3150)
);

OAI21x1_ASAP7_75t_L g3151 ( 
.A1(n_2353),
.A2(n_2367),
.B(n_2366),
.Y(n_3151)
);

OAI21x1_ASAP7_75t_L g3152 ( 
.A1(n_2366),
.A2(n_206),
.B(n_208),
.Y(n_3152)
);

BUFx2_ASAP7_75t_L g3153 ( 
.A(n_2351),
.Y(n_3153)
);

OAI21x1_ASAP7_75t_L g3154 ( 
.A1(n_2367),
.A2(n_208),
.B(n_209),
.Y(n_3154)
);

NOR2x1_ASAP7_75t_SL g3155 ( 
.A(n_2764),
.B(n_208),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2371),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2478),
.B(n_209),
.Y(n_3157)
);

OAI21x1_ASAP7_75t_L g3158 ( 
.A1(n_2564),
.A2(n_209),
.B(n_210),
.Y(n_3158)
);

HB1xp67_ASAP7_75t_L g3159 ( 
.A(n_2718),
.Y(n_3159)
);

AO21x1_ASAP7_75t_L g3160 ( 
.A1(n_2741),
.A2(n_314),
.B(n_312),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_2716),
.B(n_211),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_2716),
.B(n_212),
.Y(n_3162)
);

NAND2x1_ASAP7_75t_L g3163 ( 
.A(n_2860),
.B(n_212),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_SL g3164 ( 
.A(n_2466),
.B(n_314),
.Y(n_3164)
);

OAI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_2712),
.A2(n_213),
.B(n_214),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2389),
.Y(n_3166)
);

INVx3_ASAP7_75t_L g3167 ( 
.A(n_2764),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2856),
.B(n_213),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2482),
.B(n_214),
.Y(n_3169)
);

BUFx4_ASAP7_75t_SL g3170 ( 
.A(n_2400),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2485),
.B(n_214),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2730),
.B(n_315),
.Y(n_3172)
);

HB1xp67_ASAP7_75t_L g3173 ( 
.A(n_2734),
.Y(n_3173)
);

OAI21x1_ASAP7_75t_L g3174 ( 
.A1(n_2564),
.A2(n_215),
.B(n_216),
.Y(n_3174)
);

A2O1A1Ixp33_ASAP7_75t_L g3175 ( 
.A1(n_2674),
.A2(n_219),
.B(n_217),
.C(n_218),
.Y(n_3175)
);

NAND2x1_ASAP7_75t_L g3176 ( 
.A(n_2860),
.B(n_217),
.Y(n_3176)
);

AOI221xp5_ASAP7_75t_L g3177 ( 
.A1(n_2434),
.A2(n_220),
.B1(n_217),
.B2(n_218),
.C(n_221),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2399),
.A2(n_218),
.B(n_220),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2451),
.B(n_221),
.Y(n_3179)
);

INVx4_ASAP7_75t_L g3180 ( 
.A(n_2817),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2412),
.Y(n_3181)
);

OAI21x1_ASAP7_75t_L g3182 ( 
.A1(n_2531),
.A2(n_222),
.B(n_223),
.Y(n_3182)
);

NAND3xp33_ASAP7_75t_L g3183 ( 
.A(n_2552),
.B(n_222),
.C(n_223),
.Y(n_3183)
);

BUFx2_ASAP7_75t_L g3184 ( 
.A(n_2767),
.Y(n_3184)
);

OA21x2_ASAP7_75t_L g3185 ( 
.A1(n_2769),
.A2(n_222),
.B(n_223),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2399),
.A2(n_224),
.B(n_225),
.Y(n_3186)
);

OAI21x1_ASAP7_75t_L g3187 ( 
.A1(n_2542),
.A2(n_2514),
.B(n_2513),
.Y(n_3187)
);

INVx1_ASAP7_75t_SL g3188 ( 
.A(n_2768),
.Y(n_3188)
);

BUFx12f_ASAP7_75t_L g3189 ( 
.A(n_2829),
.Y(n_3189)
);

OA21x2_ASAP7_75t_L g3190 ( 
.A1(n_2769),
.A2(n_224),
.B(n_225),
.Y(n_3190)
);

OAI21x1_ASAP7_75t_L g3191 ( 
.A1(n_2644),
.A2(n_2630),
.B(n_2622),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_SL g3192 ( 
.A(n_2404),
.B(n_226),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_2374),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2451),
.B(n_226),
.Y(n_3194)
);

NAND3xp33_ASAP7_75t_SL g3195 ( 
.A(n_2670),
.B(n_226),
.C(n_227),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2856),
.B(n_227),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2567),
.B(n_227),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2422),
.Y(n_3198)
);

NOR2x1_ASAP7_75t_SL g3199 ( 
.A(n_2817),
.B(n_228),
.Y(n_3199)
);

BUFx6f_ASAP7_75t_L g3200 ( 
.A(n_2374),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2778),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2567),
.B(n_228),
.Y(n_3202)
);

INVx3_ASAP7_75t_L g3203 ( 
.A(n_2817),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_2374),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_2407),
.A2(n_229),
.B(n_230),
.Y(n_3205)
);

A2O1A1Ixp33_ASAP7_75t_L g3206 ( 
.A1(n_2674),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2442),
.B(n_229),
.Y(n_3207)
);

AOI22xp5_ASAP7_75t_L g3208 ( 
.A1(n_2821),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3208)
);

NAND2x1p5_ASAP7_75t_L g3209 ( 
.A(n_2813),
.B(n_232),
.Y(n_3209)
);

INVx5_ASAP7_75t_L g3210 ( 
.A(n_2516),
.Y(n_3210)
);

OAI22xp5_ASAP7_75t_L g3211 ( 
.A1(n_2778),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2442),
.B(n_233),
.Y(n_3212)
);

BUFx3_ASAP7_75t_L g3213 ( 
.A(n_2373),
.Y(n_3213)
);

NOR4xp25_ASAP7_75t_L g3214 ( 
.A(n_2854),
.B(n_236),
.C(n_234),
.D(n_235),
.Y(n_3214)
);

OAI21x1_ASAP7_75t_L g3215 ( 
.A1(n_2644),
.A2(n_237),
.B(n_238),
.Y(n_3215)
);

OAI21x1_ASAP7_75t_L g3216 ( 
.A1(n_2779),
.A2(n_237),
.B(n_238),
.Y(n_3216)
);

INVx2_ASAP7_75t_SL g3217 ( 
.A(n_2813),
.Y(n_3217)
);

CKINVDCx5p33_ASAP7_75t_R g3218 ( 
.A(n_2394),
.Y(n_3218)
);

OAI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_2779),
.A2(n_238),
.B(n_239),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2572),
.B(n_239),
.Y(n_3220)
);

OAI21xp33_ASAP7_75t_L g3221 ( 
.A1(n_2844),
.A2(n_240),
.B(n_241),
.Y(n_3221)
);

NAND3xp33_ASAP7_75t_L g3222 ( 
.A(n_2552),
.B(n_240),
.C(n_241),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_2799),
.B(n_240),
.Y(n_3223)
);

OAI21x1_ASAP7_75t_L g3224 ( 
.A1(n_2788),
.A2(n_241),
.B(n_242),
.Y(n_3224)
);

AO31x2_ASAP7_75t_L g3225 ( 
.A1(n_2788),
.A2(n_244),
.A3(n_242),
.B(n_243),
.Y(n_3225)
);

AOI21x1_ASAP7_75t_L g3226 ( 
.A1(n_2679),
.A2(n_243),
.B(n_244),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2524),
.B(n_244),
.Y(n_3227)
);

OR2x6_ASAP7_75t_L g3228 ( 
.A(n_2453),
.B(n_245),
.Y(n_3228)
);

OAI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2806),
.A2(n_246),
.B(n_247),
.Y(n_3229)
);

AO21x1_ASAP7_75t_L g3230 ( 
.A1(n_2818),
.A2(n_316),
.B(n_315),
.Y(n_3230)
);

A2O1A1Ixp33_ASAP7_75t_L g3231 ( 
.A1(n_2608),
.A2(n_248),
.B(n_246),
.C(n_247),
.Y(n_3231)
);

OAI21x1_ASAP7_75t_L g3232 ( 
.A1(n_2806),
.A2(n_247),
.B(n_248),
.Y(n_3232)
);

OAI21x1_ASAP7_75t_L g3233 ( 
.A1(n_2810),
.A2(n_249),
.B(n_250),
.Y(n_3233)
);

OAI21x1_ASAP7_75t_L g3234 ( 
.A1(n_2810),
.A2(n_249),
.B(n_250),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2819),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_2525),
.B(n_249),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_2819),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_3237)
);

BUFx3_ASAP7_75t_L g3238 ( 
.A(n_2382),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2525),
.B(n_251),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_SL g3240 ( 
.A(n_2809),
.B(n_317),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_2439),
.Y(n_3241)
);

AO21x2_ASAP7_75t_L g3242 ( 
.A1(n_2822),
.A2(n_2843),
.B(n_2839),
.Y(n_3242)
);

BUFx12f_ASAP7_75t_L g3243 ( 
.A(n_2823),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2407),
.A2(n_251),
.B(n_253),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2571),
.B(n_253),
.Y(n_3245)
);

OAI21x1_ASAP7_75t_L g3246 ( 
.A1(n_2822),
.A2(n_254),
.B(n_255),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2625),
.B(n_254),
.Y(n_3247)
);

AOI21x1_ASAP7_75t_SL g3248 ( 
.A1(n_2541),
.A2(n_255),
.B(n_256),
.Y(n_3248)
);

OAI21x1_ASAP7_75t_L g3249 ( 
.A1(n_2839),
.A2(n_255),
.B(n_256),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2445),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_2436),
.A2(n_256),
.B(n_257),
.Y(n_3251)
);

INVx2_ASAP7_75t_SL g3252 ( 
.A(n_2823),
.Y(n_3252)
);

AOI21x1_ASAP7_75t_L g3253 ( 
.A1(n_2679),
.A2(n_258),
.B(n_259),
.Y(n_3253)
);

OAI22xp5_ASAP7_75t_L g3254 ( 
.A1(n_2843),
.A2(n_2857),
.B1(n_2861),
.B2(n_2845),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2835),
.B(n_258),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_2842),
.B(n_259),
.Y(n_3256)
);

AO31x2_ASAP7_75t_L g3257 ( 
.A1(n_2845),
.A2(n_2861),
.A3(n_2863),
.B(n_2857),
.Y(n_3257)
);

AOI221x1_ASAP7_75t_L g3258 ( 
.A1(n_2601),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.C(n_263),
.Y(n_3258)
);

BUFx3_ASAP7_75t_L g3259 ( 
.A(n_2363),
.Y(n_3259)
);

AO31x2_ASAP7_75t_L g3260 ( 
.A1(n_2863),
.A2(n_263),
.A3(n_261),
.B(n_262),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_2847),
.B(n_318),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2409),
.B(n_261),
.Y(n_3262)
);

AOI22xp33_ASAP7_75t_L g3263 ( 
.A1(n_2365),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2868),
.Y(n_3264)
);

OAI21x1_ASAP7_75t_SL g3265 ( 
.A1(n_2868),
.A2(n_264),
.B(n_265),
.Y(n_3265)
);

AO31x2_ASAP7_75t_L g3266 ( 
.A1(n_2870),
.A2(n_267),
.A3(n_265),
.B(n_266),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2411),
.B(n_2610),
.Y(n_3267)
);

CKINVDCx5p33_ASAP7_75t_R g3268 ( 
.A(n_2410),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_2398),
.B(n_265),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2870),
.Y(n_3270)
);

OAI21xp33_ASAP7_75t_L g3271 ( 
.A1(n_2626),
.A2(n_266),
.B(n_267),
.Y(n_3271)
);

AOI22xp5_ASAP7_75t_L g3272 ( 
.A1(n_2815),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_2436),
.A2(n_268),
.B(n_269),
.Y(n_3273)
);

NOR2xp67_ASAP7_75t_L g3274 ( 
.A(n_2817),
.B(n_270),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2388),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2629),
.B(n_269),
.Y(n_3276)
);

OAI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_2449),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2638),
.B(n_271),
.Y(n_3278)
);

OAI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_2694),
.A2(n_272),
.B(n_273),
.Y(n_3279)
);

AO31x2_ASAP7_75t_L g3280 ( 
.A1(n_2541),
.A2(n_275),
.A3(n_273),
.B(n_274),
.Y(n_3280)
);

BUFx2_ASAP7_75t_L g3281 ( 
.A(n_2391),
.Y(n_3281)
);

AOI22xp5_ASAP7_75t_L g3282 ( 
.A1(n_2815),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_3282)
);

AOI21xp33_ASAP7_75t_L g3283 ( 
.A1(n_2547),
.A2(n_274),
.B(n_275),
.Y(n_3283)
);

AND2x6_ASAP7_75t_L g3284 ( 
.A(n_2534),
.B(n_276),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_2449),
.A2(n_276),
.B(n_277),
.Y(n_3285)
);

NAND3x1_ASAP7_75t_L g3286 ( 
.A(n_2777),
.B(n_276),
.C(n_277),
.Y(n_3286)
);

OAI22xp5_ASAP7_75t_L g3287 ( 
.A1(n_2626),
.A2(n_2628),
.B1(n_2679),
.B2(n_2675),
.Y(n_3287)
);

AOI21x1_ASAP7_75t_L g3288 ( 
.A1(n_2834),
.A2(n_277),
.B(n_278),
.Y(n_3288)
);

OAI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_2681),
.A2(n_278),
.B(n_279),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_2495),
.B(n_278),
.Y(n_3290)
);

OR2x2_ASAP7_75t_L g3291 ( 
.A(n_2455),
.B(n_279),
.Y(n_3291)
);

NOR2xp33_ASAP7_75t_L g3292 ( 
.A(n_2540),
.B(n_280),
.Y(n_3292)
);

OAI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_2681),
.A2(n_280),
.B(n_281),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2646),
.B(n_281),
.Y(n_3294)
);

OAI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_2693),
.A2(n_2566),
.B(n_2454),
.Y(n_3295)
);

OAI21x1_ASAP7_75t_L g3296 ( 
.A1(n_2421),
.A2(n_281),
.B(n_282),
.Y(n_3296)
);

OAI21x1_ASAP7_75t_L g3297 ( 
.A1(n_2421),
.A2(n_282),
.B(n_283),
.Y(n_3297)
);

OAI21x1_ASAP7_75t_L g3298 ( 
.A1(n_2503),
.A2(n_283),
.B(n_284),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2405),
.Y(n_3299)
);

INVx1_ASAP7_75t_SL g3300 ( 
.A(n_2516),
.Y(n_3300)
);

OAI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_2628),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_2392),
.A2(n_284),
.B(n_285),
.Y(n_3302)
);

OAI21x1_ASAP7_75t_L g3303 ( 
.A1(n_2503),
.A2(n_285),
.B(n_286),
.Y(n_3303)
);

BUFx6f_ASAP7_75t_L g3304 ( 
.A(n_2392),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_SL g3305 ( 
.A(n_2706),
.B(n_318),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2406),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2676),
.B(n_286),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2515),
.B(n_287),
.Y(n_3308)
);

INVxp67_ASAP7_75t_L g3309 ( 
.A(n_2417),
.Y(n_3309)
);

AO31x2_ASAP7_75t_L g3310 ( 
.A1(n_2454),
.A2(n_289),
.A3(n_287),
.B(n_288),
.Y(n_3310)
);

OAI21x1_ASAP7_75t_L g3311 ( 
.A1(n_2733),
.A2(n_2753),
.B(n_2742),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_2495),
.B(n_287),
.Y(n_3312)
);

OAI21x1_ASAP7_75t_L g3313 ( 
.A1(n_2733),
.A2(n_288),
.B(n_289),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2517),
.B(n_289),
.Y(n_3314)
);

AO21x1_ASAP7_75t_L g3315 ( 
.A1(n_2700),
.A2(n_320),
.B(n_319),
.Y(n_3315)
);

NOR2xp67_ASAP7_75t_L g3316 ( 
.A(n_2820),
.B(n_291),
.Y(n_3316)
);

AOI211x1_ASAP7_75t_L g3317 ( 
.A1(n_2584),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2606),
.B(n_290),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2533),
.B(n_290),
.Y(n_3319)
);

AOI21xp33_ASAP7_75t_L g3320 ( 
.A1(n_2473),
.A2(n_291),
.B(n_292),
.Y(n_3320)
);

OAI21x1_ASAP7_75t_L g3321 ( 
.A1(n_2742),
.A2(n_293),
.B(n_294),
.Y(n_3321)
);

AND3x2_ASAP7_75t_L g3322 ( 
.A(n_2713),
.B(n_2770),
.C(n_2723),
.Y(n_3322)
);

CKINVDCx5p33_ASAP7_75t_R g3323 ( 
.A(n_2852),
.Y(n_3323)
);

INVx5_ASAP7_75t_L g3324 ( 
.A(n_2516),
.Y(n_3324)
);

OAI21x1_ASAP7_75t_L g3325 ( 
.A1(n_2753),
.A2(n_293),
.B(n_294),
.Y(n_3325)
);

AO31x2_ASAP7_75t_L g3326 ( 
.A1(n_2687),
.A2(n_296),
.A3(n_293),
.B(n_295),
.Y(n_3326)
);

OAI21x1_ASAP7_75t_L g3327 ( 
.A1(n_2789),
.A2(n_295),
.B(n_296),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2392),
.A2(n_295),
.B(n_296),
.Y(n_3328)
);

AND2x2_ASAP7_75t_SL g3329 ( 
.A(n_2453),
.B(n_297),
.Y(n_3329)
);

OAI21x1_ASAP7_75t_L g3330 ( 
.A1(n_2789),
.A2(n_297),
.B(n_298),
.Y(n_3330)
);

CKINVDCx5p33_ASAP7_75t_R g3331 ( 
.A(n_2468),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2533),
.B(n_298),
.Y(n_3332)
);

OAI21x1_ASAP7_75t_L g3333 ( 
.A1(n_2837),
.A2(n_298),
.B(n_299),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2647),
.B(n_2654),
.Y(n_3334)
);

BUFx3_ASAP7_75t_L g3335 ( 
.A(n_3243),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_3170),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3151),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2949),
.Y(n_3338)
);

OAI21x1_ASAP7_75t_L g3339 ( 
.A1(n_2901),
.A2(n_2865),
.B(n_2837),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_2889),
.B(n_2493),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2917),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_2957),
.Y(n_3342)
);

INVx4_ASAP7_75t_SL g3343 ( 
.A(n_2905),
.Y(n_3343)
);

CKINVDCx20_ASAP7_75t_R g3344 ( 
.A(n_2920),
.Y(n_3344)
);

CKINVDCx6p67_ASAP7_75t_R g3345 ( 
.A(n_2892),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_2978),
.B(n_2526),
.Y(n_3346)
);

OAI21xp33_ASAP7_75t_SL g3347 ( 
.A1(n_3272),
.A2(n_2836),
.B(n_2354),
.Y(n_3347)
);

NOR4xp25_ASAP7_75t_L g3348 ( 
.A(n_3286),
.B(n_2765),
.C(n_2786),
.D(n_2522),
.Y(n_3348)
);

OAI21x1_ASAP7_75t_L g3349 ( 
.A1(n_3191),
.A2(n_2865),
.B(n_2642),
.Y(n_3349)
);

O2A1O1Ixp33_ASAP7_75t_SL g3350 ( 
.A1(n_2993),
.A2(n_2498),
.B(n_2486),
.C(n_2635),
.Y(n_3350)
);

CKINVDCx6p67_ASAP7_75t_R g3351 ( 
.A(n_2899),
.Y(n_3351)
);

BUFx5_ASAP7_75t_L g3352 ( 
.A(n_2891),
.Y(n_3352)
);

CKINVDCx5p33_ASAP7_75t_R g3353 ( 
.A(n_2942),
.Y(n_3353)
);

OAI21x1_ASAP7_75t_L g3354 ( 
.A1(n_3116),
.A2(n_2510),
.B(n_2530),
.Y(n_3354)
);

OAI21x1_ASAP7_75t_L g3355 ( 
.A1(n_3248),
.A2(n_2555),
.B(n_2530),
.Y(n_3355)
);

CKINVDCx20_ASAP7_75t_R g3356 ( 
.A(n_3077),
.Y(n_3356)
);

BUFx3_ASAP7_75t_L g3357 ( 
.A(n_3038),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_2949),
.Y(n_3358)
);

OAI21x1_ASAP7_75t_L g3359 ( 
.A1(n_3311),
.A2(n_2555),
.B(n_2460),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2949),
.Y(n_3360)
);

OAI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_2878),
.A2(n_2475),
.B1(n_2675),
.B2(n_2627),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_2991),
.B(n_2651),
.Y(n_3362)
);

AO21x1_ASAP7_75t_L g3363 ( 
.A1(n_2878),
.A2(n_2723),
.B(n_2713),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_L g3364 ( 
.A(n_2926),
.B(n_2653),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_2879),
.A2(n_2707),
.B1(n_2673),
.B2(n_2618),
.Y(n_3365)
);

AND2x4_ASAP7_75t_L g3366 ( 
.A(n_3096),
.B(n_2437),
.Y(n_3366)
);

INVx1_ASAP7_75t_SL g3367 ( 
.A(n_3213),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_3128),
.B(n_2910),
.Y(n_3368)
);

INVxp67_ASAP7_75t_L g3369 ( 
.A(n_3153),
.Y(n_3369)
);

OAI222xp33_ASAP7_75t_L g3370 ( 
.A1(n_3272),
.A2(n_2491),
.B1(n_2479),
.B2(n_2441),
.C1(n_2831),
.C2(n_2770),
.Y(n_3370)
);

OAI21x1_ASAP7_75t_L g3371 ( 
.A1(n_3107),
.A2(n_2471),
.B(n_2458),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3257),
.Y(n_3372)
);

OR2x6_ASAP7_75t_L g3373 ( 
.A(n_2940),
.B(n_2964),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3157),
.B(n_2831),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_3322),
.B(n_2596),
.Y(n_3375)
);

AOI21xp33_ASAP7_75t_L g3376 ( 
.A1(n_3130),
.A2(n_2678),
.B(n_2635),
.Y(n_3376)
);

AO31x2_ASAP7_75t_L g3377 ( 
.A1(n_3130),
.A2(n_2687),
.A3(n_2424),
.B(n_2432),
.Y(n_3377)
);

BUFx3_ASAP7_75t_L g3378 ( 
.A(n_3042),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3257),
.Y(n_3379)
);

OAI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3254),
.A2(n_2372),
.B(n_2507),
.Y(n_3380)
);

INVx4_ASAP7_75t_R g3381 ( 
.A(n_2888),
.Y(n_3381)
);

AO32x2_ASAP7_75t_L g3382 ( 
.A1(n_2884),
.A2(n_2491),
.A3(n_2479),
.B1(n_2665),
.B2(n_2582),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_2927),
.B(n_2526),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3137),
.B(n_2428),
.Y(n_3384)
);

OAI21x1_ASAP7_75t_L g3385 ( 
.A1(n_3017),
.A2(n_2476),
.B(n_2662),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_2972),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3267),
.B(n_2430),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2880),
.B(n_2443),
.Y(n_3388)
);

O2A1O1Ixp33_ASAP7_75t_SL g3389 ( 
.A1(n_3163),
.A2(n_2498),
.B(n_2417),
.C(n_2462),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_3005),
.B(n_2833),
.Y(n_3390)
);

OAI21x1_ASAP7_75t_L g3391 ( 
.A1(n_2918),
.A2(n_2457),
.B(n_2446),
.Y(n_3391)
);

OR2x6_ASAP7_75t_L g3392 ( 
.A(n_2940),
.B(n_2833),
.Y(n_3392)
);

OR2x6_ASAP7_75t_L g3393 ( 
.A(n_2940),
.B(n_2846),
.Y(n_3393)
);

INVx3_ASAP7_75t_L g3394 ( 
.A(n_3016),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_3291),
.B(n_2621),
.Y(n_3395)
);

INVx2_ASAP7_75t_SL g3396 ( 
.A(n_2891),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3257),
.Y(n_3397)
);

OAI21x1_ASAP7_75t_L g3398 ( 
.A1(n_3187),
.A2(n_2463),
.B(n_2692),
.Y(n_3398)
);

AND2x4_ASAP7_75t_L g3399 ( 
.A(n_3096),
.B(n_2437),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_SL g3400 ( 
.A1(n_3329),
.A2(n_2846),
.B1(n_2462),
.B2(n_2707),
.Y(n_3400)
);

INVx1_ASAP7_75t_SL g3401 ( 
.A(n_3238),
.Y(n_3401)
);

OR2x2_ASAP7_75t_L g3402 ( 
.A(n_2985),
.B(n_2427),
.Y(n_3402)
);

BUFx6f_ASAP7_75t_SL g3403 ( 
.A(n_2964),
.Y(n_3403)
);

BUFx2_ASAP7_75t_L g3404 ( 
.A(n_2928),
.Y(n_3404)
);

OAI21x1_ASAP7_75t_L g3405 ( 
.A1(n_2874),
.A2(n_2369),
.B(n_2696),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3141),
.Y(n_3406)
);

OAI21x1_ASAP7_75t_L g3407 ( 
.A1(n_2998),
.A2(n_2369),
.B(n_2696),
.Y(n_3407)
);

OAI21x1_ASAP7_75t_L g3408 ( 
.A1(n_2976),
.A2(n_2369),
.B(n_2698),
.Y(n_3408)
);

HB1xp67_ASAP7_75t_L g3409 ( 
.A(n_2939),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3152),
.Y(n_3410)
);

AO21x2_ASAP7_75t_L g3411 ( 
.A1(n_2925),
.A2(n_2581),
.B(n_2732),
.Y(n_3411)
);

AND2x4_ASAP7_75t_L g3412 ( 
.A(n_3096),
.B(n_2437),
.Y(n_3412)
);

OA21x2_ASAP7_75t_L g3413 ( 
.A1(n_2994),
.A2(n_2581),
.B(n_2536),
.Y(n_3413)
);

BUFx12f_ASAP7_75t_L g3414 ( 
.A(n_2990),
.Y(n_3414)
);

AOI221xp5_ASAP7_75t_L g3415 ( 
.A1(n_3214),
.A2(n_2909),
.B1(n_2952),
.B2(n_2884),
.C(n_3254),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3110),
.B(n_2481),
.Y(n_3416)
);

OR2x6_ASAP7_75t_L g3417 ( 
.A(n_2964),
.B(n_2416),
.Y(n_3417)
);

AOI21xp33_ASAP7_75t_SL g3418 ( 
.A1(n_3132),
.A2(n_2565),
.B(n_2574),
.Y(n_3418)
);

OAI21x1_ASAP7_75t_L g3419 ( 
.A1(n_2877),
.A2(n_2369),
.B(n_2705),
.Y(n_3419)
);

AND2x2_ASAP7_75t_L g3420 ( 
.A(n_2961),
.B(n_2427),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3154),
.Y(n_3421)
);

BUFx2_ASAP7_75t_L g3422 ( 
.A(n_2928),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_2982),
.Y(n_3423)
);

OA21x2_ASAP7_75t_L g3424 ( 
.A1(n_2994),
.A2(n_2536),
.B(n_2618),
.Y(n_3424)
);

OA21x2_ASAP7_75t_L g3425 ( 
.A1(n_3082),
.A2(n_2673),
.B(n_2710),
.Y(n_3425)
);

AND2x4_ASAP7_75t_L g3426 ( 
.A(n_3049),
.B(n_2420),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_2879),
.B(n_2420),
.Y(n_3427)
);

AOI22xp5_ASAP7_75t_L g3428 ( 
.A1(n_3046),
.A2(n_2909),
.B1(n_3287),
.B2(n_2999),
.Y(n_3428)
);

OAI21x1_ASAP7_75t_L g3429 ( 
.A1(n_2903),
.A2(n_2369),
.B(n_2496),
.Y(n_3429)
);

OAI21x1_ASAP7_75t_L g3430 ( 
.A1(n_2912),
.A2(n_2499),
.B(n_2497),
.Y(n_3430)
);

NOR2xp67_ASAP7_75t_L g3431 ( 
.A(n_3217),
.B(n_2512),
.Y(n_3431)
);

OAI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3040),
.A2(n_2527),
.B(n_2583),
.Y(n_3432)
);

AND2x2_ASAP7_75t_L g3433 ( 
.A(n_3013),
.B(n_2450),
.Y(n_3433)
);

OAI21x1_ASAP7_75t_L g3434 ( 
.A1(n_2890),
.A2(n_2501),
.B(n_2426),
.Y(n_3434)
);

CKINVDCx5p33_ASAP7_75t_R g3435 ( 
.A(n_3019),
.Y(n_3435)
);

OAI21x1_ASAP7_75t_L g3436 ( 
.A1(n_2898),
.A2(n_2426),
.B(n_2402),
.Y(n_3436)
);

OAI21xp33_ASAP7_75t_SL g3437 ( 
.A1(n_3282),
.A2(n_3139),
.B(n_2988),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_3188),
.B(n_2546),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3242),
.Y(n_3439)
);

BUFx2_ASAP7_75t_L g3440 ( 
.A(n_3281),
.Y(n_3440)
);

INVx3_ASAP7_75t_L g3441 ( 
.A(n_3016),
.Y(n_3441)
);

AOI22xp33_ASAP7_75t_L g3442 ( 
.A1(n_3287),
.A2(n_2452),
.B1(n_2450),
.B2(n_2588),
.Y(n_3442)
);

OAI21x1_ASAP7_75t_L g3443 ( 
.A1(n_3119),
.A2(n_2472),
.B(n_2402),
.Y(n_3443)
);

CKINVDCx20_ASAP7_75t_R g3444 ( 
.A(n_3218),
.Y(n_3444)
);

INVx1_ASAP7_75t_SL g3445 ( 
.A(n_3188),
.Y(n_3445)
);

OAI21x1_ASAP7_75t_L g3446 ( 
.A1(n_3125),
.A2(n_3138),
.B(n_3135),
.Y(n_3446)
);

INVx3_ASAP7_75t_L g3447 ( 
.A(n_3097),
.Y(n_3447)
);

OAI21x1_ASAP7_75t_L g3448 ( 
.A1(n_3182),
.A2(n_2474),
.B(n_2472),
.Y(n_3448)
);

OAI22xp5_ASAP7_75t_L g3449 ( 
.A1(n_3228),
.A2(n_2732),
.B1(n_2775),
.B2(n_2737),
.Y(n_3449)
);

NAND2x1p5_ASAP7_75t_L g3450 ( 
.A(n_3049),
.B(n_2820),
.Y(n_3450)
);

AO31x2_ASAP7_75t_L g3451 ( 
.A1(n_2911),
.A2(n_2709),
.A3(n_2521),
.B(n_2671),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3242),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3148),
.B(n_2557),
.Y(n_3453)
);

NOR2xp67_ASAP7_75t_L g3454 ( 
.A(n_3252),
.B(n_2570),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_L g3455 ( 
.A(n_2908),
.B(n_2598),
.Y(n_3455)
);

OAI21x1_ASAP7_75t_L g3456 ( 
.A1(n_2944),
.A2(n_2519),
.B(n_2474),
.Y(n_3456)
);

NAND2x1p5_ASAP7_75t_L g3457 ( 
.A(n_3072),
.B(n_2820),
.Y(n_3457)
);

OAI22x1_ASAP7_75t_L g3458 ( 
.A1(n_3282),
.A2(n_2452),
.B1(n_2387),
.B2(n_2420),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3192),
.A2(n_2520),
.B(n_2519),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3192),
.A2(n_2520),
.B(n_2519),
.Y(n_3460)
);

OAI21x1_ASAP7_75t_L g3461 ( 
.A1(n_2951),
.A2(n_2719),
.B(n_2520),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2904),
.Y(n_3462)
);

BUFx3_ASAP7_75t_L g3463 ( 
.A(n_3060),
.Y(n_3463)
);

AND2x2_ASAP7_75t_L g3464 ( 
.A(n_3028),
.B(n_2737),
.Y(n_3464)
);

OAI21x1_ASAP7_75t_L g3465 ( 
.A1(n_2981),
.A2(n_2735),
.B(n_2719),
.Y(n_3465)
);

OAI222xp33_ASAP7_75t_L g3466 ( 
.A1(n_3228),
.A2(n_2537),
.B1(n_2420),
.B2(n_2757),
.C1(n_2623),
.C2(n_2401),
.Y(n_3466)
);

OAI21x1_ASAP7_75t_L g3467 ( 
.A1(n_2992),
.A2(n_2795),
.B(n_2735),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_2987),
.Y(n_3468)
);

BUFx2_ASAP7_75t_L g3469 ( 
.A(n_3184),
.Y(n_3469)
);

CKINVDCx6p67_ASAP7_75t_R g3470 ( 
.A(n_3123),
.Y(n_3470)
);

BUFx2_ASAP7_75t_SL g3471 ( 
.A(n_2886),
.Y(n_3471)
);

AOI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_3195),
.A2(n_2605),
.B1(n_2652),
.B2(n_2711),
.Y(n_3472)
);

BUFx2_ASAP7_75t_L g3473 ( 
.A(n_3097),
.Y(n_3473)
);

OAI21x1_ASAP7_75t_L g3474 ( 
.A1(n_3006),
.A2(n_2869),
.B(n_2795),
.Y(n_3474)
);

HB1xp67_ASAP7_75t_L g3475 ( 
.A(n_2956),
.Y(n_3475)
);

OAI21x1_ASAP7_75t_L g3476 ( 
.A1(n_3008),
.A2(n_2871),
.B(n_2869),
.Y(n_3476)
);

BUFx8_ASAP7_75t_L g3477 ( 
.A(n_3079),
.Y(n_3477)
);

INVx3_ASAP7_75t_SL g3478 ( 
.A(n_3058),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_2915),
.Y(n_3479)
);

OAI21xp33_ASAP7_75t_L g3480 ( 
.A1(n_2923),
.A2(n_2793),
.B(n_2775),
.Y(n_3480)
);

OAI21x1_ASAP7_75t_L g3481 ( 
.A1(n_2953),
.A2(n_2872),
.B(n_2871),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3201),
.B(n_3235),
.Y(n_3482)
);

BUFx3_ASAP7_75t_L g3483 ( 
.A(n_3259),
.Y(n_3483)
);

OR2x2_ASAP7_75t_L g3484 ( 
.A(n_2985),
.B(n_2467),
.Y(n_3484)
);

AO21x2_ASAP7_75t_L g3485 ( 
.A1(n_2921),
.A2(n_2793),
.B(n_2583),
.Y(n_3485)
);

OAI21x1_ASAP7_75t_L g3486 ( 
.A1(n_2965),
.A2(n_2872),
.B(n_2871),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3036),
.Y(n_3487)
);

OAI21x1_ASAP7_75t_L g3488 ( 
.A1(n_2971),
.A2(n_2872),
.B(n_2516),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3068),
.B(n_2689),
.Y(n_3489)
);

OAI21x1_ASAP7_75t_L g3490 ( 
.A1(n_3024),
.A2(n_2597),
.B(n_2487),
.Y(n_3490)
);

OAI21x1_ASAP7_75t_L g3491 ( 
.A1(n_3034),
.A2(n_2597),
.B(n_2660),
.Y(n_3491)
);

INVx1_ASAP7_75t_SL g3492 ( 
.A(n_3331),
.Y(n_3492)
);

OA21x2_ASAP7_75t_L g3493 ( 
.A1(n_3216),
.A2(n_2563),
.B(n_2554),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_3210),
.B(n_3324),
.Y(n_3494)
);

BUFx6f_ASAP7_75t_L g3495 ( 
.A(n_2979),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_3083),
.Y(n_3496)
);

INVx2_ASAP7_75t_SL g3497 ( 
.A(n_2922),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_2937),
.Y(n_3498)
);

OAI21x1_ASAP7_75t_L g3499 ( 
.A1(n_3073),
.A2(n_2597),
.B(n_2660),
.Y(n_3499)
);

NAND2x1p5_ASAP7_75t_L g3500 ( 
.A(n_3113),
.B(n_2820),
.Y(n_3500)
);

AOI21xp5_ASAP7_75t_L g3501 ( 
.A1(n_3295),
.A2(n_2660),
.B(n_2404),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3264),
.B(n_2616),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_2966),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3103),
.A2(n_2594),
.B1(n_2602),
.B2(n_2591),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3270),
.B(n_2387),
.Y(n_3505)
);

OA21x2_ASAP7_75t_L g3506 ( 
.A1(n_3224),
.A2(n_2563),
.B(n_2554),
.Y(n_3506)
);

OR2x2_ASAP7_75t_L g3507 ( 
.A(n_3015),
.B(n_2509),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_2969),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3000),
.Y(n_3509)
);

OAI21x1_ASAP7_75t_L g3510 ( 
.A1(n_3075),
.A2(n_2597),
.B(n_2660),
.Y(n_3510)
);

NOR2xp33_ASAP7_75t_L g3511 ( 
.A(n_3164),
.B(n_2589),
.Y(n_3511)
);

O2A1O1Ixp33_ASAP7_75t_SL g3512 ( 
.A1(n_3176),
.A2(n_2537),
.B(n_2867),
.C(n_2483),
.Y(n_3512)
);

AND2x4_ASAP7_75t_L g3513 ( 
.A(n_3210),
.B(n_2537),
.Y(n_3513)
);

AO21x2_ASAP7_75t_L g3514 ( 
.A1(n_2907),
.A2(n_2483),
.B(n_2484),
.Y(n_3514)
);

AND2x4_ASAP7_75t_L g3515 ( 
.A(n_3210),
.B(n_2537),
.Y(n_3515)
);

OA21x2_ASAP7_75t_L g3516 ( 
.A1(n_3232),
.A2(n_2669),
.B(n_2589),
.Y(n_3516)
);

BUFx5_ASAP7_75t_L g3517 ( 
.A(n_3284),
.Y(n_3517)
);

OR2x6_ASAP7_75t_L g3518 ( 
.A(n_3228),
.B(n_2416),
.Y(n_3518)
);

INVx3_ASAP7_75t_L g3519 ( 
.A(n_3113),
.Y(n_3519)
);

AO21x2_ASAP7_75t_L g3520 ( 
.A1(n_2907),
.A2(n_2504),
.B(n_2484),
.Y(n_3520)
);

OAI21x1_ASAP7_75t_L g3521 ( 
.A1(n_3084),
.A2(n_2620),
.B(n_2586),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3092),
.Y(n_3522)
);

INVxp67_ASAP7_75t_SL g3523 ( 
.A(n_3041),
.Y(n_3523)
);

OAI21x1_ASAP7_75t_L g3524 ( 
.A1(n_3085),
.A2(n_2620),
.B(n_2586),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3022),
.Y(n_3525)
);

OAI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_2999),
.A2(n_2919),
.B1(n_3209),
.B2(n_3301),
.Y(n_3526)
);

OAI21x1_ASAP7_75t_L g3527 ( 
.A1(n_3088),
.A2(n_2586),
.B(n_2633),
.Y(n_3527)
);

NAND2x1p5_ASAP7_75t_L g3528 ( 
.A(n_3180),
.B(n_2867),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3026),
.B(n_2504),
.Y(n_3529)
);

INVx3_ASAP7_75t_L g3530 ( 
.A(n_3180),
.Y(n_3530)
);

AOI21xp33_ASAP7_75t_SL g3531 ( 
.A1(n_3149),
.A2(n_2623),
.B(n_299),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3031),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3099),
.Y(n_3533)
);

BUFx12f_ASAP7_75t_L g3534 ( 
.A(n_3189),
.Y(n_3534)
);

OAI21x1_ASAP7_75t_L g3535 ( 
.A1(n_3089),
.A2(n_2586),
.B(n_2633),
.Y(n_3535)
);

OAI21x1_ASAP7_75t_L g3536 ( 
.A1(n_3098),
.A2(n_2633),
.B(n_2603),
.Y(n_3536)
);

AND2x4_ASAP7_75t_L g3537 ( 
.A(n_3324),
.B(n_2867),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3324),
.B(n_2867),
.Y(n_3538)
);

O2A1O1Ixp33_ASAP7_75t_L g3539 ( 
.A1(n_3175),
.A2(n_2623),
.B(n_2444),
.C(n_2465),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3037),
.Y(n_3540)
);

INVx2_ASAP7_75t_L g3541 ( 
.A(n_2893),
.Y(n_3541)
);

OAI22xp5_ASAP7_75t_L g3542 ( 
.A1(n_2967),
.A2(n_2701),
.B1(n_2690),
.B2(n_2699),
.Y(n_3542)
);

OAI21x1_ASAP7_75t_L g3543 ( 
.A1(n_3233),
.A2(n_2603),
.B(n_2521),
.Y(n_3543)
);

AOI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3127),
.A2(n_2695),
.B1(n_2699),
.B2(n_2690),
.Y(n_3544)
);

AND2x4_ASAP7_75t_L g3545 ( 
.A(n_3057),
.B(n_2532),
.Y(n_3545)
);

OAI21x1_ASAP7_75t_L g3546 ( 
.A1(n_3234),
.A2(n_3249),
.B(n_3246),
.Y(n_3546)
);

AOI332xp33_ASAP7_75t_L g3547 ( 
.A1(n_3065),
.A2(n_304),
.A3(n_303),
.B1(n_299),
.B2(n_301),
.B3(n_300),
.C1(n_302),
.C2(n_319),
.Y(n_3547)
);

INVx4_ASAP7_75t_L g3548 ( 
.A(n_3057),
.Y(n_3548)
);

INVx4_ASAP7_75t_L g3549 ( 
.A(n_3094),
.Y(n_3549)
);

NAND3xp33_ASAP7_75t_L g3550 ( 
.A(n_2967),
.B(n_2699),
.C(n_2695),
.Y(n_3550)
);

NOR2xp33_ASAP7_75t_L g3551 ( 
.A(n_3159),
.B(n_2438),
.Y(n_3551)
);

NAND2xp33_ASAP7_75t_L g3552 ( 
.A(n_3284),
.B(n_2532),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3334),
.B(n_2701),
.Y(n_3553)
);

A2O1A1Ixp33_ASAP7_75t_L g3554 ( 
.A1(n_2923),
.A2(n_2695),
.B(n_2636),
.C(n_2672),
.Y(n_3554)
);

A2O1A1Ixp33_ASAP7_75t_SL g3555 ( 
.A1(n_2996),
.A2(n_3029),
.B(n_3045),
.C(n_2924),
.Y(n_3555)
);

BUFx3_ASAP7_75t_L g3556 ( 
.A(n_3003),
.Y(n_3556)
);

BUFx8_ASAP7_75t_SL g3557 ( 
.A(n_3323),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3136),
.Y(n_3558)
);

AOI22xp33_ASAP7_75t_L g3559 ( 
.A1(n_3055),
.A2(n_2636),
.B1(n_2672),
.B2(n_2532),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_2896),
.Y(n_3560)
);

CKINVDCx20_ASAP7_75t_R g3561 ( 
.A(n_3268),
.Y(n_3561)
);

OAI21x1_ASAP7_75t_L g3562 ( 
.A1(n_3010),
.A2(n_2672),
.B(n_2636),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3030),
.B(n_300),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3166),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3094),
.B(n_300),
.Y(n_3565)
);

AOI21xp33_ASAP7_75t_L g3566 ( 
.A1(n_3319),
.A2(n_302),
.B(n_303),
.Y(n_3566)
);

OAI21x1_ASAP7_75t_L g3567 ( 
.A1(n_2938),
.A2(n_304),
.B(n_303),
.Y(n_3567)
);

OAI21x1_ASAP7_75t_L g3568 ( 
.A1(n_3296),
.A2(n_304),
.B(n_302),
.Y(n_3568)
);

OAI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_2986),
.A2(n_322),
.B(n_324),
.Y(n_3569)
);

OAI221xp5_ASAP7_75t_L g3570 ( 
.A1(n_3295),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.C(n_327),
.Y(n_3570)
);

OAI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_2936),
.A2(n_325),
.B(n_327),
.Y(n_3571)
);

INVx1_ASAP7_75t_SL g3572 ( 
.A(n_3051),
.Y(n_3572)
);

AOI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_3112),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_3573)
);

AO21x2_ASAP7_75t_L g3574 ( 
.A1(n_3143),
.A2(n_331),
.B(n_333),
.Y(n_3574)
);

OAI21x1_ASAP7_75t_L g3575 ( 
.A1(n_3297),
.A2(n_333),
.B(n_334),
.Y(n_3575)
);

OR2x2_ASAP7_75t_L g3576 ( 
.A(n_3070),
.B(n_334),
.Y(n_3576)
);

OAI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_2936),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_3577)
);

AOI22xp5_ASAP7_75t_L g3578 ( 
.A1(n_3292),
.A2(n_339),
.B1(n_336),
.B2(n_338),
.Y(n_3578)
);

OAI221xp5_ASAP7_75t_L g3579 ( 
.A1(n_3271),
.A2(n_341),
.B1(n_338),
.B2(n_339),
.C(n_342),
.Y(n_3579)
);

OAI21x1_ASAP7_75t_L g3580 ( 
.A1(n_3298),
.A2(n_341),
.B(n_342),
.Y(n_3580)
);

OAI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_2963),
.A2(n_343),
.B(n_344),
.Y(n_3581)
);

A2O1A1Ixp33_ASAP7_75t_L g3582 ( 
.A1(n_2906),
.A2(n_3062),
.B(n_2931),
.C(n_3221),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3181),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3136),
.Y(n_3584)
);

BUFx2_ASAP7_75t_L g3585 ( 
.A(n_3121),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3185),
.Y(n_3586)
);

AO31x2_ASAP7_75t_L g3587 ( 
.A1(n_2945),
.A2(n_346),
.A3(n_344),
.B(n_345),
.Y(n_3587)
);

OAI21x1_ASAP7_75t_L g3588 ( 
.A1(n_3303),
.A2(n_345),
.B(n_346),
.Y(n_3588)
);

AO31x2_ASAP7_75t_L g3589 ( 
.A1(n_3160),
.A2(n_349),
.A3(n_347),
.B(n_348),
.Y(n_3589)
);

OAI21x1_ASAP7_75t_L g3590 ( 
.A1(n_3313),
.A2(n_347),
.B(n_348),
.Y(n_3590)
);

AND2x4_ASAP7_75t_L g3591 ( 
.A(n_3121),
.B(n_3167),
.Y(n_3591)
);

OAI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_2963),
.A2(n_349),
.B(n_350),
.Y(n_3592)
);

OR2x6_ASAP7_75t_L g3593 ( 
.A(n_2897),
.B(n_351),
.Y(n_3593)
);

INVx4_ASAP7_75t_L g3594 ( 
.A(n_3167),
.Y(n_3594)
);

INVx6_ASAP7_75t_L g3595 ( 
.A(n_2897),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3185),
.Y(n_3596)
);

O2A1O1Ixp33_ASAP7_75t_L g3597 ( 
.A1(n_3206),
.A2(n_3172),
.B(n_3261),
.C(n_3240),
.Y(n_3597)
);

OAI21x1_ASAP7_75t_L g3598 ( 
.A1(n_3321),
.A2(n_351),
.B(n_352),
.Y(n_3598)
);

INVx4_ASAP7_75t_L g3599 ( 
.A(n_3203),
.Y(n_3599)
);

AO21x2_ASAP7_75t_L g3600 ( 
.A1(n_3165),
.A2(n_353),
.B(n_355),
.Y(n_3600)
);

BUFx6f_ASAP7_75t_L g3601 ( 
.A(n_2979),
.Y(n_3601)
);

OAI21x1_ASAP7_75t_L g3602 ( 
.A1(n_3325),
.A2(n_355),
.B(n_356),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3190),
.Y(n_3603)
);

OAI21x1_ASAP7_75t_L g3604 ( 
.A1(n_3327),
.A2(n_356),
.B(n_357),
.Y(n_3604)
);

OAI21x1_ASAP7_75t_L g3605 ( 
.A1(n_3330),
.A2(n_358),
.B(n_359),
.Y(n_3605)
);

BUFx3_ASAP7_75t_L g3606 ( 
.A(n_3173),
.Y(n_3606)
);

O2A1O1Ixp33_ASAP7_75t_L g3607 ( 
.A1(n_3301),
.A2(n_362),
.B(n_358),
.C(n_360),
.Y(n_3607)
);

INVx3_ASAP7_75t_L g3608 ( 
.A(n_3203),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_2970),
.B(n_363),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3190),
.Y(n_3610)
);

OR2x2_ASAP7_75t_L g3611 ( 
.A(n_3071),
.B(n_363),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3280),
.Y(n_3612)
);

INVxp67_ASAP7_75t_L g3613 ( 
.A(n_3087),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3280),
.Y(n_3614)
);

AO21x2_ASAP7_75t_L g3615 ( 
.A1(n_3265),
.A2(n_364),
.B(n_365),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_3140),
.A2(n_365),
.B(n_366),
.Y(n_3616)
);

AOI221xp5_ASAP7_75t_SL g3617 ( 
.A1(n_2946),
.A2(n_370),
.B1(n_367),
.B2(n_368),
.C(n_371),
.Y(n_3617)
);

INVx2_ASAP7_75t_SL g3618 ( 
.A(n_2975),
.Y(n_3618)
);

INVx1_ASAP7_75t_SL g3619 ( 
.A(n_3090),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3280),
.Y(n_3620)
);

OAI21x1_ASAP7_75t_L g3621 ( 
.A1(n_3333),
.A2(n_367),
.B(n_368),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3309),
.B(n_371),
.Y(n_3622)
);

OAI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3183),
.A2(n_372),
.B(n_373),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3215),
.Y(n_3624)
);

INVx8_ASAP7_75t_L g3625 ( 
.A(n_2975),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3124),
.A2(n_374),
.B(n_375),
.Y(n_3626)
);

OR2x2_ASAP7_75t_L g3627 ( 
.A(n_3236),
.B(n_375),
.Y(n_3627)
);

BUFx6f_ASAP7_75t_L g3628 ( 
.A(n_2979),
.Y(n_3628)
);

OAI21x1_ASAP7_75t_L g3629 ( 
.A1(n_3115),
.A2(n_376),
.B(n_377),
.Y(n_3629)
);

AOI21xp5_ASAP7_75t_L g3630 ( 
.A1(n_3300),
.A2(n_376),
.B(n_377),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3047),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_SL g3632 ( 
.A1(n_3155),
.A2(n_378),
.B(n_379),
.Y(n_3632)
);

NAND3xp33_ASAP7_75t_L g3633 ( 
.A(n_3317),
.B(n_3222),
.C(n_3183),
.Y(n_3633)
);

OAI21x1_ASAP7_75t_L g3634 ( 
.A1(n_3018),
.A2(n_378),
.B(n_379),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3032),
.B(n_380),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3059),
.B(n_844),
.Y(n_3636)
);

AND2x4_ASAP7_75t_L g3637 ( 
.A(n_2988),
.B(n_381),
.Y(n_3637)
);

AO21x2_ASAP7_75t_L g3638 ( 
.A1(n_3165),
.A2(n_381),
.B(n_382),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3047),
.Y(n_3639)
);

AO31x2_ASAP7_75t_L g3640 ( 
.A1(n_3315),
.A2(n_384),
.A3(n_382),
.B(n_383),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3198),
.Y(n_3641)
);

OAI21x1_ASAP7_75t_L g3642 ( 
.A1(n_3100),
.A2(n_384),
.B(n_386),
.Y(n_3642)
);

OAI21x1_ASAP7_75t_SL g3643 ( 
.A1(n_3199),
.A2(n_386),
.B(n_387),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3241),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3250),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3095),
.B(n_387),
.Y(n_3646)
);

OAI21x1_ASAP7_75t_L g3647 ( 
.A1(n_2902),
.A2(n_389),
.B(n_390),
.Y(n_3647)
);

OAI21x1_ASAP7_75t_L g3648 ( 
.A1(n_3101),
.A2(n_389),
.B(n_390),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_3275),
.Y(n_3649)
);

AND2x4_ASAP7_75t_L g3650 ( 
.A(n_3139),
.B(n_391),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3290),
.B(n_391),
.Y(n_3651)
);

INVx3_ASAP7_75t_L g3652 ( 
.A(n_3142),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3047),
.Y(n_3653)
);

OAI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3158),
.A2(n_394),
.B(n_395),
.Y(n_3654)
);

AND2x4_ASAP7_75t_L g3655 ( 
.A(n_3274),
.B(n_395),
.Y(n_3655)
);

OA21x2_ASAP7_75t_L g3656 ( 
.A1(n_2913),
.A2(n_396),
.B(n_397),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3086),
.B(n_843),
.Y(n_3657)
);

OAI21x1_ASAP7_75t_L g3658 ( 
.A1(n_3174),
.A2(n_3011),
.B(n_3014),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3299),
.Y(n_3659)
);

NOR2xp67_ASAP7_75t_L g3660 ( 
.A(n_2959),
.B(n_396),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3306),
.Y(n_3661)
);

OAI21x1_ASAP7_75t_SL g3662 ( 
.A1(n_3009),
.A2(n_3114),
.B(n_3226),
.Y(n_3662)
);

AO21x2_ASAP7_75t_L g3663 ( 
.A1(n_2913),
.A2(n_397),
.B(n_398),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3007),
.Y(n_3664)
);

AOI31xp67_ASAP7_75t_L g3665 ( 
.A1(n_2881),
.A2(n_2883),
.A3(n_3332),
.B(n_3194),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3007),
.Y(n_3666)
);

CKINVDCx20_ASAP7_75t_R g3667 ( 
.A(n_3106),
.Y(n_3667)
);

A2O1A1Ixp33_ASAP7_75t_L g3668 ( 
.A1(n_2906),
.A2(n_400),
.B(n_398),
.C(n_399),
.Y(n_3668)
);

OAI21x1_ASAP7_75t_L g3669 ( 
.A1(n_3288),
.A2(n_2882),
.B(n_2934),
.Y(n_3669)
);

OAI21x1_ASAP7_75t_L g3670 ( 
.A1(n_2882),
.A2(n_399),
.B(n_400),
.Y(n_3670)
);

OAI22xp33_ASAP7_75t_L g3671 ( 
.A1(n_3222),
.A2(n_404),
.B1(n_401),
.B2(n_402),
.Y(n_3671)
);

BUFx12f_ASAP7_75t_L g3672 ( 
.A(n_3284),
.Y(n_3672)
);

NOR2xp67_ASAP7_75t_L g3673 ( 
.A(n_3318),
.B(n_405),
.Y(n_3673)
);

HB1xp67_ASAP7_75t_L g3674 ( 
.A(n_3312),
.Y(n_3674)
);

AO21x2_ASAP7_75t_L g3675 ( 
.A1(n_2924),
.A2(n_405),
.B(n_406),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_3007),
.Y(n_3676)
);

INVx1_ASAP7_75t_SL g3677 ( 
.A(n_3223),
.Y(n_3677)
);

CKINVDCx20_ASAP7_75t_R g3678 ( 
.A(n_3080),
.Y(n_3678)
);

OAI21x1_ASAP7_75t_L g3679 ( 
.A1(n_2895),
.A2(n_406),
.B(n_407),
.Y(n_3679)
);

OAI21x1_ASAP7_75t_SL g3680 ( 
.A1(n_3253),
.A2(n_407),
.B(n_408),
.Y(n_3680)
);

AND2x4_ASAP7_75t_L g3681 ( 
.A(n_3274),
.B(n_409),
.Y(n_3681)
);

CKINVDCx16_ASAP7_75t_R g3682 ( 
.A(n_3080),
.Y(n_3682)
);

INVx1_ASAP7_75t_SL g3683 ( 
.A(n_3255),
.Y(n_3683)
);

NOR2x1_ASAP7_75t_R g3684 ( 
.A(n_3305),
.B(n_2989),
.Y(n_3684)
);

AO21x1_ASAP7_75t_L g3685 ( 
.A1(n_2914),
.A2(n_409),
.B(n_410),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3269),
.B(n_410),
.Y(n_3686)
);

OAI21x1_ASAP7_75t_L g3687 ( 
.A1(n_2900),
.A2(n_411),
.B(n_412),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3326),
.Y(n_3688)
);

OR2x2_ASAP7_75t_L g3689 ( 
.A(n_3239),
.B(n_411),
.Y(n_3689)
);

OA21x2_ASAP7_75t_L g3690 ( 
.A1(n_3219),
.A2(n_413),
.B(n_414),
.Y(n_3690)
);

AOI21xp5_ASAP7_75t_SL g3691 ( 
.A1(n_2914),
.A2(n_3062),
.B(n_3150),
.Y(n_3691)
);

AO21x2_ASAP7_75t_L g3692 ( 
.A1(n_3219),
.A2(n_414),
.B(n_415),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_3221),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_3256),
.Y(n_3694)
);

AND2x2_ASAP7_75t_L g3695 ( 
.A(n_3161),
.B(n_418),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3025),
.Y(n_3696)
);

OAI22xp5_ASAP7_75t_L g3697 ( 
.A1(n_3208),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_3697)
);

INVx6_ASAP7_75t_L g3698 ( 
.A(n_3284),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3326),
.Y(n_3699)
);

AOI21xp5_ASAP7_75t_L g3700 ( 
.A1(n_3300),
.A2(n_420),
.B(n_422),
.Y(n_3700)
);

O2A1O1Ixp33_ASAP7_75t_SL g3701 ( 
.A1(n_2947),
.A2(n_424),
.B(n_422),
.C(n_423),
.Y(n_3701)
);

NAND3xp33_ASAP7_75t_L g3702 ( 
.A(n_3317),
.B(n_423),
.C(n_424),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3220),
.B(n_843),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_SL g3704 ( 
.A(n_3316),
.B(n_425),
.Y(n_3704)
);

OAI22xp5_ASAP7_75t_L g3705 ( 
.A1(n_3208),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_3705)
);

AND2x4_ASAP7_75t_L g3706 ( 
.A(n_3316),
.B(n_426),
.Y(n_3706)
);

OAI21x1_ASAP7_75t_L g3707 ( 
.A1(n_2973),
.A2(n_427),
.B(n_429),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3227),
.B(n_842),
.Y(n_3708)
);

AO21x2_ASAP7_75t_L g3709 ( 
.A1(n_3229),
.A2(n_842),
.B(n_429),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_L g3710 ( 
.A(n_3278),
.B(n_3294),
.Y(n_3710)
);

OAI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3025),
.A2(n_430),
.B(n_431),
.Y(n_3711)
);

OA21x2_ASAP7_75t_L g3712 ( 
.A1(n_3229),
.A2(n_431),
.B(n_432),
.Y(n_3712)
);

OAI21x1_ASAP7_75t_L g3713 ( 
.A1(n_3302),
.A2(n_432),
.B(n_433),
.Y(n_3713)
);

OAI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3277),
.A2(n_435),
.B1(n_433),
.B2(n_434),
.Y(n_3714)
);

OAI21xp5_ASAP7_75t_L g3715 ( 
.A1(n_3144),
.A2(n_434),
.B(n_435),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3326),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3066),
.Y(n_3717)
);

AND2x4_ASAP7_75t_L g3718 ( 
.A(n_3279),
.B(n_436),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_L g3719 ( 
.A1(n_3283),
.A2(n_440),
.B1(n_437),
.B2(n_438),
.Y(n_3719)
);

AO21x2_ASAP7_75t_L g3720 ( 
.A1(n_3133),
.A2(n_841),
.B(n_437),
.Y(n_3720)
);

OA21x2_ASAP7_75t_L g3721 ( 
.A1(n_3045),
.A2(n_2968),
.B(n_2958),
.Y(n_3721)
);

CKINVDCx12_ASAP7_75t_R g3722 ( 
.A(n_3162),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_3307),
.B(n_440),
.Y(n_3723)
);

AOI31xp33_ASAP7_75t_L g3724 ( 
.A1(n_3277),
.A2(n_443),
.A3(n_441),
.B(n_442),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3033),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_2930),
.Y(n_3726)
);

OAI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_3279),
.A2(n_444),
.B1(n_441),
.B2(n_443),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_SL g3728 ( 
.A(n_2995),
.B(n_445),
.Y(n_3728)
);

OAI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_2941),
.A2(n_447),
.B(n_448),
.Y(n_3729)
);

HB1xp67_ASAP7_75t_L g3730 ( 
.A(n_3409),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3338),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3338),
.Y(n_3732)
);

BUFx4f_ASAP7_75t_SL g3733 ( 
.A(n_3477),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3682),
.B(n_3340),
.Y(n_3734)
);

NAND2x1_ASAP7_75t_L g3735 ( 
.A(n_3698),
.B(n_3118),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3462),
.Y(n_3736)
);

AOI221x1_ASAP7_75t_L g3737 ( 
.A1(n_3531),
.A2(n_3145),
.B1(n_3002),
.B2(n_3023),
.C(n_2954),
.Y(n_3737)
);

AOI21xp5_ASAP7_75t_L g3738 ( 
.A1(n_3501),
.A2(n_2887),
.B(n_3200),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3341),
.Y(n_3739)
);

OAI22xp5_ASAP7_75t_L g3740 ( 
.A1(n_3400),
.A2(n_3150),
.B1(n_3237),
.B2(n_3211),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3482),
.B(n_3214),
.Y(n_3741)
);

BUFx4f_ASAP7_75t_SL g3742 ( 
.A(n_3477),
.Y(n_3742)
);

AND2x6_ASAP7_75t_L g3743 ( 
.A(n_3366),
.B(n_3142),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3649),
.B(n_3168),
.Y(n_3744)
);

AND2x4_ASAP7_75t_L g3745 ( 
.A(n_3548),
.B(n_3142),
.Y(n_3745)
);

AOI22xp5_ASAP7_75t_L g3746 ( 
.A1(n_3361),
.A2(n_3004),
.B1(n_3108),
.B2(n_3027),
.Y(n_3746)
);

OAI22xp33_ASAP7_75t_L g3747 ( 
.A1(n_3724),
.A2(n_3258),
.B1(n_3211),
.B2(n_3237),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3342),
.Y(n_3748)
);

AOI221xp5_ASAP7_75t_SL g3749 ( 
.A1(n_3526),
.A2(n_2962),
.B1(n_3263),
.B2(n_3078),
.C(n_3177),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3661),
.B(n_3196),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3386),
.Y(n_3751)
);

AOI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3363),
.A2(n_3078),
.B1(n_2948),
.B2(n_2954),
.Y(n_3752)
);

OAI22xp5_ASAP7_75t_L g3753 ( 
.A1(n_3428),
.A2(n_2933),
.B1(n_3023),
.B2(n_3002),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3462),
.Y(n_3754)
);

INVx4_ASAP7_75t_L g3755 ( 
.A(n_3625),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3479),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3479),
.Y(n_3757)
);

OAI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3365),
.A2(n_3593),
.B1(n_3698),
.B2(n_3518),
.Y(n_3758)
);

OAI221xp5_ASAP7_75t_L g3759 ( 
.A1(n_3380),
.A2(n_3056),
.B1(n_3048),
.B2(n_3283),
.C(n_3133),
.Y(n_3759)
);

AND2x4_ASAP7_75t_L g3760 ( 
.A(n_3548),
.B(n_3156),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3423),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3498),
.B(n_3061),
.Y(n_3762)
);

INVx3_ASAP7_75t_L g3763 ( 
.A(n_3450),
.Y(n_3763)
);

INVx6_ASAP7_75t_L g3764 ( 
.A(n_3534),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3498),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3468),
.Y(n_3766)
);

OAI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3347),
.A2(n_3102),
.B(n_2950),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3503),
.B(n_3061),
.Y(n_3768)
);

AND2x4_ASAP7_75t_L g3769 ( 
.A(n_3549),
.B(n_3156),
.Y(n_3769)
);

CKINVDCx6p67_ASAP7_75t_R g3770 ( 
.A(n_3335),
.Y(n_3770)
);

INVx4_ASAP7_75t_L g3771 ( 
.A(n_3625),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3503),
.Y(n_3772)
);

AOI21xp33_ASAP7_75t_L g3773 ( 
.A1(n_3555),
.A2(n_3597),
.B(n_3539),
.Y(n_3773)
);

OAI22xp33_ASAP7_75t_L g3774 ( 
.A1(n_3593),
.A2(n_2933),
.B1(n_3293),
.B2(n_3289),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3487),
.Y(n_3775)
);

OAI22xp33_ASAP7_75t_SL g3776 ( 
.A1(n_3595),
.A2(n_2943),
.B1(n_2916),
.B2(n_3197),
.Y(n_3776)
);

AOI221xp5_ASAP7_75t_SL g3777 ( 
.A1(n_3678),
.A2(n_3449),
.B1(n_3415),
.B2(n_3667),
.C(n_3455),
.Y(n_3777)
);

AOI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3403),
.A2(n_3230),
.B1(n_3320),
.B2(n_2958),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3368),
.B(n_3202),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3403),
.A2(n_2968),
.B1(n_2885),
.B2(n_2995),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3374),
.B(n_3289),
.Y(n_3781)
);

INVx3_ASAP7_75t_L g3782 ( 
.A(n_3549),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3508),
.Y(n_3783)
);

AOI22xp33_ASAP7_75t_L g3784 ( 
.A1(n_3718),
.A2(n_3001),
.B1(n_3044),
.B2(n_3293),
.Y(n_3784)
);

INVx3_ASAP7_75t_L g3785 ( 
.A(n_3594),
.Y(n_3785)
);

BUFx4f_ASAP7_75t_L g3786 ( 
.A(n_3417),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3563),
.B(n_3001),
.Y(n_3787)
);

AOI22xp33_ASAP7_75t_L g3788 ( 
.A1(n_3718),
.A2(n_3044),
.B1(n_3212),
.B2(n_3207),
.Y(n_3788)
);

BUFx5_ASAP7_75t_L g3789 ( 
.A(n_3426),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3496),
.Y(n_3790)
);

CKINVDCx11_ASAP7_75t_R g3791 ( 
.A(n_3356),
.Y(n_3791)
);

NAND3xp33_ASAP7_75t_SL g3792 ( 
.A(n_3547),
.B(n_3231),
.C(n_3035),
.Y(n_3792)
);

OAI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3518),
.A2(n_3179),
.B1(n_3245),
.B2(n_3147),
.Y(n_3793)
);

AND2x4_ASAP7_75t_L g3794 ( 
.A(n_3594),
.B(n_3193),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3509),
.B(n_3033),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3686),
.B(n_3076),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3509),
.Y(n_3797)
);

NAND2xp33_ASAP7_75t_SL g3798 ( 
.A(n_3458),
.B(n_3193),
.Y(n_3798)
);

NAND2x1p5_ASAP7_75t_L g3799 ( 
.A(n_3336),
.B(n_3193),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3651),
.B(n_3076),
.Y(n_3800)
);

NAND2x1_ASAP7_75t_L g3801 ( 
.A(n_3599),
.B(n_3200),
.Y(n_3801)
);

NAND3xp33_ASAP7_75t_L g3802 ( 
.A(n_3550),
.B(n_3109),
.C(n_3105),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3420),
.B(n_3076),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3525),
.Y(n_3804)
);

NAND3xp33_ASAP7_75t_SL g3805 ( 
.A(n_3344),
.B(n_2974),
.C(n_3146),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3525),
.B(n_3033),
.Y(n_3806)
);

INVxp67_ASAP7_75t_L g3807 ( 
.A(n_3440),
.Y(n_3807)
);

BUFx6f_ASAP7_75t_L g3808 ( 
.A(n_3473),
.Y(n_3808)
);

OAI21x1_ASAP7_75t_L g3809 ( 
.A1(n_3669),
.A2(n_3328),
.B(n_3091),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3672),
.A2(n_3012),
.B1(n_3043),
.B2(n_2977),
.Y(n_3810)
);

INVx2_ASAP7_75t_SL g3811 ( 
.A(n_3381),
.Y(n_3811)
);

OR2x2_ASAP7_75t_L g3812 ( 
.A(n_3523),
.B(n_3093),
.Y(n_3812)
);

AOI22xp33_ASAP7_75t_L g3813 ( 
.A1(n_3480),
.A2(n_3053),
.B1(n_3054),
.B2(n_3052),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_SL g3814 ( 
.A(n_3517),
.B(n_3200),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3520),
.A2(n_3067),
.B1(n_3064),
.B2(n_3069),
.Y(n_3815)
);

NOR2xp33_ASAP7_75t_L g3816 ( 
.A(n_3553),
.B(n_3364),
.Y(n_3816)
);

AOI22xp33_ASAP7_75t_SL g3817 ( 
.A1(n_3595),
.A2(n_3186),
.B1(n_3205),
.B2(n_3178),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3532),
.Y(n_3818)
);

HB1xp67_ASAP7_75t_L g3819 ( 
.A(n_3475),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3532),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3540),
.B(n_3093),
.Y(n_3821)
);

BUFx2_ASAP7_75t_L g3822 ( 
.A(n_3404),
.Y(n_3822)
);

CKINVDCx8_ASAP7_75t_R g3823 ( 
.A(n_3471),
.Y(n_3823)
);

INVx2_ASAP7_75t_SL g3824 ( 
.A(n_3357),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3433),
.B(n_3093),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3540),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3520),
.A2(n_3251),
.B1(n_3273),
.B2(n_3244),
.Y(n_3827)
);

AND2x2_ASAP7_75t_L g3828 ( 
.A(n_3674),
.B(n_3117),
.Y(n_3828)
);

INVx3_ASAP7_75t_L g3829 ( 
.A(n_3599),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3659),
.Y(n_3830)
);

OAI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3417),
.A2(n_3285),
.B1(n_2876),
.B2(n_2875),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3619),
.B(n_3117),
.Y(n_3832)
);

HB1xp67_ASAP7_75t_L g3833 ( 
.A(n_3402),
.Y(n_3833)
);

BUFx6f_ASAP7_75t_L g3834 ( 
.A(n_3426),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3659),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3522),
.Y(n_3836)
);

AOI22xp33_ASAP7_75t_L g3837 ( 
.A1(n_3464),
.A2(n_3247),
.B1(n_3131),
.B2(n_3129),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3533),
.Y(n_3838)
);

INVx2_ASAP7_75t_SL g3839 ( 
.A(n_3345),
.Y(n_3839)
);

NAND2xp33_ASAP7_75t_SL g3840 ( 
.A(n_3422),
.B(n_3204),
.Y(n_3840)
);

BUFx2_ASAP7_75t_L g3841 ( 
.A(n_3352),
.Y(n_3841)
);

INVx1_ASAP7_75t_SL g3842 ( 
.A(n_3351),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3392),
.A2(n_2983),
.B1(n_2997),
.B2(n_2980),
.Y(n_3843)
);

HB1xp67_ASAP7_75t_L g3844 ( 
.A(n_3469),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3677),
.B(n_3117),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3564),
.Y(n_3846)
);

OAI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_3373),
.A2(n_3020),
.B1(n_2929),
.B2(n_2932),
.Y(n_3847)
);

INVx2_ASAP7_75t_SL g3848 ( 
.A(n_3470),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3541),
.Y(n_3849)
);

AOI22xp33_ASAP7_75t_L g3850 ( 
.A1(n_3514),
.A2(n_2935),
.B1(n_2955),
.B2(n_2894),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3646),
.B(n_3683),
.Y(n_3851)
);

OAI22xp5_ASAP7_75t_L g3852 ( 
.A1(n_3392),
.A2(n_2960),
.B1(n_3126),
.B2(n_3120),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3583),
.Y(n_3853)
);

NAND3xp33_ASAP7_75t_SL g3854 ( 
.A(n_3348),
.B(n_3276),
.C(n_3134),
.Y(n_3854)
);

OAI221xp5_ASAP7_75t_L g3855 ( 
.A1(n_3472),
.A2(n_3021),
.B1(n_3063),
.B2(n_3050),
.C(n_3039),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3641),
.Y(n_3856)
);

NOR2xp33_ASAP7_75t_L g3857 ( 
.A(n_3497),
.B(n_3074),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3695),
.B(n_3122),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3358),
.Y(n_3859)
);

AOI22xp33_ASAP7_75t_SL g3860 ( 
.A1(n_3517),
.A2(n_3304),
.B1(n_3204),
.B2(n_3081),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3613),
.B(n_3611),
.Y(n_3861)
);

INVx2_ASAP7_75t_SL g3862 ( 
.A(n_3378),
.Y(n_3862)
);

CKINVDCx11_ASAP7_75t_R g3863 ( 
.A(n_3414),
.Y(n_3863)
);

AOI22xp33_ASAP7_75t_L g3864 ( 
.A1(n_3514),
.A2(n_3262),
.B1(n_3104),
.B2(n_3111),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_SL g3865 ( 
.A1(n_3517),
.A2(n_3304),
.B1(n_3204),
.B2(n_3171),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3346),
.B(n_3122),
.Y(n_3866)
);

AOI22xp33_ASAP7_75t_L g3867 ( 
.A1(n_3376),
.A2(n_3169),
.B1(n_3314),
.B2(n_3308),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_3557),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3383),
.B(n_3122),
.Y(n_3869)
);

AND2x2_ASAP7_75t_L g3870 ( 
.A(n_3396),
.B(n_3225),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3560),
.Y(n_3871)
);

AO22x2_ASAP7_75t_L g3872 ( 
.A1(n_3372),
.A2(n_3225),
.B1(n_3266),
.B2(n_3260),
.Y(n_3872)
);

AOI21xp33_ASAP7_75t_L g3873 ( 
.A1(n_3432),
.A2(n_3304),
.B(n_2984),
.Y(n_3873)
);

AND2x2_ASAP7_75t_SL g3874 ( 
.A(n_3552),
.B(n_3225),
.Y(n_3874)
);

AOI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3710),
.A2(n_3310),
.B1(n_3260),
.B2(n_3266),
.Y(n_3875)
);

AND2x2_ASAP7_75t_L g3876 ( 
.A(n_3565),
.B(n_3260),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3565),
.B(n_3266),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3644),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3390),
.B(n_3694),
.Y(n_3879)
);

BUFx6f_ASAP7_75t_L g3880 ( 
.A(n_3495),
.Y(n_3880)
);

BUFx3_ASAP7_75t_L g3881 ( 
.A(n_3463),
.Y(n_3881)
);

OAI211xp5_ASAP7_75t_L g3882 ( 
.A1(n_3660),
.A2(n_3310),
.B(n_2930),
.C(n_2984),
.Y(n_3882)
);

OAI221xp5_ASAP7_75t_L g3883 ( 
.A1(n_3442),
.A2(n_3310),
.B1(n_2930),
.B2(n_2984),
.C(n_451),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3645),
.Y(n_3884)
);

AOI221xp5_ASAP7_75t_L g3885 ( 
.A1(n_3691),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.C(n_452),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3453),
.Y(n_3886)
);

AOI22xp33_ASAP7_75t_L g3887 ( 
.A1(n_3485),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_3887)
);

AOI221xp5_ASAP7_75t_L g3888 ( 
.A1(n_3727),
.A2(n_3384),
.B1(n_3714),
.B2(n_3566),
.C(n_3387),
.Y(n_3888)
);

OR2x2_ASAP7_75t_L g3889 ( 
.A(n_3445),
.B(n_453),
.Y(n_3889)
);

AO31x2_ASAP7_75t_L g3890 ( 
.A1(n_3726),
.A2(n_456),
.A3(n_454),
.B(n_455),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3502),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3358),
.Y(n_3892)
);

AND2x4_ASAP7_75t_L g3893 ( 
.A(n_3394),
.B(n_456),
.Y(n_3893)
);

BUFx3_ASAP7_75t_L g3894 ( 
.A(n_3483),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3606),
.B(n_457),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_L g3896 ( 
.A1(n_3485),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_3896)
);

AND2x4_ASAP7_75t_L g3897 ( 
.A(n_3394),
.B(n_458),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3618),
.B(n_841),
.Y(n_3898)
);

OR2x2_ASAP7_75t_L g3899 ( 
.A(n_3507),
.B(n_459),
.Y(n_3899)
);

BUFx3_ASAP7_75t_L g3900 ( 
.A(n_3556),
.Y(n_3900)
);

AOI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_3489),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3352),
.B(n_461),
.Y(n_3902)
);

AOI22xp5_ASAP7_75t_SL g3903 ( 
.A1(n_3375),
.A2(n_466),
.B1(n_463),
.B2(n_465),
.Y(n_3903)
);

CKINVDCx5p33_ASAP7_75t_R g3904 ( 
.A(n_3353),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3352),
.Y(n_3905)
);

OAI221xp5_ASAP7_75t_L g3906 ( 
.A1(n_3504),
.A2(n_470),
.B1(n_466),
.B2(n_468),
.C(n_471),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3430),
.Y(n_3907)
);

OR2x6_ASAP7_75t_L g3908 ( 
.A(n_3373),
.B(n_468),
.Y(n_3908)
);

INVx3_ASAP7_75t_L g3909 ( 
.A(n_3537),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_3352),
.Y(n_3910)
);

INVx2_ASAP7_75t_L g3911 ( 
.A(n_3352),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3393),
.A2(n_473),
.B1(n_470),
.B2(n_472),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3438),
.B(n_3367),
.Y(n_3913)
);

AND2x4_ASAP7_75t_L g3914 ( 
.A(n_3441),
.B(n_472),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3401),
.B(n_473),
.Y(n_3915)
);

NAND2xp33_ASAP7_75t_R g3916 ( 
.A(n_3393),
.B(n_474),
.Y(n_3916)
);

AOI221xp5_ASAP7_75t_SL g3917 ( 
.A1(n_3505),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.C(n_477),
.Y(n_3917)
);

AND2x4_ASAP7_75t_L g3918 ( 
.A(n_3441),
.B(n_475),
.Y(n_3918)
);

OAI22x1_ASAP7_75t_L g3919 ( 
.A1(n_3369),
.A2(n_479),
.B1(n_476),
.B2(n_478),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3484),
.Y(n_3920)
);

OAI22xp5_ASAP7_75t_L g3921 ( 
.A1(n_3693),
.A2(n_482),
.B1(n_480),
.B2(n_481),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3388),
.B(n_480),
.Y(n_3922)
);

HB1xp67_ASAP7_75t_L g3923 ( 
.A(n_3585),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3702),
.Y(n_3924)
);

AOI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3685),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_3925)
);

OAI22xp5_ASAP7_75t_L g3926 ( 
.A1(n_3570),
.A2(n_3668),
.B1(n_3633),
.B2(n_3582),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3558),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3416),
.B(n_483),
.Y(n_3928)
);

OAI21x1_ASAP7_75t_L g3929 ( 
.A1(n_3465),
.A2(n_484),
.B(n_485),
.Y(n_3929)
);

INVx1_ASAP7_75t_SL g3930 ( 
.A(n_3572),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3576),
.B(n_3529),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3558),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3511),
.B(n_486),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3584),
.Y(n_3934)
);

OR2x2_ASAP7_75t_L g3935 ( 
.A(n_3635),
.B(n_487),
.Y(n_3935)
);

NAND3xp33_ASAP7_75t_SL g3936 ( 
.A(n_3457),
.B(n_487),
.C(n_488),
.Y(n_3936)
);

AND2x4_ASAP7_75t_SL g3937 ( 
.A(n_3447),
.B(n_489),
.Y(n_3937)
);

NAND2xp33_ASAP7_75t_SL g3938 ( 
.A(n_3447),
.B(n_490),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_SL g3939 ( 
.A1(n_3517),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_SL g3940 ( 
.A1(n_3571),
.A2(n_491),
.B(n_492),
.Y(n_3940)
);

AOI21xp33_ASAP7_75t_L g3941 ( 
.A1(n_3684),
.A2(n_3542),
.B(n_3411),
.Y(n_3941)
);

INVx2_ASAP7_75t_L g3942 ( 
.A(n_3584),
.Y(n_3942)
);

BUFx4_ASAP7_75t_SL g3943 ( 
.A(n_3444),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3622),
.B(n_840),
.Y(n_3944)
);

NOR2xp33_ASAP7_75t_L g3945 ( 
.A(n_3395),
.B(n_3492),
.Y(n_3945)
);

INVx2_ASAP7_75t_SL g3946 ( 
.A(n_3343),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3551),
.B(n_840),
.Y(n_3947)
);

AND2x4_ASAP7_75t_L g3948 ( 
.A(n_3519),
.B(n_495),
.Y(n_3948)
);

OAI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3581),
.A2(n_495),
.B(n_497),
.Y(n_3949)
);

NAND3xp33_ASAP7_75t_SL g3950 ( 
.A(n_3418),
.B(n_498),
.C(n_500),
.Y(n_3950)
);

AOI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3413),
.A2(n_502),
.B1(n_498),
.B2(n_501),
.Y(n_3951)
);

AOI221xp5_ASAP7_75t_SL g3952 ( 
.A1(n_3370),
.A2(n_503),
.B1(n_501),
.B2(n_502),
.C(n_504),
.Y(n_3952)
);

AOI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3413),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_3953)
);

INVx4_ASAP7_75t_L g3954 ( 
.A(n_3343),
.Y(n_3954)
);

BUFx10_ASAP7_75t_L g3955 ( 
.A(n_3435),
.Y(n_3955)
);

AOI22xp33_ASAP7_75t_L g3956 ( 
.A1(n_3697),
.A2(n_3705),
.B1(n_3721),
.B2(n_3517),
.Y(n_3956)
);

BUFx2_ASAP7_75t_L g3957 ( 
.A(n_3519),
.Y(n_3957)
);

AOI22xp33_ASAP7_75t_L g3958 ( 
.A1(n_3721),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3958)
);

INVx2_ASAP7_75t_SL g3959 ( 
.A(n_3591),
.Y(n_3959)
);

NOR2xp33_ASAP7_75t_L g3960 ( 
.A(n_3362),
.B(n_506),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3723),
.A2(n_3424),
.B1(n_3427),
.B2(n_3411),
.Y(n_3961)
);

AOI22xp33_ASAP7_75t_L g3962 ( 
.A1(n_3424),
.A2(n_510),
.B1(n_507),
.B2(n_509),
.Y(n_3962)
);

OR2x6_ASAP7_75t_L g3963 ( 
.A(n_3454),
.B(n_3431),
.Y(n_3963)
);

HB1xp67_ASAP7_75t_L g3964 ( 
.A(n_3591),
.Y(n_3964)
);

AO21x2_ASAP7_75t_L g3965 ( 
.A1(n_3662),
.A2(n_509),
.B(n_510),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3586),
.Y(n_3966)
);

AOI22xp33_ASAP7_75t_L g3967 ( 
.A1(n_3728),
.A2(n_513),
.B1(n_511),
.B2(n_512),
.Y(n_3967)
);

OAI22xp5_ASAP7_75t_L g3968 ( 
.A1(n_3573),
.A2(n_514),
.B1(n_511),
.B2(n_513),
.Y(n_3968)
);

INVx1_ASAP7_75t_SL g3969 ( 
.A(n_3478),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3636),
.B(n_514),
.Y(n_3970)
);

AOI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3459),
.A2(n_515),
.B(n_516),
.Y(n_3971)
);

HB1xp67_ASAP7_75t_L g3972 ( 
.A(n_3530),
.Y(n_3972)
);

BUFx3_ASAP7_75t_L g3973 ( 
.A(n_3561),
.Y(n_3973)
);

BUFx2_ASAP7_75t_L g3974 ( 
.A(n_3530),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3586),
.Y(n_3975)
);

OAI22xp5_ASAP7_75t_L g3976 ( 
.A1(n_3578),
.A2(n_520),
.B1(n_517),
.B2(n_519),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3596),
.Y(n_3977)
);

CKINVDCx20_ASAP7_75t_R g3978 ( 
.A(n_3722),
.Y(n_3978)
);

OAI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3592),
.A2(n_517),
.B(n_519),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3623),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.Y(n_3980)
);

AOI22xp5_ASAP7_75t_L g3981 ( 
.A1(n_3609),
.A2(n_525),
.B1(n_522),
.B2(n_524),
.Y(n_3981)
);

NAND2xp33_ASAP7_75t_SL g3982 ( 
.A(n_3366),
.B(n_525),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3596),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3673),
.B(n_526),
.Y(n_3984)
);

A2O1A1Ixp33_ASAP7_75t_L g3985 ( 
.A1(n_3437),
.A2(n_528),
.B(n_526),
.C(n_527),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3603),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3603),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3610),
.Y(n_3988)
);

OR2x6_ASAP7_75t_L g3989 ( 
.A(n_3500),
.B(n_527),
.Y(n_3989)
);

NAND3xp33_ASAP7_75t_SL g3990 ( 
.A(n_3607),
.B(n_528),
.C(n_529),
.Y(n_3990)
);

INVx3_ASAP7_75t_L g3991 ( 
.A(n_3537),
.Y(n_3991)
);

OAI22xp5_ASAP7_75t_L g3992 ( 
.A1(n_3579),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_3992)
);

AOI22xp33_ASAP7_75t_L g3993 ( 
.A1(n_3729),
.A2(n_534),
.B1(n_531),
.B2(n_533),
.Y(n_3993)
);

CKINVDCx5p33_ASAP7_75t_R g3994 ( 
.A(n_3637),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_SL g3995 ( 
.A1(n_3637),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_L g3996 ( 
.A1(n_3650),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_3996)
);

OAI22xp5_ASAP7_75t_L g3997 ( 
.A1(n_3559),
.A2(n_3719),
.B1(n_3650),
.B2(n_3681),
.Y(n_3997)
);

AOI221xp5_ASAP7_75t_L g3998 ( 
.A1(n_3466),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.C(n_539),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3657),
.B(n_539),
.Y(n_3999)
);

OA21x2_ASAP7_75t_L g4000 ( 
.A1(n_3554),
.A2(n_540),
.B(n_541),
.Y(n_4000)
);

INVx3_ASAP7_75t_L g4001 ( 
.A(n_3528),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3655),
.A2(n_3706),
.B1(n_3681),
.B2(n_3577),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3610),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3655),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_4004)
);

OAI21x1_ASAP7_75t_L g4005 ( 
.A1(n_3467),
.A2(n_542),
.B(n_543),
.Y(n_4005)
);

AOI21x1_ASAP7_75t_L g4006 ( 
.A1(n_3494),
.A2(n_544),
.B(n_546),
.Y(n_4006)
);

AOI22xp33_ASAP7_75t_L g4007 ( 
.A1(n_3706),
.A2(n_547),
.B1(n_544),
.B2(n_546),
.Y(n_4007)
);

AOI211x1_ASAP7_75t_L g4008 ( 
.A1(n_3703),
.A2(n_549),
.B(n_547),
.C(n_548),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3627),
.B(n_3689),
.Y(n_4009)
);

AND2x4_ASAP7_75t_L g4010 ( 
.A(n_3399),
.B(n_548),
.Y(n_4010)
);

AND2x4_ASAP7_75t_L g4011 ( 
.A(n_3399),
.B(n_550),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3725),
.Y(n_4012)
);

AOI22xp33_ASAP7_75t_L g4013 ( 
.A1(n_3616),
.A2(n_3425),
.B1(n_3615),
.B2(n_3574),
.Y(n_4013)
);

OAI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3715),
.A2(n_838),
.B(n_550),
.Y(n_4014)
);

OAI221xp5_ASAP7_75t_L g4015 ( 
.A1(n_3617),
.A2(n_554),
.B1(n_551),
.B2(n_553),
.C(n_555),
.Y(n_4015)
);

AO21x2_ASAP7_75t_L g4016 ( 
.A1(n_3680),
.A2(n_553),
.B(n_554),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3708),
.B(n_556),
.Y(n_4017)
);

AND2x2_ASAP7_75t_L g4018 ( 
.A(n_3545),
.B(n_3608),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3545),
.B(n_556),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3717),
.Y(n_4020)
);

AOI22xp33_ASAP7_75t_L g4021 ( 
.A1(n_3425),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3725),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3717),
.Y(n_4023)
);

OAI221xp5_ASAP7_75t_L g4024 ( 
.A1(n_3544),
.A2(n_3569),
.B1(n_3704),
.B2(n_3630),
.C(n_3700),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3688),
.Y(n_4025)
);

NOR3xp33_ASAP7_75t_SL g4026 ( 
.A(n_3671),
.B(n_557),
.C(n_558),
.Y(n_4026)
);

OR2x2_ASAP7_75t_L g4027 ( 
.A(n_3608),
.B(n_559),
.Y(n_4027)
);

CKINVDCx5p33_ASAP7_75t_R g4028 ( 
.A(n_3412),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3360),
.B(n_560),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3688),
.Y(n_4030)
);

AOI21xp5_ASAP7_75t_SL g4031 ( 
.A1(n_3412),
.A2(n_560),
.B(n_561),
.Y(n_4031)
);

INVx3_ASAP7_75t_L g4032 ( 
.A(n_3513),
.Y(n_4032)
);

CKINVDCx6p67_ASAP7_75t_R g4033 ( 
.A(n_3538),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3439),
.Y(n_4034)
);

INVxp67_ASAP7_75t_SL g4035 ( 
.A(n_3696),
.Y(n_4035)
);

INVx6_ASAP7_75t_L g4036 ( 
.A(n_3513),
.Y(n_4036)
);

CKINVDCx20_ASAP7_75t_R g4037 ( 
.A(n_3495),
.Y(n_4037)
);

INVxp67_ASAP7_75t_L g4038 ( 
.A(n_3663),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3439),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_L g4040 ( 
.A(n_3360),
.B(n_561),
.Y(n_4040)
);

INVx3_ASAP7_75t_L g4041 ( 
.A(n_3515),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3382),
.B(n_562),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_3452),
.Y(n_4043)
);

INVx5_ASAP7_75t_L g4044 ( 
.A(n_3601),
.Y(n_4044)
);

AOI21x1_ASAP7_75t_L g4045 ( 
.A1(n_3699),
.A2(n_562),
.B(n_563),
.Y(n_4045)
);

CKINVDCx6p67_ASAP7_75t_R g4046 ( 
.A(n_3515),
.Y(n_4046)
);

AND2x4_ASAP7_75t_L g4047 ( 
.A(n_3652),
.B(n_563),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3574),
.A2(n_567),
.B1(n_564),
.B2(n_566),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_L g4049 ( 
.A1(n_3615),
.A2(n_568),
.B1(n_564),
.B2(n_567),
.Y(n_4049)
);

AND2x4_ASAP7_75t_L g4050 ( 
.A(n_3652),
.B(n_569),
.Y(n_4050)
);

OAI22xp5_ASAP7_75t_L g4051 ( 
.A1(n_3690),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_4051)
);

CKINVDCx11_ASAP7_75t_R g4052 ( 
.A(n_3601),
.Y(n_4052)
);

CKINVDCx5p33_ASAP7_75t_R g4053 ( 
.A(n_3601),
.Y(n_4053)
);

AOI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3740),
.A2(n_3638),
.B1(n_3709),
.B2(n_3663),
.Y(n_4054)
);

OAI22xp5_ASAP7_75t_L g4055 ( 
.A1(n_3780),
.A2(n_3690),
.B1(n_3712),
.B2(n_3656),
.Y(n_4055)
);

OR2x2_ASAP7_75t_L g4056 ( 
.A(n_3730),
.B(n_3377),
.Y(n_4056)
);

OAI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3774),
.A2(n_3712),
.B1(n_3656),
.B2(n_3624),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3736),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3754),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_L g4060 ( 
.A1(n_3753),
.A2(n_3709),
.B1(n_3692),
.B2(n_3675),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3739),
.Y(n_4061)
);

INVx2_ASAP7_75t_SL g4062 ( 
.A(n_3881),
.Y(n_4062)
);

AOI221xp5_ASAP7_75t_L g4063 ( 
.A1(n_3747),
.A2(n_3701),
.B1(n_3716),
.B2(n_3699),
.C(n_3676),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_3851),
.B(n_3382),
.Y(n_4064)
);

NAND3xp33_ASAP7_75t_L g4065 ( 
.A(n_3777),
.B(n_3716),
.C(n_3666),
.Y(n_4065)
);

OAI221xp5_ASAP7_75t_L g4066 ( 
.A1(n_3888),
.A2(n_3666),
.B1(n_3676),
.B2(n_3664),
.C(n_3389),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3792),
.A2(n_3720),
.B1(n_3632),
.B2(n_3643),
.Y(n_4067)
);

OAI21xp5_ASAP7_75t_L g4068 ( 
.A1(n_3985),
.A2(n_3665),
.B(n_3626),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3756),
.Y(n_4069)
);

INVx3_ASAP7_75t_L g4070 ( 
.A(n_3782),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3805),
.A2(n_3720),
.B1(n_3638),
.B2(n_3600),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_3759),
.A2(n_3506),
.B1(n_3493),
.B2(n_3631),
.Y(n_4072)
);

BUFx2_ASAP7_75t_L g4073 ( 
.A(n_3808),
.Y(n_4073)
);

OAI221xp5_ASAP7_75t_L g4074 ( 
.A1(n_3778),
.A2(n_3664),
.B1(n_3653),
.B2(n_3639),
.C(n_3631),
.Y(n_4074)
);

AOI222xp33_ASAP7_75t_L g4075 ( 
.A1(n_3786),
.A2(n_3787),
.B1(n_3781),
.B2(n_3758),
.C1(n_3919),
.C2(n_3825),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3757),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3803),
.A2(n_3506),
.B1(n_3493),
.B2(n_3639),
.Y(n_4077)
);

OAI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3916),
.A2(n_3516),
.B1(n_3624),
.B2(n_3410),
.Y(n_4078)
);

OAI221xp5_ASAP7_75t_L g4079 ( 
.A1(n_3773),
.A2(n_3653),
.B1(n_3614),
.B2(n_3620),
.C(n_3612),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3784),
.A2(n_3516),
.B1(n_3372),
.B2(n_3397),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3765),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_3748),
.Y(n_4082)
);

AOI22xp33_ASAP7_75t_L g4083 ( 
.A1(n_3998),
.A2(n_3614),
.B1(n_3620),
.B2(n_3612),
.Y(n_4083)
);

OAI22xp33_ASAP7_75t_L g4084 ( 
.A1(n_3908),
.A2(n_3410),
.B1(n_3421),
.B2(n_3406),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3751),
.Y(n_4085)
);

AO21x2_ASAP7_75t_L g4086 ( 
.A1(n_3873),
.A2(n_3452),
.B(n_3421),
.Y(n_4086)
);

NAND3xp33_ASAP7_75t_L g4087 ( 
.A(n_3875),
.B(n_3397),
.C(n_3379),
.Y(n_4087)
);

INVx5_ASAP7_75t_SL g4088 ( 
.A(n_3770),
.Y(n_4088)
);

AOI22xp33_ASAP7_75t_L g4089 ( 
.A1(n_3990),
.A2(n_3406),
.B1(n_3379),
.B2(n_3679),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3796),
.A2(n_3687),
.B1(n_3707),
.B2(n_3713),
.Y(n_4090)
);

OR2x2_ASAP7_75t_L g4091 ( 
.A(n_3819),
.B(n_3377),
.Y(n_4091)
);

AOI222xp33_ASAP7_75t_L g4092 ( 
.A1(n_3786),
.A2(n_3711),
.B1(n_3568),
.B2(n_3654),
.C1(n_3634),
.C2(n_3580),
.Y(n_4092)
);

OAI22xp5_ASAP7_75t_L g4093 ( 
.A1(n_4002),
.A2(n_3752),
.B1(n_3908),
.B2(n_3989),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3772),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3833),
.B(n_3377),
.Y(n_4095)
);

HB1xp67_ASAP7_75t_L g4096 ( 
.A(n_3808),
.Y(n_4096)
);

INVx5_ASAP7_75t_SL g4097 ( 
.A(n_3963),
.Y(n_4097)
);

AOI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3749),
.A2(n_3350),
.B1(n_3512),
.B2(n_3543),
.Y(n_4098)
);

AOI211xp5_ASAP7_75t_L g4099 ( 
.A1(n_4031),
.A2(n_3648),
.B(n_3588),
.C(n_3590),
.Y(n_4099)
);

OA21x2_ASAP7_75t_L g4100 ( 
.A1(n_3738),
.A2(n_3670),
.B(n_3436),
.Y(n_4100)
);

OR2x6_ASAP7_75t_L g4101 ( 
.A(n_3963),
.B(n_3954),
.Y(n_4101)
);

OAI22xp5_ASAP7_75t_L g4102 ( 
.A1(n_3989),
.A2(n_3337),
.B1(n_3460),
.B2(n_3628),
.Y(n_4102)
);

OAI22xp5_ASAP7_75t_L g4103 ( 
.A1(n_3995),
.A2(n_3337),
.B1(n_3628),
.B2(n_3382),
.Y(n_4103)
);

AOI22xp33_ASAP7_75t_L g4104 ( 
.A1(n_3800),
.A2(n_3355),
.B1(n_3647),
.B2(n_3546),
.Y(n_4104)
);

OAI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_3952),
.A2(n_3598),
.B(n_3575),
.Y(n_4105)
);

OAI221xp5_ASAP7_75t_L g4106 ( 
.A1(n_3746),
.A2(n_3628),
.B1(n_3589),
.B2(n_3587),
.C(n_3640),
.Y(n_4106)
);

INVx1_ASAP7_75t_SL g4107 ( 
.A(n_3894),
.Y(n_4107)
);

OAI221xp5_ASAP7_75t_L g4108 ( 
.A1(n_3850),
.A2(n_3589),
.B1(n_3587),
.B2(n_3640),
.C(n_3451),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_L g4109 ( 
.A1(n_3931),
.A2(n_3602),
.B1(n_3605),
.B2(n_3604),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_3891),
.B(n_3451),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_3886),
.B(n_3451),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3783),
.Y(n_4112)
);

A2O1A1Ixp33_ASAP7_75t_SL g4113 ( 
.A1(n_3857),
.A2(n_3587),
.B(n_3589),
.C(n_3640),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3858),
.A2(n_3621),
.B1(n_3567),
.B2(n_3658),
.Y(n_4114)
);

OA21x2_ASAP7_75t_L g4115 ( 
.A1(n_4038),
.A2(n_3434),
.B(n_3474),
.Y(n_4115)
);

CKINVDCx20_ASAP7_75t_R g4116 ( 
.A(n_3733),
.Y(n_4116)
);

AO21x2_ASAP7_75t_L g4117 ( 
.A1(n_3854),
.A2(n_3476),
.B(n_3481),
.Y(n_4117)
);

OAI221xp5_ASAP7_75t_L g4118 ( 
.A1(n_3855),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.C(n_574),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3797),
.Y(n_4119)
);

OAI22xp5_ASAP7_75t_L g4120 ( 
.A1(n_3994),
.A2(n_3499),
.B1(n_3510),
.B2(n_3491),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_L g4121 ( 
.A1(n_3950),
.A2(n_3642),
.B1(n_3408),
.B2(n_3371),
.Y(n_4121)
);

OAI21x1_ASAP7_75t_SL g4122 ( 
.A1(n_3954),
.A2(n_573),
.B(n_576),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3936),
.A2(n_3629),
.B1(n_3391),
.B2(n_3490),
.Y(n_4123)
);

OAI211xp5_ASAP7_75t_L g4124 ( 
.A1(n_3823),
.A2(n_3488),
.B(n_3407),
.C(n_3405),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_3920),
.B(n_3398),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3804),
.Y(n_4126)
);

OAI221xp5_ASAP7_75t_L g4127 ( 
.A1(n_3903),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.C(n_580),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3939),
.A2(n_3429),
.B1(n_3536),
.B2(n_3535),
.Y(n_4128)
);

OAI322xp33_ASAP7_75t_L g4129 ( 
.A1(n_3741),
.A2(n_3922),
.A3(n_3845),
.B1(n_3812),
.B2(n_3928),
.C1(n_4009),
.C2(n_3866),
.Y(n_4129)
);

AND2x4_ASAP7_75t_L g4130 ( 
.A(n_3782),
.B(n_3339),
.Y(n_4130)
);

AOI21xp5_ASAP7_75t_L g4131 ( 
.A1(n_3840),
.A2(n_3524),
.B(n_3521),
.Y(n_4131)
);

AO21x1_ASAP7_75t_L g4132 ( 
.A1(n_3938),
.A2(n_3527),
.B(n_3354),
.Y(n_4132)
);

BUFx4f_ASAP7_75t_SL g4133 ( 
.A(n_3842),
.Y(n_4133)
);

OAI22xp5_ASAP7_75t_L g4134 ( 
.A1(n_4046),
.A2(n_3419),
.B1(n_3359),
.B2(n_3562),
.Y(n_4134)
);

AO21x2_ASAP7_75t_L g4135 ( 
.A1(n_3882),
.A2(n_3486),
.B(n_3448),
.Y(n_4135)
);

A2O1A1Ixp33_ASAP7_75t_L g4136 ( 
.A1(n_3982),
.A2(n_3446),
.B(n_3456),
.C(n_3443),
.Y(n_4136)
);

OAI21xp5_ASAP7_75t_SL g4137 ( 
.A1(n_3737),
.A2(n_578),
.B(n_579),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_3779),
.B(n_582),
.Y(n_4138)
);

OAI22xp5_ASAP7_75t_L g4139 ( 
.A1(n_3980),
.A2(n_3461),
.B1(n_3385),
.B2(n_3349),
.Y(n_4139)
);

OAI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_3940),
.A2(n_582),
.B(n_583),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_L g4141 ( 
.A1(n_3828),
.A2(n_586),
.B1(n_584),
.B2(n_585),
.Y(n_4141)
);

AOI22xp33_ASAP7_75t_L g4142 ( 
.A1(n_3847),
.A2(n_588),
.B1(n_584),
.B2(n_587),
.Y(n_4142)
);

BUFx3_ASAP7_75t_L g4143 ( 
.A(n_3742),
.Y(n_4143)
);

OAI22xp33_ASAP7_75t_L g4144 ( 
.A1(n_3735),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3818),
.Y(n_4145)
);

OAI22xp5_ASAP7_75t_L g4146 ( 
.A1(n_3996),
.A2(n_591),
.B1(n_589),
.B2(n_590),
.Y(n_4146)
);

AOI221xp5_ASAP7_75t_L g4147 ( 
.A1(n_3926),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.C(n_594),
.Y(n_4147)
);

OAI21x1_ASAP7_75t_L g4148 ( 
.A1(n_3809),
.A2(n_592),
.B(n_595),
.Y(n_4148)
);

HB1xp67_ASAP7_75t_L g4149 ( 
.A(n_3808),
.Y(n_4149)
);

AOI222xp33_ASAP7_75t_L g4150 ( 
.A1(n_3885),
.A2(n_596),
.B1(n_597),
.B2(n_598),
.C1(n_599),
.C2(n_601),
.Y(n_4150)
);

AOI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_3997),
.A2(n_601),
.B1(n_596),
.B2(n_598),
.Y(n_4151)
);

NAND3xp33_ASAP7_75t_L g4152 ( 
.A(n_3917),
.B(n_603),
.C(n_604),
.Y(n_4152)
);

AND2x4_ASAP7_75t_L g4153 ( 
.A(n_3785),
.B(n_604),
.Y(n_4153)
);

INVx3_ASAP7_75t_L g4154 ( 
.A(n_3785),
.Y(n_4154)
);

OAI22xp5_ASAP7_75t_L g4155 ( 
.A1(n_4004),
.A2(n_609),
.B1(n_605),
.B2(n_608),
.Y(n_4155)
);

AOI22xp33_ASAP7_75t_L g4156 ( 
.A1(n_3816),
.A2(n_609),
.B1(n_605),
.B2(n_608),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_3849),
.B(n_610),
.Y(n_4157)
);

OAI21xp5_ASAP7_75t_L g4158 ( 
.A1(n_4051),
.A2(n_610),
.B(n_611),
.Y(n_4158)
);

OR2x2_ASAP7_75t_L g4159 ( 
.A(n_3844),
.B(n_612),
.Y(n_4159)
);

INVx2_ASAP7_75t_SL g4160 ( 
.A(n_3811),
.Y(n_4160)
);

OAI22xp5_ASAP7_75t_L g4161 ( 
.A1(n_4007),
.A2(n_615),
.B1(n_613),
.B2(n_614),
.Y(n_4161)
);

OAI22xp33_ASAP7_75t_L g4162 ( 
.A1(n_3755),
.A2(n_838),
.B1(n_616),
.B2(n_613),
.Y(n_4162)
);

AOI222xp33_ASAP7_75t_L g4163 ( 
.A1(n_3960),
.A2(n_615),
.B1(n_620),
.B2(n_621),
.C1(n_622),
.C2(n_623),
.Y(n_4163)
);

AOI22xp33_ASAP7_75t_L g4164 ( 
.A1(n_3906),
.A2(n_624),
.B1(n_620),
.B2(n_621),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3871),
.B(n_625),
.Y(n_4165)
);

AO21x2_ASAP7_75t_L g4166 ( 
.A1(n_4029),
.A2(n_625),
.B(n_626),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3820),
.Y(n_4167)
);

AOI22xp33_ASAP7_75t_L g4168 ( 
.A1(n_3793),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_4168)
);

OAI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3755),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_3861),
.B(n_837),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_SL g4171 ( 
.A1(n_3829),
.A2(n_632),
.B1(n_629),
.B2(n_630),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3826),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3878),
.B(n_632),
.Y(n_4173)
);

AND2x2_ASAP7_75t_L g4174 ( 
.A(n_3913),
.B(n_634),
.Y(n_4174)
);

OAI322xp33_ASAP7_75t_L g4175 ( 
.A1(n_3869),
.A2(n_635),
.A3(n_636),
.B1(n_637),
.B2(n_638),
.C1(n_639),
.C2(n_640),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_3761),
.Y(n_4176)
);

OR2x2_ASAP7_75t_L g4177 ( 
.A(n_3923),
.B(n_635),
.Y(n_4177)
);

OAI22xp5_ASAP7_75t_L g4178 ( 
.A1(n_3788),
.A2(n_638),
.B1(n_636),
.B2(n_637),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_3766),
.Y(n_4179)
);

OAI22xp5_ASAP7_75t_L g4180 ( 
.A1(n_3993),
.A2(n_644),
.B1(n_642),
.B2(n_643),
.Y(n_4180)
);

OAI221xp5_ASAP7_75t_L g4181 ( 
.A1(n_3837),
.A2(n_3852),
.B1(n_3843),
.B2(n_3864),
.C(n_3901),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3830),
.Y(n_4182)
);

OAI22xp5_ASAP7_75t_L g4183 ( 
.A1(n_4026),
.A2(n_646),
.B1(n_643),
.B2(n_644),
.Y(n_4183)
);

OAI22xp33_ASAP7_75t_L g4184 ( 
.A1(n_3771),
.A2(n_837),
.B1(n_649),
.B2(n_647),
.Y(n_4184)
);

OAI211xp5_ASAP7_75t_L g4185 ( 
.A1(n_3941),
.A2(n_650),
.B(n_647),
.C(n_648),
.Y(n_4185)
);

AOI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_3831),
.A2(n_3912),
.B1(n_3976),
.B2(n_3810),
.Y(n_4186)
);

CKINVDCx5p33_ASAP7_75t_R g4187 ( 
.A(n_3863),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3884),
.B(n_648),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_3822),
.B(n_836),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_3832),
.B(n_836),
.Y(n_4190)
);

OAI22xp33_ASAP7_75t_L g4191 ( 
.A1(n_3771),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_4191)
);

CKINVDCx5p33_ASAP7_75t_R g4192 ( 
.A(n_3791),
.Y(n_4192)
);

AOI22xp33_ASAP7_75t_SL g4193 ( 
.A1(n_3829),
.A2(n_653),
.B1(n_651),
.B2(n_652),
.Y(n_4193)
);

OAI221xp5_ASAP7_75t_L g4194 ( 
.A1(n_3961),
.A2(n_654),
.B1(n_655),
.B2(n_657),
.C(n_658),
.Y(n_4194)
);

AOI33xp33_ASAP7_75t_L g4195 ( 
.A1(n_3944),
.A2(n_3947),
.A3(n_4049),
.B1(n_4048),
.B2(n_3925),
.B3(n_3984),
.Y(n_4195)
);

OAI21xp33_ASAP7_75t_L g4196 ( 
.A1(n_4013),
.A2(n_655),
.B(n_657),
.Y(n_4196)
);

NOR2xp33_ASAP7_75t_SL g4197 ( 
.A(n_3839),
.B(n_658),
.Y(n_4197)
);

AOI22xp33_ASAP7_75t_L g4198 ( 
.A1(n_3876),
.A2(n_662),
.B1(n_659),
.B2(n_660),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_3835),
.B(n_659),
.Y(n_4199)
);

AOI221xp5_ASAP7_75t_L g4200 ( 
.A1(n_4008),
.A2(n_662),
.B1(n_663),
.B2(n_664),
.C(n_665),
.Y(n_4200)
);

AOI22xp33_ASAP7_75t_L g4201 ( 
.A1(n_3877),
.A2(n_668),
.B1(n_666),
.B2(n_667),
.Y(n_4201)
);

INVx3_ASAP7_75t_L g4202 ( 
.A(n_3957),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3801),
.A2(n_666),
.B(n_667),
.Y(n_4203)
);

A2O1A1Ixp33_ASAP7_75t_L g4204 ( 
.A1(n_3937),
.A2(n_671),
.B(n_669),
.C(n_670),
.Y(n_4204)
);

INVxp67_ASAP7_75t_SL g4205 ( 
.A(n_3972),
.Y(n_4205)
);

AO21x2_ASAP7_75t_L g4206 ( 
.A1(n_4040),
.A2(n_669),
.B(n_671),
.Y(n_4206)
);

OAI211xp5_ASAP7_75t_L g4207 ( 
.A1(n_3981),
.A2(n_675),
.B(n_673),
.C(n_674),
.Y(n_4207)
);

AOI22xp33_ASAP7_75t_L g4208 ( 
.A1(n_3817),
.A2(n_677),
.B1(n_673),
.B2(n_676),
.Y(n_4208)
);

HB1xp67_ASAP7_75t_L g4209 ( 
.A(n_3974),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3775),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_3790),
.Y(n_4211)
);

OR2x2_ASAP7_75t_L g4212 ( 
.A(n_3807),
.B(n_676),
.Y(n_4212)
);

NOR2xp33_ASAP7_75t_L g4213 ( 
.A(n_3734),
.B(n_835),
.Y(n_4213)
);

HB1xp67_ASAP7_75t_L g4214 ( 
.A(n_3964),
.Y(n_4214)
);

AOI22xp33_ASAP7_75t_L g4215 ( 
.A1(n_4015),
.A2(n_680),
.B1(n_678),
.B2(n_679),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_3836),
.B(n_678),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_3956),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_4217)
);

OAI221xp5_ASAP7_75t_L g4218 ( 
.A1(n_3933),
.A2(n_681),
.B1(n_683),
.B2(n_684),
.C(n_686),
.Y(n_4218)
);

AOI211xp5_ASAP7_75t_L g4219 ( 
.A1(n_3776),
.A2(n_686),
.B(n_683),
.C(n_684),
.Y(n_4219)
);

AND2x4_ASAP7_75t_L g4220 ( 
.A(n_3841),
.B(n_687),
.Y(n_4220)
);

AOI221xp5_ASAP7_75t_L g4221 ( 
.A1(n_3970),
.A2(n_688),
.B1(n_689),
.B2(n_690),
.C(n_691),
.Y(n_4221)
);

OAI211xp5_ASAP7_75t_L g4222 ( 
.A1(n_3887),
.A2(n_690),
.B(n_688),
.C(n_689),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_3838),
.B(n_692),
.Y(n_4223)
);

OAI21xp33_ASAP7_75t_L g4224 ( 
.A1(n_3874),
.A2(n_692),
.B(n_695),
.Y(n_4224)
);

AOI21xp33_ASAP7_75t_L g4225 ( 
.A1(n_3924),
.A2(n_695),
.B(n_696),
.Y(n_4225)
);

OAI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_3893),
.A2(n_3897),
.B1(n_3918),
.B2(n_3914),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_SL g4227 ( 
.A(n_3798),
.B(n_697),
.Y(n_4227)
);

OAI21xp5_ASAP7_75t_SL g4228 ( 
.A1(n_3946),
.A2(n_698),
.B(n_699),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3846),
.Y(n_4229)
);

INVx2_ASAP7_75t_SL g4230 ( 
.A(n_3900),
.Y(n_4230)
);

AOI22xp33_ASAP7_75t_L g4231 ( 
.A1(n_3949),
.A2(n_702),
.B1(n_700),
.B2(n_701),
.Y(n_4231)
);

OAI211xp5_ASAP7_75t_L g4232 ( 
.A1(n_3896),
.A2(n_705),
.B(n_703),
.C(n_704),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3853),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_3856),
.B(n_834),
.Y(n_4234)
);

INVx4_ASAP7_75t_L g4235 ( 
.A(n_3743),
.Y(n_4235)
);

AOI22xp33_ASAP7_75t_L g4236 ( 
.A1(n_3979),
.A2(n_705),
.B1(n_703),
.B2(n_704),
.Y(n_4236)
);

NOR2xp33_ASAP7_75t_L g4237 ( 
.A(n_3824),
.B(n_706),
.Y(n_4237)
);

INVx1_ASAP7_75t_SL g4238 ( 
.A(n_3978),
.Y(n_4238)
);

AOI22xp33_ASAP7_75t_L g4239 ( 
.A1(n_3968),
.A2(n_709),
.B1(n_707),
.B2(n_708),
.Y(n_4239)
);

AOI221xp5_ASAP7_75t_L g4240 ( 
.A1(n_3999),
.A2(n_710),
.B1(n_712),
.B2(n_713),
.C(n_714),
.Y(n_4240)
);

OR2x2_ASAP7_75t_L g4241 ( 
.A(n_3930),
.B(n_3744),
.Y(n_4241)
);

O2A1O1Ixp33_ASAP7_75t_SL g4242 ( 
.A1(n_3848),
.A2(n_716),
.B(n_710),
.C(n_712),
.Y(n_4242)
);

INVx3_ASAP7_75t_L g4243 ( 
.A(n_3745),
.Y(n_4243)
);

OR2x2_ASAP7_75t_L g4244 ( 
.A(n_3750),
.B(n_717),
.Y(n_4244)
);

INVx2_ASAP7_75t_L g4245 ( 
.A(n_3942),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3975),
.Y(n_4246)
);

AOI22xp33_ASAP7_75t_L g4247 ( 
.A1(n_4042),
.A2(n_719),
.B1(n_717),
.B2(n_718),
.Y(n_4247)
);

AO21x2_ASAP7_75t_L g4248 ( 
.A1(n_3907),
.A2(n_718),
.B(n_720),
.Y(n_4248)
);

AOI22xp33_ASAP7_75t_L g4249 ( 
.A1(n_4014),
.A2(n_722),
.B1(n_720),
.B2(n_721),
.Y(n_4249)
);

OAI221xp5_ASAP7_75t_L g4250 ( 
.A1(n_3867),
.A2(n_721),
.B1(n_722),
.B2(n_723),
.C(n_724),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_4003),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_3927),
.Y(n_4252)
);

AOI221xp5_ASAP7_75t_L g4253 ( 
.A1(n_4017),
.A2(n_723),
.B1(n_725),
.B2(n_726),
.C(n_727),
.Y(n_4253)
);

AND2x2_ASAP7_75t_L g4254 ( 
.A(n_3879),
.B(n_728),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3932),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3870),
.B(n_4018),
.Y(n_4256)
);

AOI221xp5_ASAP7_75t_L g4257 ( 
.A1(n_3883),
.A2(n_728),
.B1(n_731),
.B2(n_732),
.C(n_733),
.Y(n_4257)
);

AOI22xp33_ASAP7_75t_L g4258 ( 
.A1(n_4024),
.A2(n_733),
.B1(n_734),
.B2(n_735),
.Y(n_4258)
);

AND2x4_ASAP7_75t_L g4259 ( 
.A(n_3909),
.B(n_734),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_3893),
.A2(n_735),
.B1(n_736),
.B2(n_737),
.Y(n_4260)
);

AOI221xp5_ASAP7_75t_L g4261 ( 
.A1(n_3895),
.A2(n_737),
.B1(n_738),
.B2(n_739),
.C(n_740),
.Y(n_4261)
);

AOI221xp5_ASAP7_75t_L g4262 ( 
.A1(n_3872),
.A2(n_738),
.B1(n_739),
.B2(n_740),
.C(n_741),
.Y(n_4262)
);

NOR2x1_ASAP7_75t_L g4263 ( 
.A(n_3897),
.B(n_741),
.Y(n_4263)
);

OAI221xp5_ASAP7_75t_L g4264 ( 
.A1(n_3813),
.A2(n_742),
.B1(n_743),
.B2(n_746),
.C(n_747),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_3959),
.B(n_834),
.Y(n_4265)
);

AOI22xp5_ASAP7_75t_L g4266 ( 
.A1(n_3914),
.A2(n_3918),
.B1(n_3948),
.B2(n_4010),
.Y(n_4266)
);

OAI22xp33_ASAP7_75t_L g4267 ( 
.A1(n_4033),
.A2(n_742),
.B1(n_743),
.B2(n_746),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_4209),
.B(n_3762),
.Y(n_4268)
);

INVx2_ASAP7_75t_L g4269 ( 
.A(n_4245),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4058),
.Y(n_4270)
);

INVx1_ASAP7_75t_L g4271 ( 
.A(n_4059),
.Y(n_4271)
);

INVxp67_ASAP7_75t_SL g4272 ( 
.A(n_4205),
.Y(n_4272)
);

AOI22xp5_ASAP7_75t_L g4273 ( 
.A1(n_4093),
.A2(n_3948),
.B1(n_4011),
.B2(n_4010),
.Y(n_4273)
);

INVxp67_ASAP7_75t_SL g4274 ( 
.A(n_4056),
.Y(n_4274)
);

AOI22xp33_ASAP7_75t_L g4275 ( 
.A1(n_4181),
.A2(n_3767),
.B1(n_3827),
.B2(n_3802),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4256),
.B(n_3934),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4246),
.Y(n_4277)
);

BUFx2_ASAP7_75t_L g4278 ( 
.A(n_4101),
.Y(n_4278)
);

HB1xp67_ASAP7_75t_L g4279 ( 
.A(n_4096),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4069),
.Y(n_4280)
);

INVx3_ASAP7_75t_L g4281 ( 
.A(n_4070),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4064),
.B(n_3966),
.Y(n_4282)
);

AND2x4_ASAP7_75t_L g4283 ( 
.A(n_4202),
.B(n_3731),
.Y(n_4283)
);

HB1xp67_ASAP7_75t_L g4284 ( 
.A(n_4149),
.Y(n_4284)
);

INVx3_ASAP7_75t_L g4285 ( 
.A(n_4070),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4202),
.B(n_4214),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4076),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_4190),
.B(n_3768),
.Y(n_4288)
);

AND2x2_ASAP7_75t_L g4289 ( 
.A(n_4241),
.B(n_3977),
.Y(n_4289)
);

OA21x2_ASAP7_75t_L g4290 ( 
.A1(n_4136),
.A2(n_3821),
.B(n_3806),
.Y(n_4290)
);

OR2x2_ASAP7_75t_L g4291 ( 
.A(n_4091),
.B(n_3795),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4251),
.Y(n_4292)
);

AND2x4_ASAP7_75t_L g4293 ( 
.A(n_4243),
.B(n_3731),
.Y(n_4293)
);

BUFx2_ASAP7_75t_L g4294 ( 
.A(n_4101),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4081),
.Y(n_4295)
);

AND2x2_ASAP7_75t_L g4296 ( 
.A(n_4073),
.B(n_3983),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4094),
.Y(n_4297)
);

HB1xp67_ASAP7_75t_L g4298 ( 
.A(n_4061),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_4082),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4112),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4085),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4176),
.Y(n_4302)
);

AO21x2_ASAP7_75t_L g4303 ( 
.A1(n_4084),
.A2(n_4045),
.B(n_3965),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4119),
.Y(n_4304)
);

HB1xp67_ASAP7_75t_L g4305 ( 
.A(n_4179),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4211),
.Y(n_4306)
);

AO31x2_ASAP7_75t_L g4307 ( 
.A1(n_4132),
.A2(n_4057),
.A3(n_4080),
.B(n_4055),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4126),
.B(n_3872),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4145),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4252),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4255),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4167),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4172),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4210),
.Y(n_4314)
);

HB1xp67_ASAP7_75t_L g4315 ( 
.A(n_4229),
.Y(n_4315)
);

OR2x2_ASAP7_75t_L g4316 ( 
.A(n_4233),
.B(n_3732),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4182),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4110),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4125),
.B(n_4012),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4111),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4174),
.B(n_3986),
.Y(n_4321)
);

AND2x2_ASAP7_75t_L g4322 ( 
.A(n_4243),
.B(n_3987),
.Y(n_4322)
);

NOR2xp33_ASAP7_75t_L g4323 ( 
.A(n_4129),
.B(n_4159),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_4075),
.B(n_4022),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_4254),
.B(n_4154),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4154),
.Y(n_4326)
);

INVx2_ASAP7_75t_SL g4327 ( 
.A(n_4062),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4115),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_4095),
.B(n_3732),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4115),
.Y(n_4330)
);

OR2x2_ASAP7_75t_L g4331 ( 
.A(n_4107),
.B(n_4226),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4170),
.B(n_3988),
.Y(n_4332)
);

BUFx3_ASAP7_75t_L g4333 ( 
.A(n_4230),
.Y(n_4333)
);

NOR2x1_ASAP7_75t_L g4334 ( 
.A(n_4143),
.B(n_4037),
.Y(n_4334)
);

INVx3_ASAP7_75t_SL g4335 ( 
.A(n_4116),
.Y(n_4335)
);

OR2x2_ASAP7_75t_L g4336 ( 
.A(n_4177),
.B(n_3859),
.Y(n_4336)
);

OR2x2_ASAP7_75t_L g4337 ( 
.A(n_4087),
.B(n_3859),
.Y(n_4337)
);

INVx5_ASAP7_75t_L g4338 ( 
.A(n_4097),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4189),
.B(n_4023),
.Y(n_4339)
);

OR2x2_ASAP7_75t_L g4340 ( 
.A(n_4138),
.B(n_3892),
.Y(n_4340)
);

OAI221xp5_ASAP7_75t_L g4341 ( 
.A1(n_4228),
.A2(n_3951),
.B1(n_3953),
.B2(n_3962),
.C(n_3958),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4199),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4130),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_4130),
.Y(n_4344)
);

NOR2xp67_ASAP7_75t_L g4345 ( 
.A(n_4235),
.B(n_3862),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4266),
.B(n_3915),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4157),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4220),
.B(n_4020),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_4220),
.B(n_3892),
.Y(n_4349)
);

HB1xp67_ASAP7_75t_L g4350 ( 
.A(n_4086),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4165),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4212),
.Y(n_4352)
);

BUFx2_ASAP7_75t_L g4353 ( 
.A(n_4235),
.Y(n_4353)
);

AND2x2_ASAP7_75t_L g4354 ( 
.A(n_4160),
.B(n_3909),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4216),
.Y(n_4355)
);

HB1xp67_ASAP7_75t_L g4356 ( 
.A(n_4086),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_4153),
.B(n_3991),
.Y(n_4357)
);

INVx3_ASAP7_75t_L g4358 ( 
.A(n_4153),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4100),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4100),
.Y(n_4360)
);

INVx2_ASAP7_75t_L g4361 ( 
.A(n_4135),
.Y(n_4361)
);

NAND2x1p5_ASAP7_75t_L g4362 ( 
.A(n_4259),
.B(n_4044),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4135),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4223),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4234),
.Y(n_4365)
);

NOR2x1p5_ASAP7_75t_L g4366 ( 
.A(n_4187),
.B(n_4028),
.Y(n_4366)
);

OAI211xp5_ASAP7_75t_L g4367 ( 
.A1(n_4137),
.A2(n_3899),
.B(n_4052),
.C(n_4001),
.Y(n_4367)
);

OR2x2_ASAP7_75t_L g4368 ( 
.A(n_4244),
.B(n_4034),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4315),
.Y(n_4369)
);

OAI221xp5_ASAP7_75t_L g4370 ( 
.A1(n_4273),
.A2(n_4197),
.B1(n_4127),
.B2(n_4186),
.C(n_4140),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4298),
.Y(n_4371)
);

AOI221xp5_ASAP7_75t_L g4372 ( 
.A1(n_4323),
.A2(n_4218),
.B1(n_4213),
.B2(n_4118),
.C(n_4175),
.Y(n_4372)
);

AOI221xp5_ASAP7_75t_L g4373 ( 
.A1(n_4323),
.A2(n_4103),
.B1(n_4267),
.B2(n_4162),
.C(n_4184),
.Y(n_4373)
);

AOI222xp33_ASAP7_75t_L g4374 ( 
.A1(n_4324),
.A2(n_4262),
.B1(n_4261),
.B2(n_4152),
.C1(n_4237),
.C2(n_4133),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_4276),
.B(n_4054),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_L g4376 ( 
.A1(n_4367),
.A2(n_4227),
.B(n_4224),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4275),
.A2(n_4063),
.B1(n_4196),
.B2(n_4217),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4315),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4270),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_L g4380 ( 
.A(n_4335),
.B(n_4238),
.Y(n_4380)
);

OR2x2_ASAP7_75t_L g4381 ( 
.A(n_4291),
.B(n_4039),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4298),
.Y(n_4382)
);

OR2x2_ASAP7_75t_L g4383 ( 
.A(n_4272),
.B(n_4043),
.Y(n_4383)
);

OAI211xp5_ASAP7_75t_SL g4384 ( 
.A1(n_4275),
.A2(n_4163),
.B(n_4219),
.C(n_4195),
.Y(n_4384)
);

HB1xp67_ASAP7_75t_L g4385 ( 
.A(n_4305),
.Y(n_4385)
);

OR2x2_ASAP7_75t_L g4386 ( 
.A(n_4272),
.B(n_4025),
.Y(n_4386)
);

OAI33xp33_ASAP7_75t_L g4387 ( 
.A1(n_4331),
.A2(n_4191),
.A3(n_4169),
.B1(n_4183),
.B2(n_4260),
.B3(n_4078),
.Y(n_4387)
);

OR2x2_ASAP7_75t_L g4388 ( 
.A(n_4268),
.B(n_4030),
.Y(n_4388)
);

AOI22xp33_ASAP7_75t_L g4389 ( 
.A1(n_4346),
.A2(n_4151),
.B1(n_4257),
.B2(n_4194),
.Y(n_4389)
);

BUFx2_ASAP7_75t_L g4390 ( 
.A(n_4333),
.Y(n_4390)
);

BUFx6f_ASAP7_75t_L g4391 ( 
.A(n_4338),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4271),
.Y(n_4392)
);

NOR2xp33_ASAP7_75t_R g4393 ( 
.A(n_4335),
.B(n_3868),
.Y(n_4393)
);

NOR2xp33_ASAP7_75t_L g4394 ( 
.A(n_4333),
.B(n_4192),
.Y(n_4394)
);

INVxp67_ASAP7_75t_L g4395 ( 
.A(n_4279),
.Y(n_4395)
);

OAI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_4367),
.A2(n_4263),
.B(n_4204),
.Y(n_4396)
);

OR2x2_ASAP7_75t_L g4397 ( 
.A(n_4274),
.B(n_4035),
.Y(n_4397)
);

NAND3xp33_ASAP7_75t_L g4398 ( 
.A(n_4279),
.B(n_4065),
.C(n_4071),
.Y(n_4398)
);

OR2x2_ASAP7_75t_L g4399 ( 
.A(n_4274),
.B(n_4074),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4286),
.B(n_4077),
.Y(n_4400)
);

AOI221xp5_ASAP7_75t_L g4401 ( 
.A1(n_4342),
.A2(n_4250),
.B1(n_4178),
.B2(n_4264),
.C(n_4240),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4289),
.B(n_4325),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4305),
.Y(n_4403)
);

OA21x2_ASAP7_75t_L g4404 ( 
.A1(n_4328),
.A2(n_4124),
.B(n_4131),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4282),
.B(n_4113),
.Y(n_4405)
);

INVxp67_ASAP7_75t_SL g4406 ( 
.A(n_4284),
.Y(n_4406)
);

AOI221xp5_ASAP7_75t_L g4407 ( 
.A1(n_4347),
.A2(n_4253),
.B1(n_4221),
.B2(n_4225),
.C(n_4142),
.Y(n_4407)
);

OA21x2_ASAP7_75t_L g4408 ( 
.A1(n_4328),
.A2(n_4072),
.B(n_4068),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_4284),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_4299),
.Y(n_4410)
);

INVxp67_ASAP7_75t_L g4411 ( 
.A(n_4327),
.Y(n_4411)
);

NOR2xp33_ASAP7_75t_L g4412 ( 
.A(n_4278),
.B(n_4294),
.Y(n_4412)
);

OAI22xp5_ASAP7_75t_L g4413 ( 
.A1(n_4345),
.A2(n_4097),
.B1(n_4088),
.B2(n_4259),
.Y(n_4413)
);

AOI22xp33_ASAP7_75t_SL g4414 ( 
.A1(n_4358),
.A2(n_4088),
.B1(n_4102),
.B2(n_4120),
.Y(n_4414)
);

INVx1_ASAP7_75t_SL g4415 ( 
.A(n_4334),
.Y(n_4415)
);

AOI22xp5_ASAP7_75t_L g4416 ( 
.A1(n_4341),
.A2(n_4207),
.B1(n_4011),
.B2(n_4185),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4299),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4301),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_4301),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_4341),
.A2(n_4067),
.B1(n_4150),
.B2(n_4158),
.Y(n_4420)
);

OAI21x1_ASAP7_75t_L g4421 ( 
.A1(n_4330),
.A2(n_4134),
.B(n_4128),
.Y(n_4421)
);

OR2x2_ASAP7_75t_L g4422 ( 
.A(n_4329),
.B(n_4079),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4302),
.Y(n_4423)
);

OAI33xp33_ASAP7_75t_L g4424 ( 
.A1(n_4352),
.A2(n_4144),
.A3(n_4161),
.B1(n_4146),
.B2(n_4155),
.B3(n_3889),
.Y(n_4424)
);

NOR2xp33_ASAP7_75t_R g4425 ( 
.A(n_4338),
.B(n_3764),
.Y(n_4425)
);

OR2x6_ASAP7_75t_L g4426 ( 
.A(n_4362),
.B(n_3764),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4280),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4287),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4354),
.B(n_3945),
.Y(n_4429)
);

NAND3xp33_ASAP7_75t_L g4430 ( 
.A(n_4350),
.B(n_4356),
.C(n_4351),
.Y(n_4430)
);

NOR2xp33_ASAP7_75t_R g4431 ( 
.A(n_4338),
.B(n_3904),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4302),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4295),
.Y(n_4433)
);

AOI221xp5_ASAP7_75t_L g4434 ( 
.A1(n_4308),
.A2(n_4242),
.B1(n_4147),
.B2(n_4200),
.C(n_4106),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4297),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4318),
.B(n_4060),
.Y(n_4436)
);

AOI21xp33_ASAP7_75t_L g4437 ( 
.A1(n_4337),
.A2(n_4122),
.B(n_3935),
.Y(n_4437)
);

AOI22xp33_ASAP7_75t_L g4438 ( 
.A1(n_4358),
.A2(n_4066),
.B1(n_4208),
.B2(n_4258),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4320),
.B(n_4114),
.Y(n_4439)
);

AOI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_4349),
.A2(n_4288),
.B1(n_4364),
.B2(n_4355),
.Y(n_4440)
);

OAI22xp5_ASAP7_75t_SL g4441 ( 
.A1(n_4338),
.A2(n_3969),
.B1(n_3973),
.B2(n_3943),
.Y(n_4441)
);

BUFx3_ASAP7_75t_L g4442 ( 
.A(n_4362),
.Y(n_4442)
);

NAND3xp33_ASAP7_75t_L g4443 ( 
.A(n_4350),
.B(n_4099),
.C(n_4108),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4310),
.Y(n_4444)
);

INVx3_ASAP7_75t_L g4445 ( 
.A(n_4281),
.Y(n_4445)
);

AO21x2_ASAP7_75t_L g4446 ( 
.A1(n_4361),
.A2(n_4117),
.B(n_4105),
.Y(n_4446)
);

AOI31xp33_ASAP7_75t_L g4447 ( 
.A1(n_4357),
.A2(n_4171),
.A3(n_4193),
.B(n_3799),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4397),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4402),
.B(n_4343),
.Y(n_4449)
);

OR2x2_ASAP7_75t_L g4450 ( 
.A(n_4385),
.B(n_4319),
.Y(n_4450)
);

AOI211x1_ASAP7_75t_SL g4451 ( 
.A1(n_4384),
.A2(n_4363),
.B(n_4361),
.C(n_4330),
.Y(n_4451)
);

AOI22xp33_ASAP7_75t_L g4452 ( 
.A1(n_4387),
.A2(n_4365),
.B1(n_4321),
.B2(n_4332),
.Y(n_4452)
);

INVx2_ASAP7_75t_L g4453 ( 
.A(n_4383),
.Y(n_4453)
);

INVx2_ASAP7_75t_SL g4454 ( 
.A(n_4390),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4369),
.Y(n_4455)
);

HB1xp67_ASAP7_75t_L g4456 ( 
.A(n_4406),
.Y(n_4456)
);

INVx2_ASAP7_75t_L g4457 ( 
.A(n_4369),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4400),
.B(n_4343),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4422),
.B(n_4339),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4378),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4379),
.Y(n_4461)
);

OAI321xp33_ASAP7_75t_L g4462 ( 
.A1(n_4396),
.A2(n_4353),
.A3(n_4344),
.B1(n_4098),
.B2(n_4326),
.C(n_4363),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4409),
.B(n_4344),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4375),
.B(n_4314),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4440),
.B(n_4296),
.Y(n_4465)
);

OR2x2_ASAP7_75t_L g4466 ( 
.A(n_4381),
.B(n_4340),
.Y(n_4466)
);

AND2x2_ASAP7_75t_L g4467 ( 
.A(n_4371),
.B(n_4293),
.Y(n_4467)
);

INVx2_ASAP7_75t_SL g4468 ( 
.A(n_4426),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_4382),
.B(n_4293),
.Y(n_4469)
);

NAND3xp33_ASAP7_75t_L g4470 ( 
.A(n_4443),
.B(n_4356),
.C(n_4359),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4403),
.B(n_4322),
.Y(n_4471)
);

INVxp67_ASAP7_75t_SL g4472 ( 
.A(n_4395),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4392),
.Y(n_4473)
);

AND2x2_ASAP7_75t_L g4474 ( 
.A(n_4412),
.B(n_4405),
.Y(n_4474)
);

OR2x2_ASAP7_75t_L g4475 ( 
.A(n_4388),
.B(n_4336),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4408),
.B(n_4307),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4427),
.Y(n_4477)
);

AND2x2_ASAP7_75t_L g4478 ( 
.A(n_4408),
.B(n_4307),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4428),
.Y(n_4479)
);

OR2x2_ASAP7_75t_L g4480 ( 
.A(n_4386),
.B(n_4436),
.Y(n_4480)
);

AND2x2_ASAP7_75t_L g4481 ( 
.A(n_4399),
.B(n_4307),
.Y(n_4481)
);

INVx2_ASAP7_75t_SL g4482 ( 
.A(n_4426),
.Y(n_4482)
);

HB1xp67_ASAP7_75t_L g4483 ( 
.A(n_4444),
.Y(n_4483)
);

AND2x2_ASAP7_75t_L g4484 ( 
.A(n_4439),
.B(n_4307),
.Y(n_4484)
);

INVx3_ASAP7_75t_L g4485 ( 
.A(n_4442),
.Y(n_4485)
);

AND2x2_ASAP7_75t_L g4486 ( 
.A(n_4429),
.B(n_4283),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4421),
.B(n_4433),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4435),
.B(n_4283),
.Y(n_4488)
);

AND2x2_ASAP7_75t_L g4489 ( 
.A(n_4444),
.B(n_4410),
.Y(n_4489)
);

NAND2x1_ASAP7_75t_SL g4490 ( 
.A(n_4394),
.B(n_4445),
.Y(n_4490)
);

NOR2xp33_ASAP7_75t_L g4491 ( 
.A(n_4415),
.B(n_4300),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4417),
.B(n_4418),
.Y(n_4492)
);

OR2x2_ASAP7_75t_L g4493 ( 
.A(n_4419),
.B(n_4306),
.Y(n_4493)
);

OR2x2_ASAP7_75t_L g4494 ( 
.A(n_4423),
.B(n_4306),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4432),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4446),
.Y(n_4496)
);

AND2x2_ASAP7_75t_L g4497 ( 
.A(n_4445),
.B(n_4290),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4446),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4411),
.B(n_4430),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_4398),
.B(n_4314),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4404),
.Y(n_4501)
);

INVx2_ASAP7_75t_L g4502 ( 
.A(n_4404),
.Y(n_4502)
);

INVx1_ASAP7_75t_SL g4503 ( 
.A(n_4393),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4380),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4414),
.B(n_4290),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4413),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4391),
.Y(n_4507)
);

CKINVDCx16_ASAP7_75t_R g4508 ( 
.A(n_4431),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4391),
.Y(n_4509)
);

AND2x4_ASAP7_75t_L g4510 ( 
.A(n_4391),
.B(n_4281),
.Y(n_4510)
);

OR2x2_ASAP7_75t_L g4511 ( 
.A(n_4420),
.B(n_4269),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_4441),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_4425),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4416),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4370),
.Y(n_4515)
);

HB1xp67_ASAP7_75t_L g4516 ( 
.A(n_4434),
.Y(n_4516)
);

AND2x4_ASAP7_75t_L g4517 ( 
.A(n_4468),
.B(n_4285),
.Y(n_4517)
);

INVx1_ASAP7_75t_SL g4518 ( 
.A(n_4454),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4450),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4481),
.B(n_4304),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4453),
.Y(n_4521)
);

INVxp67_ASAP7_75t_SL g4522 ( 
.A(n_4456),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_4481),
.B(n_4309),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4464),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4474),
.B(n_4348),
.Y(n_4525)
);

AND2x4_ASAP7_75t_L g4526 ( 
.A(n_4468),
.B(n_4285),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4460),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_4475),
.Y(n_4528)
);

INVx2_ASAP7_75t_L g4529 ( 
.A(n_4453),
.Y(n_4529)
);

BUFx2_ASAP7_75t_SL g4530 ( 
.A(n_4482),
.Y(n_4530)
);

OR2x2_ASAP7_75t_L g4531 ( 
.A(n_4448),
.B(n_4368),
.Y(n_4531)
);

NAND2xp5_ASAP7_75t_L g4532 ( 
.A(n_4484),
.B(n_4312),
.Y(n_4532)
);

AOI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_4513),
.A2(n_4447),
.B(n_4376),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4461),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4473),
.Y(n_4535)
);

AND2x2_ASAP7_75t_L g4536 ( 
.A(n_4474),
.B(n_4290),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4477),
.Y(n_4537)
);

OR2x6_ASAP7_75t_L g4538 ( 
.A(n_4482),
.B(n_4366),
.Y(n_4538)
);

INVx3_ASAP7_75t_L g4539 ( 
.A(n_4485),
.Y(n_4539)
);

BUFx3_ASAP7_75t_L g4540 ( 
.A(n_4454),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_L g4541 ( 
.A(n_4484),
.B(n_4313),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4511),
.B(n_4317),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4514),
.B(n_4310),
.Y(n_4543)
);

AOI21xp33_ASAP7_75t_SL g4544 ( 
.A1(n_4508),
.A2(n_4437),
.B(n_4374),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_4483),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4479),
.Y(n_4546)
);

OAI21xp33_ASAP7_75t_L g4547 ( 
.A1(n_4476),
.A2(n_4377),
.B(n_4373),
.Y(n_4547)
);

INVxp67_ASAP7_75t_SL g4548 ( 
.A(n_4485),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4506),
.B(n_4311),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4500),
.B(n_4311),
.Y(n_4550)
);

INVx1_ASAP7_75t_SL g4551 ( 
.A(n_4485),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4448),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4472),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4458),
.B(n_4269),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4489),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4458),
.B(n_4277),
.Y(n_4556)
);

AND2x2_ASAP7_75t_L g4557 ( 
.A(n_4486),
.B(n_4277),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4451),
.B(n_4292),
.Y(n_4558)
);

OAI21xp5_ASAP7_75t_L g4559 ( 
.A1(n_4516),
.A2(n_4372),
.B(n_4438),
.Y(n_4559)
);

INVxp67_ASAP7_75t_SL g4560 ( 
.A(n_4501),
.Y(n_4560)
);

INVx4_ASAP7_75t_L g4561 ( 
.A(n_4510),
.Y(n_4561)
);

NOR2xp33_ASAP7_75t_R g4562 ( 
.A(n_4539),
.B(n_4512),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_L g4563 ( 
.A(n_4547),
.B(n_4515),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4530),
.B(n_4548),
.Y(n_4564)
);

INVxp67_ASAP7_75t_L g4565 ( 
.A(n_4533),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_SL g4566 ( 
.A(n_4539),
.B(n_4462),
.Y(n_4566)
);

AO22x1_ASAP7_75t_L g4567 ( 
.A1(n_4551),
.A2(n_4505),
.B1(n_4503),
.B2(n_4499),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4549),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4522),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4553),
.Y(n_4570)
);

OR2x2_ASAP7_75t_L g4571 ( 
.A(n_4532),
.B(n_4480),
.Y(n_4571)
);

AND2x2_ASAP7_75t_L g4572 ( 
.A(n_4540),
.B(n_4499),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4551),
.B(n_4487),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4532),
.B(n_4515),
.Y(n_4574)
);

CKINVDCx5p33_ASAP7_75t_R g4575 ( 
.A(n_4538),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4538),
.B(n_4517),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_4541),
.B(n_4520),
.Y(n_4577)
);

HB1xp67_ASAP7_75t_L g4578 ( 
.A(n_4518),
.Y(n_4578)
);

AND2x4_ASAP7_75t_L g4579 ( 
.A(n_4538),
.B(n_4504),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4543),
.Y(n_4580)
);

NOR2xp33_ASAP7_75t_L g4581 ( 
.A(n_4544),
.B(n_4459),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4528),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4524),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4560),
.Y(n_4584)
);

INVx1_ASAP7_75t_SL g4585 ( 
.A(n_4518),
.Y(n_4585)
);

BUFx3_ASAP7_75t_L g4586 ( 
.A(n_4517),
.Y(n_4586)
);

NAND2xp33_ASAP7_75t_R g4587 ( 
.A(n_4559),
.B(n_4505),
.Y(n_4587)
);

AND2x4_ASAP7_75t_L g4588 ( 
.A(n_4526),
.B(n_4487),
.Y(n_4588)
);

OR2x2_ASAP7_75t_L g4589 ( 
.A(n_4541),
.B(n_4466),
.Y(n_4589)
);

AND2x2_ASAP7_75t_L g4590 ( 
.A(n_4526),
.B(n_4465),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4555),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4561),
.B(n_4465),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4542),
.B(n_4452),
.Y(n_4593)
);

NOR4xp25_ASAP7_75t_SL g4594 ( 
.A(n_4519),
.B(n_4507),
.C(n_4509),
.D(n_4407),
.Y(n_4594)
);

NAND2x1p5_ASAP7_75t_L g4595 ( 
.A(n_4561),
.B(n_4510),
.Y(n_4595)
);

OAI21xp5_ASAP7_75t_L g4596 ( 
.A1(n_4559),
.A2(n_4470),
.B(n_4452),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4521),
.Y(n_4597)
);

AND3x2_ASAP7_75t_L g4598 ( 
.A(n_4536),
.B(n_4491),
.C(n_4478),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4534),
.Y(n_4599)
);

NOR2xp33_ASAP7_75t_R g4600 ( 
.A(n_4525),
.B(n_3955),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4557),
.B(n_4488),
.Y(n_4601)
);

OR2x6_ASAP7_75t_L g4602 ( 
.A(n_4558),
.B(n_4490),
.Y(n_4602)
);

NOR3xp33_ASAP7_75t_L g4603 ( 
.A(n_4558),
.B(n_4424),
.C(n_4476),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4520),
.B(n_4488),
.Y(n_4604)
);

NAND4xp25_ASAP7_75t_L g4605 ( 
.A(n_4542),
.B(n_4401),
.C(n_4389),
.D(n_4478),
.Y(n_4605)
);

AND2x2_ASAP7_75t_L g4606 ( 
.A(n_4523),
.B(n_4486),
.Y(n_4606)
);

OR2x2_ASAP7_75t_L g4607 ( 
.A(n_4523),
.B(n_4550),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4535),
.Y(n_4608)
);

OR2x2_ASAP7_75t_L g4609 ( 
.A(n_4550),
.B(n_4493),
.Y(n_4609)
);

OAI32xp33_ASAP7_75t_L g4610 ( 
.A1(n_4587),
.A2(n_4491),
.A3(n_4502),
.B1(n_4545),
.B2(n_4552),
.Y(n_4610)
);

AOI22xp33_ASAP7_75t_L g4611 ( 
.A1(n_4581),
.A2(n_4502),
.B1(n_4497),
.B2(n_4527),
.Y(n_4611)
);

NOR2xp33_ASAP7_75t_L g4612 ( 
.A(n_4575),
.B(n_4537),
.Y(n_4612)
);

OAI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4565),
.A2(n_4531),
.B1(n_4529),
.B2(n_4546),
.Y(n_4613)
);

AOI221xp5_ASAP7_75t_L g4614 ( 
.A1(n_4596),
.A2(n_4497),
.B1(n_4496),
.B2(n_4498),
.C(n_4457),
.Y(n_4614)
);

NOR2xp33_ASAP7_75t_R g4615 ( 
.A(n_4564),
.B(n_3955),
.Y(n_4615)
);

NOR3xp33_ASAP7_75t_SL g4616 ( 
.A(n_4596),
.B(n_4232),
.C(n_4222),
.Y(n_4616)
);

XOR2xp5_ASAP7_75t_L g4617 ( 
.A(n_4563),
.B(n_4510),
.Y(n_4617)
);

AOI21xp5_ASAP7_75t_L g4618 ( 
.A1(n_4567),
.A2(n_4457),
.B(n_4455),
.Y(n_4618)
);

OAI22xp5_ASAP7_75t_L g4619 ( 
.A1(n_4593),
.A2(n_4449),
.B1(n_4556),
.B2(n_4554),
.Y(n_4619)
);

OAI21xp5_ASAP7_75t_L g4620 ( 
.A1(n_4585),
.A2(n_4203),
.B(n_4496),
.Y(n_4620)
);

OAI22xp5_ASAP7_75t_L g4621 ( 
.A1(n_4595),
.A2(n_4449),
.B1(n_4469),
.B2(n_4467),
.Y(n_4621)
);

OAI22xp5_ASAP7_75t_L g4622 ( 
.A1(n_4586),
.A2(n_4469),
.B1(n_4467),
.B2(n_4455),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4569),
.Y(n_4623)
);

OAI22xp5_ASAP7_75t_L g4624 ( 
.A1(n_4579),
.A2(n_4471),
.B1(n_4463),
.B2(n_4494),
.Y(n_4624)
);

OR2x2_ASAP7_75t_L g4625 ( 
.A(n_4607),
.B(n_4495),
.Y(n_4625)
);

OAI321xp33_ASAP7_75t_L g4626 ( 
.A1(n_4605),
.A2(n_4498),
.A3(n_4168),
.B1(n_4198),
.B2(n_4201),
.C(n_4141),
.Y(n_4626)
);

OAI22xp5_ASAP7_75t_L g4627 ( 
.A1(n_4579),
.A2(n_4471),
.B1(n_4463),
.B2(n_4489),
.Y(n_4627)
);

NAND3xp33_ASAP7_75t_L g4628 ( 
.A(n_4603),
.B(n_4215),
.C(n_4156),
.Y(n_4628)
);

NOR2xp33_ASAP7_75t_L g4629 ( 
.A(n_4605),
.B(n_4492),
.Y(n_4629)
);

OAI211xp5_ASAP7_75t_L g4630 ( 
.A1(n_4562),
.A2(n_4236),
.B(n_4231),
.C(n_4249),
.Y(n_4630)
);

AOI22xp33_ASAP7_75t_SL g4631 ( 
.A1(n_4576),
.A2(n_4303),
.B1(n_4036),
.B2(n_4265),
.Y(n_4631)
);

OAI211xp5_ASAP7_75t_SL g4632 ( 
.A1(n_4566),
.A2(n_4247),
.B(n_4089),
.C(n_4164),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4585),
.B(n_4492),
.Y(n_4633)
);

OAI22xp5_ASAP7_75t_L g4634 ( 
.A1(n_4574),
.A2(n_4083),
.B1(n_4316),
.B2(n_3991),
.Y(n_4634)
);

NAND4xp25_ASAP7_75t_L g4635 ( 
.A(n_4572),
.B(n_4239),
.C(n_3967),
.D(n_4109),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4578),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4609),
.Y(n_4637)
);

NOR2xp33_ASAP7_75t_L g4638 ( 
.A(n_4584),
.B(n_4303),
.Y(n_4638)
);

OAI22xp5_ASAP7_75t_L g4639 ( 
.A1(n_4592),
.A2(n_4036),
.B1(n_4090),
.B2(n_4123),
.Y(n_4639)
);

OAI32xp33_ASAP7_75t_L g4640 ( 
.A1(n_4594),
.A2(n_4001),
.A3(n_4027),
.B1(n_3763),
.B2(n_3902),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4597),
.Y(n_4641)
);

AOI221xp5_ASAP7_75t_L g4642 ( 
.A1(n_4629),
.A2(n_4570),
.B1(n_4583),
.B2(n_4582),
.C(n_4580),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4636),
.B(n_4604),
.Y(n_4643)
);

OAI21xp5_ASAP7_75t_L g4644 ( 
.A1(n_4626),
.A2(n_4602),
.B(n_4573),
.Y(n_4644)
);

OAI21xp33_ASAP7_75t_L g4645 ( 
.A1(n_4611),
.A2(n_4602),
.B(n_4600),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4637),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4616),
.B(n_4606),
.Y(n_4647)
);

OAI32xp33_ASAP7_75t_L g4648 ( 
.A1(n_4617),
.A2(n_4594),
.A3(n_4577),
.B1(n_4571),
.B2(n_4590),
.Y(n_4648)
);

OR2x2_ASAP7_75t_L g4649 ( 
.A(n_4633),
.B(n_4589),
.Y(n_4649)
);

OR2x2_ASAP7_75t_L g4650 ( 
.A(n_4623),
.B(n_4568),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4612),
.B(n_4608),
.Y(n_4651)
);

OAI22xp5_ASAP7_75t_L g4652 ( 
.A1(n_4621),
.A2(n_4602),
.B1(n_4588),
.B2(n_4599),
.Y(n_4652)
);

NOR3xp33_ASAP7_75t_L g4653 ( 
.A(n_4626),
.B(n_4180),
.C(n_3921),
.Y(n_4653)
);

AOI221xp5_ASAP7_75t_SL g4654 ( 
.A1(n_4610),
.A2(n_4591),
.B1(n_4598),
.B2(n_4601),
.C(n_3898),
.Y(n_4654)
);

INVx1_ASAP7_75t_SL g4655 ( 
.A(n_4615),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4625),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4613),
.Y(n_4657)
);

AOI22xp33_ASAP7_75t_L g4658 ( 
.A1(n_4639),
.A2(n_4588),
.B1(n_4359),
.B2(n_4360),
.Y(n_4658)
);

AND2x4_ASAP7_75t_L g4659 ( 
.A(n_4641),
.B(n_4620),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_L g4660 ( 
.A(n_4628),
.B(n_4166),
.Y(n_4660)
);

AOI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_4632),
.A2(n_4206),
.B1(n_4166),
.B2(n_4248),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4614),
.B(n_4206),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4634),
.B(n_4360),
.Y(n_4663)
);

AOI22xp33_ASAP7_75t_L g4664 ( 
.A1(n_4631),
.A2(n_4248),
.B1(n_4041),
.B2(n_4032),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4619),
.Y(n_4665)
);

NOR2xp33_ASAP7_75t_L g4666 ( 
.A(n_4640),
.B(n_4622),
.Y(n_4666)
);

CKINVDCx5p33_ASAP7_75t_R g4667 ( 
.A(n_4655),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4657),
.B(n_4627),
.Y(n_4668)
);

AOI21xp5_ASAP7_75t_L g4669 ( 
.A1(n_4648),
.A2(n_4618),
.B(n_4638),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4646),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4665),
.B(n_4624),
.Y(n_4671)
);

XOR2x2_ASAP7_75t_L g4672 ( 
.A(n_4647),
.B(n_4630),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4642),
.B(n_4635),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4656),
.B(n_4292),
.Y(n_4674)
);

NOR2xp33_ASAP7_75t_L g4675 ( 
.A(n_4645),
.B(n_3763),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4649),
.Y(n_4676)
);

NAND3xp33_ASAP7_75t_L g4677 ( 
.A(n_4644),
.B(n_4188),
.C(n_4173),
.Y(n_4677)
);

HB1xp67_ASAP7_75t_L g4678 ( 
.A(n_4651),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4652),
.B(n_4053),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4650),
.Y(n_4680)
);

INVx1_ASAP7_75t_SL g4681 ( 
.A(n_4659),
.Y(n_4681)
);

NAND2xp33_ASAP7_75t_SL g4682 ( 
.A(n_4660),
.B(n_4019),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4643),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4653),
.B(n_4016),
.Y(n_4684)
);

AND2x2_ASAP7_75t_L g4685 ( 
.A(n_4666),
.B(n_4659),
.Y(n_4685)
);

INVx1_ASAP7_75t_L g4686 ( 
.A(n_4662),
.Y(n_4686)
);

NOR2xp33_ASAP7_75t_L g4687 ( 
.A(n_4663),
.B(n_748),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4661),
.Y(n_4688)
);

AOI21xp5_ASAP7_75t_L g4689 ( 
.A1(n_4667),
.A2(n_4658),
.B(n_4664),
.Y(n_4689)
);

NOR3xp33_ASAP7_75t_L g4690 ( 
.A(n_4681),
.B(n_4654),
.C(n_3992),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4676),
.Y(n_4691)
);

NOR5xp2_ASAP7_75t_L g4692 ( 
.A(n_4678),
.B(n_4686),
.C(n_4688),
.D(n_4670),
.E(n_4683),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4668),
.B(n_748),
.Y(n_4693)
);

XNOR2x2_ASAP7_75t_L g4694 ( 
.A(n_4672),
.B(n_3971),
.Y(n_4694)
);

AOI21xp33_ASAP7_75t_SL g4695 ( 
.A1(n_4687),
.A2(n_749),
.B(n_751),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4680),
.Y(n_4696)
);

NOR3xp33_ASAP7_75t_L g4697 ( 
.A(n_4675),
.B(n_4006),
.C(n_4047),
.Y(n_4697)
);

NOR3xp33_ASAP7_75t_L g4698 ( 
.A(n_4687),
.B(n_4050),
.C(n_4047),
.Y(n_4698)
);

NAND3xp33_ASAP7_75t_L g4699 ( 
.A(n_4669),
.B(n_4678),
.C(n_4685),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_SL g4700 ( 
.A(n_4669),
.B(n_4044),
.Y(n_4700)
);

INVxp67_ASAP7_75t_L g4701 ( 
.A(n_4684),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4671),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_SL g4703 ( 
.A(n_4673),
.B(n_4044),
.Y(n_4703)
);

OAI211xp5_ASAP7_75t_L g4704 ( 
.A1(n_4699),
.A2(n_4679),
.B(n_4677),
.C(n_4682),
.Y(n_4704)
);

AOI21xp5_ASAP7_75t_L g4705 ( 
.A1(n_4700),
.A2(n_4674),
.B(n_4050),
.Y(n_4705)
);

OAI21xp33_ASAP7_75t_SL g4706 ( 
.A1(n_4703),
.A2(n_4092),
.B(n_4148),
.Y(n_4706)
);

AOI211x1_ASAP7_75t_L g4707 ( 
.A1(n_4689),
.A2(n_3814),
.B(n_4139),
.C(n_753),
.Y(n_4707)
);

AOI32xp33_ASAP7_75t_L g4708 ( 
.A1(n_4690),
.A2(n_4021),
.A3(n_3860),
.B1(n_3815),
.B2(n_3865),
.Y(n_4708)
);

NAND3xp33_ASAP7_75t_SL g4709 ( 
.A(n_4692),
.B(n_4121),
.C(n_751),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4702),
.B(n_4696),
.Y(n_4710)
);

AOI221xp5_ASAP7_75t_L g4711 ( 
.A1(n_4691),
.A2(n_4104),
.B1(n_3910),
.B2(n_3905),
.C(n_3911),
.Y(n_4711)
);

OAI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4693),
.A2(n_4005),
.B(n_3929),
.Y(n_4712)
);

OAI21xp5_ASAP7_75t_L g4713 ( 
.A1(n_4701),
.A2(n_4695),
.B(n_4697),
.Y(n_4713)
);

OAI221xp5_ASAP7_75t_SL g4714 ( 
.A1(n_4694),
.A2(n_4041),
.B1(n_4032),
.B2(n_3743),
.C(n_3890),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4698),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4710),
.Y(n_4716)
);

CKINVDCx5p33_ASAP7_75t_R g4717 ( 
.A(n_4709),
.Y(n_4717)
);

HB1xp67_ASAP7_75t_L g4718 ( 
.A(n_4715),
.Y(n_4718)
);

NOR2xp33_ASAP7_75t_R g4719 ( 
.A(n_4713),
.B(n_752),
.Y(n_4719)
);

AOI222xp33_ASAP7_75t_L g4720 ( 
.A1(n_4706),
.A2(n_3743),
.B1(n_3794),
.B2(n_3769),
.C1(n_3745),
.C2(n_3760),
.Y(n_4720)
);

AOI22xp33_ASAP7_75t_L g4721 ( 
.A1(n_4705),
.A2(n_3834),
.B1(n_3743),
.B2(n_3789),
.Y(n_4721)
);

O2A1O1Ixp33_ASAP7_75t_L g4722 ( 
.A1(n_4704),
.A2(n_4000),
.B(n_755),
.C(n_756),
.Y(n_4722)
);

INVx1_ASAP7_75t_SL g4723 ( 
.A(n_4712),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4717),
.B(n_4711),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4716),
.B(n_4708),
.Y(n_4725)
);

AOI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4718),
.A2(n_4714),
.B(n_4707),
.Y(n_4726)
);

NAND4xp25_ASAP7_75t_L g4727 ( 
.A(n_4725),
.B(n_4726),
.C(n_4724),
.D(n_4722),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_SL g4728 ( 
.A(n_4726),
.B(n_4719),
.Y(n_4728)
);

OAI22xp33_ASAP7_75t_SL g4729 ( 
.A1(n_4725),
.A2(n_4723),
.B1(n_4720),
.B2(n_4721),
.Y(n_4729)
);

CKINVDCx5p33_ASAP7_75t_R g4730 ( 
.A(n_4728),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_4730),
.A2(n_4727),
.B(n_4729),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4731),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4732),
.Y(n_4733)
);

AOI21xp33_ASAP7_75t_L g4734 ( 
.A1(n_4733),
.A2(n_754),
.B(n_756),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4734),
.Y(n_4735)
);

AOI22xp33_ASAP7_75t_SL g4736 ( 
.A1(n_4735),
.A2(n_3834),
.B1(n_3789),
.B2(n_3880),
.Y(n_4736)
);

OAI221xp5_ASAP7_75t_R g4737 ( 
.A1(n_4736),
.A2(n_3890),
.B1(n_758),
.B2(n_759),
.C(n_760),
.Y(n_4737)
);

AOI211xp5_ASAP7_75t_L g4738 ( 
.A1(n_4737),
.A2(n_3834),
.B(n_3794),
.C(n_3769),
.Y(n_4738)
);


endmodule