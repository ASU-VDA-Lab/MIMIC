module fake_jpeg_9542_n_116 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_29),
.Y(n_48)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_32),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_13),
.B1(n_15),
.B2(n_19),
.Y(n_47)
);

AOI32xp33_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_17),
.A3(n_16),
.B1(n_12),
.B2(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_47),
.B1(n_37),
.B2(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_19),
.B1(n_18),
.B2(n_15),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_61),
.B1(n_63),
.B2(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_9),
.Y(n_79)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_12),
.B1(n_3),
.B2(n_5),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_38),
.B1(n_5),
.B2(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_78),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_48),
.C(n_40),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_55),
.C(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_39),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_61),
.B1(n_60),
.B2(n_65),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_83),
.B1(n_89),
.B2(n_73),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_69),
.B1(n_78),
.B2(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_52),
.B1(n_60),
.B2(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_69),
.B1(n_74),
.B2(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_100)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_7),
.C(n_9),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_93),
.B1(n_89),
.B2(n_83),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_86),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_94),
.C(n_98),
.Y(n_104)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_98),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_91),
.C(n_82),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_97),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_101),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_111),
.B(n_40),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_91),
.C(n_80),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_82),
.A3(n_70),
.B1(n_38),
.B2(n_58),
.C1(n_7),
.C2(n_45),
.Y(n_112)
);

OAI321xp33_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_113),
.A3(n_40),
.B1(n_53),
.B2(n_45),
.C(n_2),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_2),
.B(n_5),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_6),
.Y(n_116)
);


endmodule