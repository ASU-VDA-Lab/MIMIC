module fake_jpeg_25890_n_101 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx11_ASAP7_75t_SL g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_21),
.B1(n_18),
.B2(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_13),
.B1(n_19),
.B2(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_23),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_25),
.A2(n_18),
.B(n_15),
.C(n_13),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_45),
.B1(n_34),
.B2(n_23),
.Y(n_50)
);

AO21x2_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_27),
.B(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_46),
.B1(n_39),
.B2(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_54),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_65)
);

FAx1_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_11),
.CI(n_2),
.CON(n_51),
.SN(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_59),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_19),
.B1(n_14),
.B2(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_5),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_11),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_43),
.B1(n_46),
.B2(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_67),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_55),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_47),
.B(n_9),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_48),
.B(n_51),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_7),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_47),
.B(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_79),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_61),
.C(n_69),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_72),
.C(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_62),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_90),
.B1(n_81),
.B2(n_85),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_76),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_67),
.C(n_70),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_84),
.B1(n_80),
.B2(n_68),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_91),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

NOR2xp67_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_62),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_92),
.C(n_47),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_47),
.Y(n_101)
);


endmodule