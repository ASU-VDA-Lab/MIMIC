module fake_jpeg_28737_n_439 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_439);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_439;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_70),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_75),
.Y(n_84)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_16),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_30),
.Y(n_85)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_15),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_19),
.B(n_0),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_24),
.C(n_20),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_85),
.B(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_89),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_121),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_29),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_117),
.Y(n_130)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_54),
.B(n_30),
.CON(n_111),
.SN(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_64),
.B(n_30),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_32),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_136),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_51),
.B1(n_52),
.B2(n_48),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_137),
.B1(n_143),
.B2(n_73),
.Y(n_184)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_106),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_58),
.B1(n_63),
.B2(n_59),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_28),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_138),
.B(n_162),
.Y(n_193)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_26),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_153),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_43),
.B1(n_53),
.B2(n_56),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_65),
.B1(n_62),
.B2(n_44),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_157),
.B1(n_67),
.B2(n_68),
.Y(n_173)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_26),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_156),
.Y(n_192)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_111),
.A2(n_61),
.B1(n_60),
.B2(n_76),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_161),
.Y(n_189)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_164),
.B1(n_123),
.B2(n_98),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_119),
.CI(n_113),
.CON(n_170),
.SN(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_185),
.B(n_178),
.C(n_187),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_184),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_98),
.B1(n_120),
.B2(n_87),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_178),
.A2(n_182),
.B1(n_185),
.B2(n_188),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_114),
.B(n_118),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_138),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_120),
.B1(n_127),
.B2(n_87),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_133),
.A2(n_127),
.B1(n_99),
.B2(n_92),
.Y(n_185)
);

AOI22x1_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_114),
.B1(n_79),
.B2(n_101),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_182),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_130),
.A2(n_109),
.B1(n_104),
.B2(n_92),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_202),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_198),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_160),
.C(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_209),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_139),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_215),
.C(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_131),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_134),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_218),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_132),
.B1(n_163),
.B2(n_110),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_206),
.B1(n_168),
.B2(n_176),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_155),
.B1(n_149),
.B2(n_150),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_136),
.CI(n_129),
.CON(n_208),
.SN(n_208)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_180),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_190),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_191),
.Y(n_225)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_193),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_213),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_161),
.C(n_148),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_181),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_188),
.B(n_32),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_184),
.B1(n_173),
.B2(n_177),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_225),
.B1(n_207),
.B2(n_204),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_183),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_177),
.B1(n_104),
.B2(n_109),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_223),
.A2(n_226),
.B1(n_180),
.B2(n_198),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_177),
.B1(n_175),
.B2(n_174),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NOR4xp25_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_15),
.C(n_168),
.D(n_2),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_229),
.B(n_197),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_204),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_179),
.B(n_108),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_234),
.B(n_236),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_179),
.B(n_186),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_207),
.B(n_210),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_171),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_215),
.C(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_242),
.A2(n_248),
.B1(n_266),
.B2(n_230),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_195),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_219),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_229),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_244),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_265),
.C(n_227),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_203),
.B(n_208),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_251),
.B(n_229),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_221),
.A2(n_202),
.B1(n_214),
.B2(n_218),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_202),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_261),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_257),
.A2(n_259),
.B1(n_267),
.B2(n_235),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_171),
.B1(n_152),
.B2(n_156),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_183),
.Y(n_260)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_28),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_28),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_169),
.B1(n_147),
.B2(n_90),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_236),
.A2(n_169),
.B1(n_158),
.B2(n_162),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_222),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_280),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_222),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_277),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_220),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_259),
.B1(n_225),
.B2(n_252),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_279),
.A2(n_297),
.B1(n_242),
.B2(n_248),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_220),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_225),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_284),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_234),
.B(n_232),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_224),
.Y(n_283)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_255),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_232),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_290),
.C(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_SL g321 ( 
.A(n_286),
.B(n_257),
.C(n_237),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_287),
.A2(n_257),
.B1(n_246),
.B2(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_291),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_224),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_235),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_240),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_299),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_253),
.C(n_250),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_302),
.B(n_292),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_253),
.C(n_256),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_310),
.C(n_322),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_272),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_306),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_309),
.A2(n_321),
.B1(n_297),
.B2(n_286),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_242),
.C(n_263),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_279),
.A2(n_266),
.B1(n_226),
.B2(n_223),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_314),
.A2(n_309),
.B1(n_321),
.B2(n_298),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_287),
.A2(n_276),
.B1(n_278),
.B2(n_259),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_292),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_316),
.B(n_323),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_318),
.A2(n_295),
.B1(n_296),
.B2(n_271),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_240),
.C(n_237),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_324),
.A2(n_327),
.B1(n_319),
.B2(n_318),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_301),
.B(n_280),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_333),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_339),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_344),
.B1(n_339),
.B2(n_330),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_338),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_290),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_285),
.C(n_281),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_335),
.C(n_337),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_301),
.B(n_295),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_311),
.B(n_288),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_146),
.C(n_141),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_342),
.C(n_347),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_140),
.C(n_264),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_307),
.A2(n_264),
.B1(n_20),
.B2(n_24),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_34),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_315),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_108),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_15),
.B1(n_90),
.B2(n_38),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_303),
.C(n_317),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_350),
.A2(n_355),
.B1(n_338),
.B2(n_341),
.Y(n_372)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_302),
.C(n_319),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_353),
.Y(n_374)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_331),
.Y(n_352)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_356),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_324),
.A2(n_317),
.B1(n_164),
.B2(n_96),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_362),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_359),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_335),
.A2(n_41),
.B1(n_39),
.B2(n_38),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_333),
.B(n_24),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_164),
.C(n_38),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_367),
.C(n_340),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_347),
.B(n_32),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_366),
.A2(n_34),
.B(n_39),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_332),
.B(n_164),
.C(n_39),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_370),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_41),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_342),
.C(n_334),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_371),
.B(n_375),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_373),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_325),
.C(n_337),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_381),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_363),
.C(n_367),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_41),
.C(n_36),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_383),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_36),
.C(n_23),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_36),
.C(n_23),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_386),
.C(n_369),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_23),
.C(n_108),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_100),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_0),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_374),
.A2(n_358),
.B1(n_360),
.B2(n_352),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_392),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_SL g390 ( 
.A(n_385),
.B(n_356),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_390),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_378),
.A2(n_365),
.B1(n_359),
.B2(n_357),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_393),
.A2(n_397),
.B1(n_1),
.B2(n_4),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_34),
.C(n_26),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_373),
.C(n_384),
.Y(n_403)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_395),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_398),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_386),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_402),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_406),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_376),
.B1(n_4),
.B2(n_5),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_405),
.B(n_410),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_1),
.C(n_5),
.Y(n_409)
);

OAI21xp33_ASAP7_75t_L g420 ( 
.A1(n_409),
.A2(n_412),
.B(n_401),
.Y(n_420)
);

OAI22x1_ASAP7_75t_L g410 ( 
.A1(n_396),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_5),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_411),
.B(n_8),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_6),
.C(n_7),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_405),
.B(n_400),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_415),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_395),
.Y(n_415)
);

A2O1A1O1Ixp25_ASAP7_75t_L g416 ( 
.A1(n_404),
.A2(n_394),
.B(n_397),
.C(n_9),
.D(n_10),
.Y(n_416)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_7),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_419),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_10),
.Y(n_429)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_420),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_407),
.A2(n_8),
.B(n_10),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_422),
.B(n_14),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_425),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_421),
.B(n_8),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_426),
.Y(n_431)
);

AOI322xp5_ASAP7_75t_L g433 ( 
.A1(n_429),
.A2(n_413),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_10),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_SL g432 ( 
.A(n_427),
.B(n_417),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_432),
.A2(n_428),
.B(n_423),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_13),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g436 ( 
.A1(n_434),
.A2(n_435),
.B(n_430),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_431),
.C(n_12),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_11),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_13),
.B(n_11),
.Y(n_439)
);


endmodule