module fake_jpeg_11742_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_19),
.B(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_7),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_26),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_19),
.B1(n_15),
.B2(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_15),
.B1(n_20),
.B2(n_24),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_70),
.Y(n_88)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_18),
.Y(n_67)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_69),
.Y(n_82)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_25),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_55),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_42),
.B1(n_48),
.B2(n_52),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_12),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_72),
.C(n_17),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_35),
.B1(n_25),
.B2(n_17),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_77),
.B1(n_69),
.B2(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_22),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_57),
.B(n_16),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_76),
.B(n_55),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_94),
.C(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_102),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_83),
.B(n_91),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_105),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_83),
.B(n_85),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_78),
.B(n_79),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_89),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_110),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_98),
.B(n_99),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_98),
.B1(n_73),
.B2(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_93),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_107),
.C(n_8),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_73),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_121),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_7),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_119),
.A2(n_112),
.B(n_10),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_120),
.B(n_10),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_118),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_126),
.B(n_123),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_30),
.B(n_38),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_38),
.Y(n_129)
);


endmodule