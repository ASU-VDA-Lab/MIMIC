module real_jpeg_14457_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_25),
.C(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_4),
.B(n_43),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_4),
.B(n_23),
.C(n_29),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_48),
.C(n_58),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_102),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_100),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_84),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_14),
.B(n_84),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_65),
.C(n_72),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_15),
.A2(n_16),
.B1(n_65),
.B2(n_66),
.Y(n_180)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_45),
.B2(n_64),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_17),
.A2(n_18),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_17),
.A2(n_18),
.B1(n_75),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_33),
.B2(n_44),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_44),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_19),
.A2(n_20),
.B1(n_56),
.B2(n_67),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_19),
.B(n_79),
.C(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_19),
.A2(n_20),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_20),
.B(n_67),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_20),
.A2(n_67),
.B(n_129),
.C(n_134),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_31),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

OA22x2_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_24),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_25),
.B(n_133),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_28),
.Y(n_152)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_29),
.A2(n_30),
.B1(n_58),
.B2(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_29),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_32),
.B(n_97),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_32),
.B(n_51),
.Y(n_160)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_33),
.A2(n_44),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI211xp5_ASAP7_75t_SL g116 ( 
.A1(n_44),
.A2(n_56),
.B(n_83),
.C(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_45),
.A2(n_74),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_56),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_46),
.A2(n_56),
.B1(n_67),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_51),
.B1(n_54),
.B2(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_49),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_49),
.B(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_56),
.A2(n_67),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_56),
.A2(n_67),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_56),
.A2(n_67),
.B1(n_146),
.B2(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_56),
.B(n_79),
.C(n_150),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_56),
.B(n_136),
.C(n_140),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_63),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_67),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_72),
.A2(n_73),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_82),
.Y(n_73)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_80),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_79),
.A2(n_80),
.B1(n_111),
.B2(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_79),
.B(n_131),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_79),
.A2(n_80),
.B1(n_149),
.B2(n_153),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_79),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_79),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_80),
.B(n_162),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_99),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_87),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_98),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_123),
.B(n_176),
.C(n_181),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_113),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_105),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_107),
.B1(n_129),
.B2(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_115),
.B(n_119),
.C(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_170),
.B(n_175),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_142),
.B(n_169),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_165),
.B(n_168),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_154),
.B(n_164),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);


endmodule