module fake_jpeg_13493_n_526 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_4),
.B(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_62),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_74),
.B(n_110),
.Y(n_159)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_77),
.B(n_93),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g179 ( 
.A(n_80),
.Y(n_179)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_86),
.Y(n_124)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_34),
.B(n_16),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g161 ( 
.A(n_94),
.Y(n_161)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_22),
.Y(n_101)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_16),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_109),
.Y(n_133)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_108),
.Y(n_172)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_38),
.B(n_15),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_111),
.Y(n_196)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_59),
.B1(n_32),
.B2(n_26),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_34),
.B(n_13),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_116),
.Y(n_176)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_53),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_37),
.Y(n_181)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_122),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_138),
.B(n_148),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_81),
.A2(n_59),
.B1(n_42),
.B2(n_41),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_178),
.B1(n_186),
.B2(n_194),
.Y(n_203)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_53),
.B1(n_36),
.B2(n_29),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_150),
.A2(n_179),
.B(n_189),
.C(n_127),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_80),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_154),
.B(n_158),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_94),
.A2(n_32),
.B(n_26),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_156),
.B(n_23),
.C(n_2),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_93),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_77),
.A2(n_114),
.B1(n_48),
.B2(n_38),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_192),
.B1(n_28),
.B2(n_26),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_113),
.B(n_48),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_183),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_105),
.A2(n_59),
.B1(n_42),
.B2(n_41),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_43),
.B1(n_28),
.B2(n_27),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_103),
.A2(n_37),
.B1(n_36),
.B2(n_39),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_27),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_40),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_68),
.A2(n_111),
.B1(n_90),
.B2(n_112),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_40),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_190),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_60),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_62),
.B(n_35),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_115),
.A2(n_35),
.B1(n_54),
.B2(n_30),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_67),
.B(n_54),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_71),
.A2(n_58),
.B1(n_52),
.B2(n_44),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_73),
.B(n_43),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_157),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_76),
.A2(n_58),
.B1(n_52),
.B2(n_44),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_162),
.B1(n_186),
.B2(n_142),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_198),
.Y(n_314)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_110),
.A3(n_100),
.B1(n_99),
.B2(n_89),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_199),
.B(n_206),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_200),
.B(n_204),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_202),
.B(n_213),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_161),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_205),
.A2(n_220),
.B1(n_223),
.B2(n_251),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_144),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_85),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_207),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_209),
.B(n_217),
.Y(n_275)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_84),
.B1(n_79),
.B2(n_78),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_212),
.A2(n_243),
.B1(n_221),
.B2(n_225),
.Y(n_304)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_214),
.Y(n_281)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_155),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_156),
.A2(n_26),
.B1(n_23),
.B2(n_3),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_219),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_149),
.A2(n_26),
.B1(n_23),
.B2(n_13),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_23),
.B1(n_2),
.B2(n_5),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_125),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_224),
.B(n_235),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_225),
.A2(n_262),
.B(n_179),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_152),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_226),
.Y(n_279)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_229),
.Y(n_299)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_179),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_231),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_124),
.B(n_1),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_232),
.B(n_246),
.Y(n_273)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_126),
.B(n_1),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_233),
.Y(n_270)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_128),
.Y(n_234)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_134),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_130),
.Y(n_236)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_152),
.A2(n_1),
.B1(n_6),
.B2(n_7),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_237),
.B(n_238),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_136),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_240),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_178),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_241),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_242),
.B(n_249),
.Y(n_306)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_160),
.Y(n_245)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_129),
.B(n_133),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_141),
.B(n_173),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_257),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_147),
.Y(n_248)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_166),
.Y(n_249)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_160),
.Y(n_250)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_177),
.B1(n_168),
.B2(n_145),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_167),
.B(n_191),
.C(n_127),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_252),
.B(n_247),
.CI(n_202),
.CON(n_315),
.SN(n_315)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_253),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_134),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_254),
.B(n_255),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_136),
.B(n_132),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g256 ( 
.A1(n_150),
.A2(n_185),
.B1(n_153),
.B2(n_131),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_256),
.A2(n_263),
.B1(n_151),
.B2(n_165),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_185),
.B(n_140),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_258),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_259),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_189),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_143),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_123),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_261),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_137),
.A2(n_145),
.B1(n_168),
.B2(n_164),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_137),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_264),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_205),
.A2(n_131),
.B1(n_140),
.B2(n_123),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_265),
.A2(n_295),
.B1(n_297),
.B2(n_302),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_269),
.A2(n_308),
.B(n_219),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_164),
.B1(n_171),
.B2(n_146),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_278),
.A2(n_301),
.B1(n_305),
.B2(n_255),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_201),
.B(n_146),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_310),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_220),
.A2(n_151),
.B1(n_171),
.B2(n_165),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_233),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_208),
.A2(n_189),
.B1(n_196),
.B2(n_170),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_203),
.A2(n_170),
.B1(n_196),
.B2(n_199),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_304),
.A2(n_310),
.B1(n_316),
.B2(n_318),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_208),
.A2(n_213),
.B1(n_221),
.B2(n_256),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_231),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_242),
.A2(n_223),
.B1(n_201),
.B2(n_202),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_234),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_256),
.A2(n_262),
.B1(n_207),
.B2(n_255),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_256),
.A2(n_207),
.B1(n_233),
.B2(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_320),
.Y(n_374)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_322),
.B(n_328),
.Y(n_369)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_269),
.Y(n_324)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_324),
.Y(n_368)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_325),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_338),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_327),
.A2(n_340),
.B1(n_353),
.B2(n_285),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_244),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_211),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_330),
.B(n_332),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_331),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_306),
.B(n_216),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_268),
.B(n_252),
.C(n_215),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_350),
.C(n_270),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_222),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_335),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_282),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_317),
.Y(n_336)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_336),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_337),
.B(n_349),
.C(n_356),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_275),
.B(n_227),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_341),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_290),
.A2(n_229),
.B1(n_258),
.B2(n_260),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_249),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_342),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_268),
.B(n_254),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_345),
.Y(n_367)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_348),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_240),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_291),
.B(n_214),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_296),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_352),
.Y(n_381)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_286),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_279),
.A2(n_253),
.B1(n_248),
.B2(n_239),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_355),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_274),
.A2(n_302),
.B1(n_304),
.B2(n_318),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_307),
.B(n_236),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_298),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_358),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_230),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_307),
.A2(n_228),
.B(n_264),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_337),
.C(n_278),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_373),
.C(n_325),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_347),
.A2(n_300),
.B(n_309),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_370),
.A2(n_371),
.B(n_280),
.Y(n_413)
);

A2O1A1Ixp33_ASAP7_75t_SL g371 ( 
.A1(n_347),
.A2(n_309),
.B(n_279),
.C(n_297),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_333),
.C(n_358),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_362),
.Y(n_411)
);

AO22x1_ASAP7_75t_SL g378 ( 
.A1(n_324),
.A2(n_266),
.B1(n_307),
.B2(n_267),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_392),
.Y(n_397)
);

AO22x1_ASAP7_75t_L g379 ( 
.A1(n_341),
.A2(n_272),
.B1(n_266),
.B2(n_315),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_379),
.B(n_356),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_326),
.A2(n_272),
.B1(n_267),
.B2(n_270),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_382),
.A2(n_385),
.B1(n_393),
.B2(n_344),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_327),
.A2(n_309),
.B1(n_312),
.B2(n_311),
.Y(n_385)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_287),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_323),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_343),
.B(n_293),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_349),
.A2(n_313),
.B1(n_311),
.B2(n_245),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_337),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_402),
.C(n_415),
.Y(n_422)
);

A2O1A1O1Ixp25_ASAP7_75t_L g429 ( 
.A1(n_395),
.A2(n_417),
.B(n_397),
.C(n_406),
.D(n_407),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_381),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_398),
.Y(n_426)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_399),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_400),
.A2(n_401),
.B1(n_410),
.B2(n_365),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_386),
.A2(n_344),
.B1(n_335),
.B2(n_319),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_363),
.B(n_322),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_366),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_412),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_405),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_320),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_406),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_329),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_407),
.B(n_408),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_364),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_409),
.A2(n_419),
.B1(n_420),
.B2(n_380),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_411),
.A2(n_414),
.B(n_379),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_391),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_413),
.A2(n_371),
.B(n_376),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_375),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_370),
.A2(n_339),
.B1(n_351),
.B2(n_345),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_418),
.B1(n_390),
.B2(n_384),
.Y(n_425)
);

OA21x2_ASAP7_75t_SL g417 ( 
.A1(n_389),
.A2(n_354),
.B(n_352),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_386),
.A2(n_336),
.B1(n_321),
.B2(n_313),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_374),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_287),
.C(n_280),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_383),
.C(n_375),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_379),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_432),
.C(n_433),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_427),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_428),
.A2(n_430),
.B1(n_445),
.B2(n_414),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_429),
.A2(n_436),
.B(n_441),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_401),
.A2(n_388),
.B1(n_368),
.B2(n_360),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_361),
.C(n_378),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_360),
.B1(n_369),
.B2(n_387),
.Y(n_434)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_434),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_361),
.C(n_378),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_437),
.C(n_417),
.Y(n_461)
);

A2O1A1O1Ixp25_ASAP7_75t_L g436 ( 
.A1(n_395),
.A2(n_368),
.B(n_371),
.C(n_384),
.D(n_380),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_371),
.C(n_390),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_416),
.A2(n_371),
.B1(n_393),
.B2(n_376),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_372),
.B1(n_346),
.B2(n_276),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_400),
.A2(n_413),
.B1(n_397),
.B2(n_398),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_421),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_453),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_441),
.A2(n_403),
.B(n_411),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_447),
.A2(n_462),
.B(n_452),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_411),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_438),
.Y(n_451)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_404),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_443),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_455),
.Y(n_471)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_440),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_399),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_432),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_458),
.A2(n_426),
.B1(n_457),
.B2(n_448),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_420),
.B1(n_405),
.B2(n_419),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_460),
.A2(n_464),
.B1(n_445),
.B2(n_426),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_461),
.A2(n_437),
.B(n_429),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_423),
.A2(n_409),
.B(n_418),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_439),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_463),
.B(n_465),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_293),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_473),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_467),
.B(n_468),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_433),
.Y(n_468)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_480),
.C(n_449),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_424),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_439),
.C(n_430),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_477),
.Y(n_491)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_444),
.C(n_425),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_479),
.A2(n_314),
.B1(n_299),
.B2(n_288),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_442),
.C(n_372),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_481),
.A2(n_461),
.B1(n_449),
.B2(n_452),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_494),
.Y(n_503)
);

XOR2x1_ASAP7_75t_SL g483 ( 
.A(n_466),
.B(n_450),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_492),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_457),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_486),
.B(n_488),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_487),
.B(n_474),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_471),
.B(n_442),
.Y(n_488)
);

AOI21x1_ASAP7_75t_L g492 ( 
.A1(n_481),
.A2(n_450),
.B(n_447),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_462),
.C(n_464),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_472),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_491),
.B(n_476),
.C(n_477),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_498),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_490),
.B(n_475),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_500),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_480),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_502),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_467),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_489),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_495),
.B(n_496),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_483),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_505),
.A2(n_508),
.B(n_271),
.Y(n_518)
);

AOI322xp5_ASAP7_75t_L g507 ( 
.A1(n_499),
.A2(n_482),
.A3(n_485),
.B1(n_468),
.B2(n_473),
.C1(n_314),
.C2(n_303),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_511),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_503),
.B(n_485),
.C(n_299),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_210),
.B1(n_250),
.B2(n_198),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_512),
.B(n_288),
.Y(n_514)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_514),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_509),
.B(n_294),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_511),
.B(n_303),
.C(n_512),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_294),
.Y(n_516)
);

OAI21x1_ASAP7_75t_SL g519 ( 
.A1(n_516),
.A2(n_517),
.B(n_518),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_271),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_519),
.B(n_277),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_513),
.C(n_517),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_523),
.Y(n_524)
);

MAJx2_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_277),
.C(n_248),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_248),
.Y(n_526)
);


endmodule