module real_aes_8190_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g468 ( .A(n_1), .Y(n_468) );
INVx1_ASAP7_75t_L g252 ( .A(n_2), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_3), .A2(n_37), .B1(n_202), .B2(n_507), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_4), .B(n_445), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g213 ( .A1(n_5), .A2(n_135), .B(n_214), .Y(n_213) );
XNOR2xp5_ASAP7_75t_L g119 ( .A(n_6), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_6), .B(n_157), .Y(n_493) );
AND2x6_ASAP7_75t_L g140 ( .A(n_7), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_8), .A2(n_134), .B(n_142), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_9), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_9), .B(n_38), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_10), .B(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g219 ( .A(n_11), .Y(n_219) );
INVx1_ASAP7_75t_L g132 ( .A(n_12), .Y(n_132) );
INVx1_ASAP7_75t_L g462 ( .A(n_13), .Y(n_462) );
INVx1_ASAP7_75t_L g152 ( .A(n_14), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_15), .B(n_226), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_16), .B(n_158), .Y(n_495) );
AO32x2_ASAP7_75t_L g541 ( .A1(n_17), .A2(n_157), .A3(n_173), .B1(n_481), .B2(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_18), .B(n_202), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_19), .B(n_169), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_20), .B(n_158), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_21), .A2(n_49), .B1(n_202), .B2(n_507), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_22), .B(n_135), .Y(n_162) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_23), .A2(n_78), .B1(n_202), .B2(n_226), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_24), .B(n_202), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_25), .B(n_212), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_26), .A2(n_149), .B(n_151), .C(n_153), .Y(n_148) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_28), .B(n_128), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_29), .B(n_184), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_30), .A2(n_102), .B1(n_734), .B2(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_30), .Y(n_735) );
INVx1_ASAP7_75t_L g231 ( .A(n_31), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_32), .B(n_128), .Y(n_519) );
INVx2_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_34), .B(n_202), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_35), .B(n_128), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_36), .A2(n_140), .B(n_145), .C(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g114 ( .A(n_38), .Y(n_114) );
INVx1_ASAP7_75t_L g229 ( .A(n_39), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_40), .B(n_184), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_41), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_41), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_42), .B(n_202), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_43), .A2(n_88), .B1(n_154), .B2(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_44), .B(n_202), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_45), .B(n_202), .Y(n_463) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_46), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_47), .B(n_467), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_48), .B(n_135), .Y(n_203) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_50), .A2(n_60), .B1(n_202), .B2(n_226), .Y(n_499) );
OAI22xp5_ASAP7_75t_SL g430 ( .A1(n_51), .A2(n_431), .B1(n_434), .B2(n_435), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_51), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_52), .A2(n_145), .B1(n_226), .B2(n_228), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_53), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_54), .B(n_202), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_55), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_56), .B(n_202), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_57), .A2(n_217), .B(n_218), .C(n_220), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_58), .Y(n_188) );
INVx1_ASAP7_75t_L g215 ( .A(n_59), .Y(n_215) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_62), .A2(n_733), .B1(n_736), .B2(n_737), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_62), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_63), .B(n_202), .Y(n_469) );
INVx1_ASAP7_75t_L g131 ( .A(n_64), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_65), .A2(n_77), .B1(n_432), .B2(n_433), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_65), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
AO32x2_ASAP7_75t_L g504 ( .A1(n_67), .A2(n_157), .A3(n_194), .B1(n_481), .B2(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g479 ( .A(n_68), .Y(n_479) );
INVx1_ASAP7_75t_L g514 ( .A(n_69), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_SL g239 ( .A1(n_70), .A2(n_169), .B(n_220), .C(n_240), .Y(n_239) );
INVxp67_ASAP7_75t_L g241 ( .A(n_71), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_72), .B(n_226), .Y(n_515) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_74), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_75), .A2(n_105), .B1(n_115), .B2(n_747), .Y(n_104) );
INVx1_ASAP7_75t_L g179 ( .A(n_76), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_77), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_79), .A2(n_140), .B(n_145), .C(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_80), .B(n_507), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_81), .B(n_226), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_82), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_84), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_85), .B(n_226), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_86), .A2(n_140), .B(n_145), .C(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g440 ( .A(n_87), .B(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g450 ( .A(n_87), .B(n_442), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_89), .A2(n_103), .B1(n_226), .B2(n_227), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_90), .B(n_128), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_91), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_92), .A2(n_140), .B(n_145), .C(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_93), .Y(n_205) );
INVx1_ASAP7_75t_L g238 ( .A(n_94), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g143 ( .A(n_95), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_96), .B(n_166), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_97), .B(n_226), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_98), .B(n_157), .Y(n_156) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_99), .A2(n_449), .B1(n_728), .B2(n_729), .C1(n_738), .C2(n_741), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_101), .A2(n_135), .B(n_237), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_102), .Y(n_734) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g748 ( .A(n_106), .Y(n_748) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g442 ( .A(n_108), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g727 ( .A(n_109), .B(n_442), .Y(n_727) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_109), .B(n_441), .Y(n_743) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_118), .B(n_447), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g746 ( .A(n_117), .Y(n_746) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_437), .B(n_444), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_429), .B1(n_430), .B2(n_436), .Y(n_120) );
INVx2_ASAP7_75t_SL g436 ( .A(n_121), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_121), .A2(n_450), .B1(n_452), .B2(n_739), .Y(n_738) );
OR4x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_325), .C(n_384), .D(n_411), .Y(n_121) );
NAND3xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_267), .C(n_292), .Y(n_122) );
O2A1O1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_190), .B(n_210), .C(n_243), .Y(n_123) );
AOI211xp5_ASAP7_75t_SL g415 ( .A1(n_124), .A2(n_416), .B(n_418), .C(n_421), .Y(n_415) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_159), .Y(n_124) );
INVx1_ASAP7_75t_L g290 ( .A(n_125), .Y(n_290) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g265 ( .A(n_126), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g297 ( .A(n_126), .Y(n_297) );
AND2x2_ASAP7_75t_L g352 ( .A(n_126), .B(n_321), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_126), .B(n_208), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_126), .B(n_209), .Y(n_410) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g271 ( .A(n_127), .Y(n_271) );
AND2x2_ASAP7_75t_L g314 ( .A(n_127), .B(n_177), .Y(n_314) );
AND2x2_ASAP7_75t_L g332 ( .A(n_127), .B(n_209), .Y(n_332) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_133), .B(n_156), .Y(n_127) );
INVx1_ASAP7_75t_L g189 ( .A(n_128), .Y(n_189) );
INVx2_ASAP7_75t_L g194 ( .A(n_128), .Y(n_194) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_128), .A2(n_512), .B(n_519), .Y(n_511) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_128), .A2(n_521), .B(n_529), .Y(n_520) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_L g158 ( .A(n_129), .B(n_130), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
BUFx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_136), .B(n_140), .Y(n_180) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g467 ( .A(n_137), .Y(n_467) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
INVx1_ASAP7_75t_L g227 ( .A(n_138), .Y(n_227) );
INVx1_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx3_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
INVx4_ASAP7_75t_SL g155 ( .A(n_140), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_140), .A2(n_461), .B(n_465), .Y(n_460) );
BUFx3_ASAP7_75t_L g481 ( .A(n_140), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_140), .A2(n_487), .B(n_490), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_140), .A2(n_513), .B(n_516), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_140), .A2(n_522), .B(n_526), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_148), .C(n_155), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_144), .A2(n_155), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_144), .A2(n_155), .B(n_238), .C(n_239), .Y(n_237) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_146), .Y(n_202) );
INVx1_ASAP7_75t_L g507 ( .A(n_146), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_149), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g464 ( .A(n_149), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_149), .A2(n_517), .B(n_518), .Y(n_516) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g228 ( .A1(n_150), .A2(n_229), .B1(n_230), .B2(n_231), .Y(n_228) );
INVx2_ASAP7_75t_L g230 ( .A(n_150), .Y(n_230) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
OAI22xp33_ASAP7_75t_L g224 ( .A1(n_155), .A2(n_180), .B1(n_225), .B2(n_232), .Y(n_224) );
INVx4_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_157), .A2(n_236), .B(n_242), .Y(n_235) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_157), .A2(n_486), .B(n_493), .Y(n_485) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
INVx4_ASAP7_75t_L g264 ( .A(n_159), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g319 ( .A1(n_159), .A2(n_320), .B(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_L g400 ( .A(n_159), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_177), .Y(n_159) );
INVx1_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
AND2x2_ASAP7_75t_L g269 ( .A(n_160), .B(n_209), .Y(n_269) );
OR2x2_ASAP7_75t_L g298 ( .A(n_160), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g312 ( .A(n_160), .Y(n_312) );
INVx3_ASAP7_75t_L g321 ( .A(n_160), .Y(n_321) );
AND2x2_ASAP7_75t_L g331 ( .A(n_160), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g364 ( .A(n_160), .B(n_270), .Y(n_364) );
AND2x2_ASAP7_75t_L g388 ( .A(n_160), .B(n_344), .Y(n_388) );
OR2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_174), .Y(n_160) );
AOI21xp5_ASAP7_75t_SL g161 ( .A1(n_162), .A2(n_163), .B(n_172), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_170), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_166), .A2(n_252), .B(n_253), .C(n_254), .Y(n_251) );
INVx2_ASAP7_75t_L g470 ( .A(n_166), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_166), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_166), .A2(n_488), .B(n_489), .Y(n_487) );
O2A1O1Ixp5_ASAP7_75t_SL g513 ( .A1(n_166), .A2(n_220), .B(n_514), .C(n_515), .Y(n_513) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_167), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_167), .B(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g505 ( .A1(n_167), .A2(n_184), .B1(n_506), .B2(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g525 ( .A(n_169), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_170), .A2(n_183), .B(n_185), .Y(n_182) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_172), .A2(n_460), .B(n_471), .Y(n_459) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_172), .A2(n_474), .B(n_482), .Y(n_473) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_173), .A2(n_224), .B(n_233), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_173), .B(n_234), .Y(n_233) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_173), .A2(n_248), .B(n_255), .Y(n_247) );
NOR2xp33_ASAP7_75t_SL g174 ( .A(n_175), .B(n_176), .Y(n_174) );
INVx3_ASAP7_75t_L g212 ( .A(n_176), .Y(n_212) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_176), .B(n_481), .C(n_497), .Y(n_496) );
AO21x1_ASAP7_75t_L g575 ( .A1(n_176), .A2(n_497), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g209 ( .A(n_177), .Y(n_209) );
AND2x2_ASAP7_75t_L g424 ( .A(n_177), .B(n_266), .Y(n_424) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_186), .B(n_187), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g248 ( .A1(n_180), .A2(n_249), .B(n_250), .Y(n_248) );
INVx4_ASAP7_75t_L g200 ( .A(n_184), .Y(n_200) );
INVx2_ASAP7_75t_L g217 ( .A(n_184), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_184), .A2(n_470), .B1(n_498), .B2(n_499), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_184), .A2(n_470), .B1(n_543), .B2(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_189), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_189), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_206), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_192), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g344 ( .A(n_192), .B(n_332), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_192), .B(n_321), .Y(n_406) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g266 ( .A(n_193), .Y(n_266) );
AND2x2_ASAP7_75t_L g270 ( .A(n_193), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g311 ( .A(n_193), .B(n_312), .Y(n_311) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_204), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_203), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_201), .Y(n_197) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g220 ( .A(n_202), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_206), .B(n_307), .Y(n_329) );
INVx1_ASAP7_75t_L g368 ( .A(n_206), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_206), .B(n_295), .Y(n_412) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
AND2x2_ASAP7_75t_L g275 ( .A(n_207), .B(n_270), .Y(n_275) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_209), .B(n_266), .Y(n_299) );
INVx1_ASAP7_75t_L g378 ( .A(n_209), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g402 ( .A1(n_210), .A2(n_317), .A3(n_377), .B1(n_403), .B2(n_405), .C1(n_407), .C2(n_409), .Y(n_402) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_211), .B(n_222), .Y(n_210) );
AND2x2_ASAP7_75t_L g257 ( .A(n_211), .B(n_235), .Y(n_257) );
INVx1_ASAP7_75t_SL g260 ( .A(n_211), .Y(n_260) );
AND2x2_ASAP7_75t_L g262 ( .A(n_211), .B(n_223), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_211), .B(n_279), .Y(n_285) );
INVx2_ASAP7_75t_L g304 ( .A(n_211), .Y(n_304) );
AND2x2_ASAP7_75t_L g317 ( .A(n_211), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g355 ( .A(n_211), .B(n_279), .Y(n_355) );
BUFx2_ASAP7_75t_L g372 ( .A(n_211), .Y(n_372) );
AND2x2_ASAP7_75t_L g386 ( .A(n_211), .B(n_246), .Y(n_386) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_221), .Y(n_211) );
O2A1O1Ixp5_ASAP7_75t_L g478 ( .A1(n_217), .A2(n_466), .B(n_479), .C(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_217), .A2(n_527), .B(n_528), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_222), .B(n_274), .Y(n_301) );
AND2x2_ASAP7_75t_L g428 ( .A(n_222), .B(n_304), .Y(n_428) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_235), .Y(n_222) );
OR2x2_ASAP7_75t_L g273 ( .A(n_223), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
AND2x2_ASAP7_75t_L g324 ( .A(n_223), .B(n_247), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_223), .B(n_372), .Y(n_371) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_223), .Y(n_408) );
INVx2_ASAP7_75t_L g254 ( .A(n_226), .Y(n_254) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g259 ( .A(n_235), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g281 ( .A(n_235), .Y(n_281) );
BUFx2_ASAP7_75t_L g287 ( .A(n_235), .Y(n_287) );
AND2x2_ASAP7_75t_L g306 ( .A(n_235), .B(n_279), .Y(n_306) );
INVx3_ASAP7_75t_L g318 ( .A(n_235), .Y(n_318) );
OR2x2_ASAP7_75t_L g328 ( .A(n_235), .B(n_279), .Y(n_328) );
AOI31xp33_ASAP7_75t_SL g243 ( .A1(n_244), .A2(n_258), .A3(n_261), .B(n_263), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_257), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_245), .B(n_280), .Y(n_291) );
OR2x2_ASAP7_75t_L g315 ( .A(n_245), .B(n_285), .Y(n_315) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_246), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g336 ( .A(n_246), .B(n_328), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_246), .B(n_318), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_246), .B(n_354), .Y(n_353) );
NAND2x1_ASAP7_75t_L g381 ( .A(n_246), .B(n_317), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_246), .B(n_372), .Y(n_382) );
AND2x2_ASAP7_75t_L g394 ( .A(n_246), .B(n_279), .Y(n_394) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g274 ( .A(n_247), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_254), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g340 ( .A(n_257), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_257), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_259), .B(n_335), .Y(n_369) );
AND2x4_ASAP7_75t_L g280 ( .A(n_260), .B(n_281), .Y(n_280) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g359 ( .A(n_265), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_265), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g307 ( .A(n_266), .B(n_297), .Y(n_307) );
AND2x2_ASAP7_75t_L g401 ( .A(n_266), .B(n_271), .Y(n_401) );
INVx1_ASAP7_75t_L g426 ( .A(n_266), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .B1(n_275), .B2(n_276), .C(n_282), .Y(n_267) );
CKINVDCx14_ASAP7_75t_R g288 ( .A(n_268), .Y(n_288) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_269), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_272), .B(n_323), .Y(n_342) );
INVx3_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g391 ( .A(n_273), .B(n_287), .Y(n_391) );
AND2x2_ASAP7_75t_L g305 ( .A(n_274), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g335 ( .A(n_274), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_274), .B(n_318), .Y(n_363) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_274), .B(n_375), .C(n_406), .Y(n_405) );
AOI211xp5_ASAP7_75t_SL g338 ( .A1(n_275), .A2(n_339), .B(n_341), .C(n_349), .Y(n_338) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g327 ( .A1(n_277), .A2(n_328), .B1(n_329), .B2(n_330), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_278), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_278), .B(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g420 ( .A(n_280), .B(n_394), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_288), .B1(n_289), .B2(n_291), .Y(n_282) );
NOR2xp33_ASAP7_75t_SL g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_286), .B(n_335), .Y(n_366) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_289), .A2(n_381), .B1(n_412), .B2(n_419), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_300), .B1(n_302), .B2(n_307), .C(n_308), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_298), .A2(n_309), .B1(n_315), .B2(n_316), .C(n_319), .Y(n_308) );
INVx1_ASAP7_75t_L g351 ( .A(n_299), .Y(n_351) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_SL g323 ( .A(n_304), .Y(n_323) );
OR2x2_ASAP7_75t_L g396 ( .A(n_304), .B(n_328), .Y(n_396) );
AND2x2_ASAP7_75t_L g398 ( .A(n_304), .B(n_306), .Y(n_398) );
INVx1_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
AOI21xp33_ASAP7_75t_SL g367 ( .A1(n_310), .A2(n_368), .B(n_369), .Y(n_367) );
OR2x2_ASAP7_75t_L g374 ( .A(n_310), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g348 ( .A(n_311), .B(n_332), .Y(n_348) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp33_ASAP7_75t_SL g365 ( .A(n_316), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_317), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_318), .B(n_354), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_321), .A2(n_334), .B(n_336), .C(n_337), .Y(n_333) );
NAND2x1_ASAP7_75t_SL g358 ( .A(n_321), .B(n_359), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_322), .A2(n_371), .B1(n_373), .B2(n_376), .Y(n_370) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_324), .B(n_414), .Y(n_413) );
NAND5xp2_ASAP7_75t_L g325 ( .A(n_326), .B(n_338), .C(n_356), .D(n_370), .E(n_379), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_327), .B(n_333), .Y(n_326) );
INVx1_ASAP7_75t_L g383 ( .A(n_329), .Y(n_383) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_331), .A2(n_350), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_332), .B(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_335), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_335), .B(n_401), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_345), .B2(n_347), .Y(n_341) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x2_ASAP7_75t_L g423 ( .A(n_352), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B1(n_364), .B2(n_365), .C(n_367), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g407 ( .A(n_362), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g414 ( .A(n_372), .Y(n_414) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI21xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_382), .B(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_387), .B(n_389), .C(n_402), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g411 ( .A1(n_387), .A2(n_412), .B(n_413), .C(n_415), .Y(n_411) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_391), .B(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .B(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
CKINVDCx14_ASAP7_75t_R g435 ( .A(n_431), .Y(n_435) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_436), .A2(n_450), .B1(n_451), .B2(n_727), .Y(n_449) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_440), .Y(n_446) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_444), .B(n_448), .C(n_744), .Y(n_447) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR5x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_618), .C(n_676), .D(n_712), .E(n_719), .Y(n_454) );
NAND3xp33_ASAP7_75t_SL g455 ( .A(n_456), .B(n_564), .C(n_588), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_500), .B1(n_530), .B2(n_535), .C(n_545), .Y(n_456) );
OAI21xp5_ASAP7_75t_SL g698 ( .A1(n_457), .A2(n_699), .B(n_701), .Y(n_698) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_483), .Y(n_457) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_458), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_472), .Y(n_458) );
INVx2_ASAP7_75t_L g534 ( .A(n_459), .Y(n_534) );
AND2x2_ASAP7_75t_L g547 ( .A(n_459), .B(n_485), .Y(n_547) );
AND2x2_ASAP7_75t_L g601 ( .A(n_459), .B(n_484), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_459), .B(n_473), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_468), .B(n_469), .C(n_470), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_470), .A2(n_491), .B(n_492), .Y(n_490) );
AND2x2_ASAP7_75t_L g634 ( .A(n_472), .B(n_575), .Y(n_634) );
AND2x2_ASAP7_75t_L g667 ( .A(n_472), .B(n_485), .Y(n_667) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g574 ( .A(n_473), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g587 ( .A(n_473), .B(n_485), .Y(n_587) );
AND2x2_ASAP7_75t_L g594 ( .A(n_473), .B(n_575), .Y(n_594) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_473), .Y(n_603) );
AND2x2_ASAP7_75t_L g610 ( .A(n_473), .B(n_484), .Y(n_610) );
INVx1_ASAP7_75t_L g641 ( .A(n_473), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_478), .B(n_481), .Y(n_474) );
INVx1_ASAP7_75t_L g617 ( .A(n_483), .Y(n_617) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_494), .Y(n_483) );
INVx2_ASAP7_75t_L g573 ( .A(n_484), .Y(n_573) );
AND2x2_ASAP7_75t_L g595 ( .A(n_484), .B(n_534), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_484), .B(n_641), .Y(n_646) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_485), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g718 ( .A(n_485), .B(n_682), .Y(n_718) );
INVx2_ASAP7_75t_L g532 ( .A(n_494), .Y(n_532) );
INVx3_ASAP7_75t_L g633 ( .A(n_494), .Y(n_633) );
OR2x2_ASAP7_75t_L g663 ( .A(n_494), .B(n_664), .Y(n_663) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_494), .B(n_573), .Y(n_689) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g576 ( .A(n_495), .Y(n_576) );
AOI33xp33_ASAP7_75t_L g709 ( .A1(n_500), .A2(n_547), .A3(n_561), .B1(n_633), .B2(n_710), .B3(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_509), .Y(n_501) );
OR2x2_ASAP7_75t_L g562 ( .A(n_502), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_502), .B(n_559), .Y(n_621) );
OR2x2_ASAP7_75t_L g674 ( .A(n_502), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g600 ( .A(n_503), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g625 ( .A(n_503), .B(n_509), .Y(n_625) );
AND2x2_ASAP7_75t_L g692 ( .A(n_503), .B(n_537), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_503), .A2(n_592), .B(n_718), .Y(n_717) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g539 ( .A(n_504), .Y(n_539) );
INVx1_ASAP7_75t_L g552 ( .A(n_504), .Y(n_552) );
AND2x2_ASAP7_75t_L g571 ( .A(n_504), .B(n_541), .Y(n_571) );
AND2x2_ASAP7_75t_L g620 ( .A(n_504), .B(n_540), .Y(n_620) );
INVx2_ASAP7_75t_SL g662 ( .A(n_509), .Y(n_662) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
INVx2_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
INVx1_ASAP7_75t_L g713 ( .A(n_510), .Y(n_713) );
AND2x2_ASAP7_75t_L g726 ( .A(n_510), .B(n_607), .Y(n_726) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g553 ( .A(n_511), .Y(n_553) );
OR2x2_ASAP7_75t_L g559 ( .A(n_511), .B(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_511), .Y(n_570) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_520), .Y(n_537) );
AND2x2_ASAP7_75t_L g554 ( .A(n_520), .B(n_540), .Y(n_554) );
INVx1_ASAP7_75t_L g560 ( .A(n_520), .Y(n_560) );
INVx1_ASAP7_75t_L g567 ( .A(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g592 ( .A(n_520), .B(n_541), .Y(n_592) );
INVx2_ASAP7_75t_L g608 ( .A(n_520), .Y(n_608) );
AND2x2_ASAP7_75t_L g701 ( .A(n_520), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_520), .B(n_582), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_525), .Y(n_522) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
INVx1_ASAP7_75t_L g585 ( .A(n_532), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_532), .B(n_616), .Y(n_682) );
INVx1_ASAP7_75t_SL g642 ( .A(n_533), .Y(n_642) );
INVx2_ASAP7_75t_L g563 ( .A(n_534), .Y(n_563) );
AND2x2_ASAP7_75t_L g632 ( .A(n_534), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g648 ( .A(n_534), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
INVx1_ASAP7_75t_L g710 ( .A(n_536), .Y(n_710) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g565 ( .A(n_538), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g668 ( .A(n_538), .B(n_658), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_538), .A2(n_679), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AND2x2_ASAP7_75t_L g581 ( .A(n_539), .B(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
INVx1_ASAP7_75t_L g630 ( .A(n_539), .Y(n_630) );
OR2x2_ASAP7_75t_L g694 ( .A(n_540), .B(n_553), .Y(n_694) );
NOR2xp67_ASAP7_75t_L g702 ( .A(n_540), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g607 ( .A(n_541), .B(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g614 ( .A(n_541), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_548), .B1(n_555), .B2(n_557), .Y(n_545) );
OR2x2_ASAP7_75t_L g624 ( .A(n_546), .B(n_574), .Y(n_624) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_547), .A2(n_666), .B1(n_668), .B2(n_669), .C1(n_670), .C2(n_673), .Y(n_665) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g612 ( .A(n_551), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_SL g566 ( .A(n_553), .B(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_553), .Y(n_637) );
AND2x2_ASAP7_75t_L g685 ( .A(n_553), .B(n_554), .Y(n_685) );
INVx1_ASAP7_75t_L g703 ( .A(n_553), .Y(n_703) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g669 ( .A(n_556), .B(n_595), .Y(n_669) );
AND2x2_ASAP7_75t_L g711 ( .A(n_556), .B(n_587), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_558), .B(n_606), .Y(n_693) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_559), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g586 ( .A(n_563), .B(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g654 ( .A(n_563), .Y(n_654) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .B(n_572), .C(n_577), .Y(n_564) );
INVxp67_ASAP7_75t_L g578 ( .A(n_565), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_566), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_566), .B(n_613), .Y(n_708) );
BUFx3_ASAP7_75t_L g672 ( .A(n_567), .Y(n_672) );
INVx1_ASAP7_75t_L g579 ( .A(n_568), .Y(n_579) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g598 ( .A(n_570), .B(n_592), .Y(n_598) );
INVx1_ASAP7_75t_SL g638 ( .A(n_571), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g628 ( .A(n_573), .Y(n_628) );
AND2x2_ASAP7_75t_L g651 ( .A(n_573), .B(n_634), .Y(n_651) );
INVx1_ASAP7_75t_SL g622 ( .A(n_574), .Y(n_622) );
INVx1_ASAP7_75t_L g649 ( .A(n_575), .Y(n_649) );
AOI31xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .A3(n_580), .B(n_583), .Y(n_577) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g670 ( .A(n_581), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g644 ( .A(n_582), .Y(n_644) );
BUFx2_ASAP7_75t_L g658 ( .A(n_582), .Y(n_658) );
AND2x2_ASAP7_75t_L g686 ( .A(n_582), .B(n_607), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g659 ( .A(n_586), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_587), .B(n_654), .Y(n_700) );
AND2x2_ASAP7_75t_L g707 ( .A(n_587), .B(n_633), .Y(n_707) );
AOI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_593), .B(n_596), .C(n_611), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_593), .A2(n_620), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_619) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g627 ( .A(n_594), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g664 ( .A(n_595), .Y(n_664) );
OAI32xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .A3(n_602), .B1(n_604), .B2(n_609), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_598), .A2(n_651), .B(n_652), .C(n_655), .Y(n_650) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_606), .A2(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g675 ( .A(n_607), .Y(n_675) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_612), .B(n_615), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_613), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g661 ( .A(n_613), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g678 ( .A(n_615), .Y(n_678) );
OR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND4xp25_ASAP7_75t_SL g618 ( .A(n_619), .B(n_631), .C(n_650), .D(n_665), .Y(n_618) );
AND2x2_ASAP7_75t_L g657 ( .A(n_620), .B(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g679 ( .A(n_620), .B(n_672), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_622), .B(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_626), .B2(n_629), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_624), .A2(n_675), .B1(n_706), .B2(n_708), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_624), .A2(n_713), .B(n_714), .C(n_717), .Y(n_712) );
INVx2_ASAP7_75t_L g683 ( .A(n_625), .Y(n_683) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI222xp33_ASAP7_75t_L g677 ( .A1(n_627), .A2(n_661), .B1(n_678), .B2(n_679), .C1(n_680), .C2(n_683), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B(n_635), .C(n_639), .Y(n_631) );
INVx1_ASAP7_75t_L g697 ( .A(n_632), .Y(n_697) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_636), .A2(n_640), .B1(n_643), .B2(n_645), .Y(n_639) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g666 ( .A(n_648), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g724 ( .A(n_651), .Y(n_724) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B1(n_660), .B2(n_663), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_658), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g715 ( .A(n_663), .Y(n_715) );
INVx1_ASAP7_75t_L g696 ( .A(n_667), .Y(n_696) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_669), .Y(n_723) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND5xp2_ASAP7_75t_L g676 ( .A(n_677), .B(n_684), .C(n_698), .D(n_704), .E(n_709), .Y(n_676) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B(n_687), .C(n_690), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI31xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .A3(n_694), .B(n_695), .Y(n_690) );
INVx1_ASAP7_75t_L g716 ( .A(n_692), .Y(n_716) );
OR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI222xp33_ASAP7_75t_L g719 ( .A1(n_706), .A2(n_708), .B1(n_720), .B2(n_723), .C1(n_724), .C2(n_725), .Y(n_719) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g740 ( .A(n_727), .Y(n_740) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g736 ( .A(n_733), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
endmodule