module fake_netlist_5_2437_n_1290 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1290);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1290;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1286;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_12),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_33),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_82),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_17),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_8),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_98),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_90),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_26),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_69),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_141),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_55),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_174),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_16),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_60),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_187),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_28),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_23),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_176),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_139),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_162),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_115),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_118),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_163),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_38),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_2),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_10),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_5),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_46),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_6),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_47),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_42),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_6),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_56),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_92),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_52),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_86),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_181),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_32),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_27),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_100),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_29),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_146),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_49),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_105),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_122),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_33),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_38),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_34),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_23),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_67),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_119),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_160),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_126),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_167),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_85),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_68),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_95),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_24),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_63),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_102),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_188),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_75),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_103),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_70),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_145),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_148),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_191),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_19),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_21),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_177),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_136),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_170),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_183),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_50),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_42),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_182),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_88),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_171),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_110),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_114),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_4),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_64),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_150),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_59),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_127),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_78),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_149),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_157),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_72),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_65),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_158),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_41),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_179),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_44),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_133),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_1),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_113),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_125),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_8),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_186),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_45),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_45),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_41),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_14),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_28),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_87),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_200),
.B(n_0),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_213),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_236),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_196),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_264),
.B(n_0),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_236),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

BUFx6f_ASAP7_75t_SL g334 ( 
.A(n_247),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_206),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_216),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_201),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_210),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_203),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_1),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_242),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_210),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_264),
.B(n_3),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_3),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_316),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_238),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_249),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_214),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_215),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_238),
.B(n_4),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_221),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_319),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_223),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_216),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_275),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_228),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_292),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_275),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_249),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_206),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_288),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_199),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_283),
.B(n_5),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_300),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_197),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_198),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_202),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_205),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_280),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_231),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_280),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_204),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_247),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_284),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_233),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_284),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_241),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_211),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_244),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_217),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_245),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_265),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_253),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_268),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_218),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_222),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_219),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_289),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_292),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_207),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_227),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_269),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_220),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_229),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_227),
.B(n_7),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_289),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_232),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_313),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_271),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_313),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_240),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_274),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_246),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_292),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_281),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_225),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_209),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_226),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_336),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_328),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_334),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_389),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_339),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_389),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_338),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_259),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_398),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_353),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_354),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_337),
.B(n_279),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_323),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_362),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_325),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_326),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_356),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_345),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_368),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_393),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_407),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_331),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_358),
.B(n_248),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_332),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_347),
.A2(n_411),
.B(n_396),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_361),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_377),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_335),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_382),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_333),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_384),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_352),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_352),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_386),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_341),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_342),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_359),
.B(n_307),
.Y(n_463)
);

BUFx10_ASAP7_75t_L g464 ( 
.A(n_334),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_346),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_360),
.B(n_307),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_388),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_372),
.B(n_257),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_390),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_364),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_R g472 ( 
.A(n_391),
.B(n_286),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_349),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_363),
.B(n_230),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_350),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_399),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_357),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_406),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_409),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_R g484 ( 
.A(n_412),
.B(n_287),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_379),
.B(n_266),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_385),
.B(n_267),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_413),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_443),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_451),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_418),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_322),
.C(n_329),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_451),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_477),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_433),
.B(n_351),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_433),
.B(n_392),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_461),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

BUFx10_ASAP7_75t_L g504 ( 
.A(n_428),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_446),
.B(n_397),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_461),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_431),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_461),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_422),
.B(n_414),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_487),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_473),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_473),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_421),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_473),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_468),
.B(n_394),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_470),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_468),
.A2(n_355),
.B1(n_348),
.B2(n_410),
.Y(n_520)
);

INVx4_ASAP7_75t_SL g521 ( 
.A(n_420),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_452),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_423),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_470),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_424),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_460),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_468),
.B(n_400),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_463),
.B(n_343),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_422),
.B(n_365),
.Y(n_530)
);

BUFx6f_ASAP7_75t_SL g531 ( 
.A(n_464),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_473),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_470),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_463),
.B(n_466),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_429),
.B(n_324),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_470),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_468),
.B(n_265),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_424),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_483),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_477),
.A2(n_432),
.B1(n_449),
.B2(n_439),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_472),
.B(n_415),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_486),
.B(n_265),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_486),
.B(n_401),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_474),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_486),
.A2(n_404),
.B1(n_408),
.B2(n_369),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_474),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_423),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_416),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_417),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_486),
.B(n_366),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_484),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_417),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_466),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_489),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_537),
.A2(n_453),
.B1(n_455),
.B2(n_450),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_493),
.A2(n_482),
.B1(n_481),
.B2(n_479),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_559),
.A2(n_520),
.B1(n_547),
.B2(n_539),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_559),
.B(n_458),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_489),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_490),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_559),
.A2(n_448),
.B1(n_297),
.B2(n_315),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_SL g569 ( 
.A(n_523),
.B(n_376),
.C(n_364),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_540),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_496),
.A2(n_467),
.B1(n_469),
.B2(n_413),
.Y(n_571)
);

OAI22x1_ASAP7_75t_SL g572 ( 
.A1(n_512),
.A2(n_330),
.B1(n_327),
.B2(n_403),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_491),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_542),
.Y(n_575)
);

NAND3xp33_ASAP7_75t_SL g576 ( 
.A(n_523),
.B(n_378),
.C(n_376),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_549),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_497),
.B(n_448),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_513),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_476),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_535),
.B(n_441),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_496),
.B(n_464),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_517),
.B(n_419),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_528),
.B(n_548),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_549),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_490),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_527),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_513),
.B(n_464),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_500),
.B(n_419),
.Y(n_589)
);

AND2x6_ASAP7_75t_SL g590 ( 
.A(n_506),
.B(n_327),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_488),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_556),
.A2(n_518),
.B(n_502),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_529),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_529),
.B(n_442),
.Y(n_594)
);

BUFx6f_ASAP7_75t_SL g595 ( 
.A(n_492),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_514),
.B(n_426),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_514),
.B(n_426),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_529),
.B(n_367),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_557),
.B(n_415),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_557),
.B(n_344),
.Y(n_600)
);

OAI221xp5_ASAP7_75t_L g601 ( 
.A1(n_550),
.A2(n_402),
.B1(n_478),
.B2(n_475),
.C(n_465),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_488),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_502),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_516),
.B(n_532),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_544),
.B(n_344),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_516),
.B(n_270),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_546),
.B(n_378),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_539),
.A2(n_277),
.B1(n_305),
.B2(n_294),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_492),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_529),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_529),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_551),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_494),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_532),
.B(n_464),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_553),
.B(n_276),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_551),
.B(n_292),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_494),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_553),
.B(n_554),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_501),
.B(n_292),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_554),
.B(n_278),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_555),
.B(n_435),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_539),
.B(n_435),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_502),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_530),
.B(n_381),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_515),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_539),
.B(n_437),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_539),
.A2(n_295),
.B1(n_224),
.B2(n_293),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_511),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_515),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_437),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_504),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_539),
.B(n_438),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_547),
.B(n_438),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_547),
.B(n_445),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_519),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_558),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_558),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_547),
.B(n_445),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_547),
.B(n_495),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_547),
.B(n_447),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_495),
.B(n_370),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_547),
.B(n_447),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_498),
.B(n_371),
.C(n_454),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_498),
.B(n_454),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_499),
.B(n_459),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_524),
.A2(n_306),
.B1(n_321),
.B2(n_312),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_501),
.B(n_292),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_499),
.B(n_459),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_524),
.B(n_503),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_503),
.A2(n_480),
.B(n_478),
.C(n_475),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_531),
.B(n_381),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_491),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_510),
.B(n_462),
.Y(n_656)
);

NAND2x1_ASAP7_75t_L g657 ( 
.A(n_518),
.B(n_427),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_510),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_504),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_578),
.A2(n_507),
.B(n_533),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_581),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_603),
.A2(n_534),
.B(n_518),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_584),
.B(n_534),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_653),
.A2(n_480),
.B(n_462),
.C(n_465),
.Y(n_664)
);

AO21x1_ASAP7_75t_L g665 ( 
.A1(n_619),
.A2(n_538),
.B(n_534),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_581),
.B(n_504),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_563),
.B(n_508),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_653),
.A2(n_507),
.B(n_545),
.C(n_552),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_603),
.A2(n_538),
.B(n_505),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_568),
.A2(n_536),
.B(n_533),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_593),
.B(n_508),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_640),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_564),
.B(n_538),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_570),
.B(n_509),
.Y(n_675)
);

AOI21x1_ASAP7_75t_L g676 ( 
.A1(n_657),
.A2(n_541),
.B(n_536),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_603),
.A2(n_505),
.B(n_491),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_579),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_604),
.A2(n_541),
.B(n_545),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_658),
.Y(n_680)
);

O2A1O1Ixp5_ASAP7_75t_L g681 ( 
.A1(n_606),
.A2(n_552),
.B(n_543),
.C(n_509),
.Y(n_681)
);

O2A1O1Ixp5_ASAP7_75t_L g682 ( 
.A1(n_616),
.A2(n_543),
.B(n_509),
.C(n_526),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_592),
.A2(n_543),
.B(n_526),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_574),
.A2(n_282),
.B(n_234),
.C(n_235),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_655),
.Y(n_685)
);

OAI321xp33_ASAP7_75t_L g686 ( 
.A1(n_601),
.A2(n_434),
.A3(n_430),
.B1(n_427),
.B2(n_334),
.C(n_247),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_655),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_624),
.A2(n_505),
.B(n_491),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_640),
.Y(n_689)
);

AOI221xp5_ASAP7_75t_L g690 ( 
.A1(n_605),
.A2(n_256),
.B1(n_296),
.B2(n_237),
.C(n_239),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_575),
.B(n_526),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_624),
.A2(n_505),
.B(n_491),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_589),
.B(n_525),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_609),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_560),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_591),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_621),
.B(n_525),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_593),
.A2(n_383),
.B1(n_395),
.B2(n_403),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_610),
.A2(n_261),
.B(n_314),
.C(n_243),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_580),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_624),
.A2(n_505),
.B(n_522),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_655),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_580),
.B(n_525),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_652),
.A2(n_522),
.B(n_434),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_560),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_618),
.A2(n_430),
.B(n_383),
.C(n_395),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_591),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_573),
.A2(n_522),
.B(n_298),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_583),
.A2(n_522),
.B(n_308),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g710 ( 
.A1(n_655),
.A2(n_522),
.B(n_310),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_587),
.B(n_508),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_655),
.A2(n_522),
.B(n_304),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_577),
.B(n_585),
.Y(n_713)
);

A2O1A1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_610),
.A2(n_317),
.B(n_251),
.C(n_254),
.Y(n_714)
);

AOI221xp5_ASAP7_75t_L g715 ( 
.A1(n_607),
.A2(n_262),
.B1(n_309),
.B2(n_405),
.C(n_330),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_602),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_571),
.B(n_405),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_657),
.A2(n_302),
.B(n_521),
.Y(n_718)
);

OAI21xp33_ASAP7_75t_L g719 ( 
.A1(n_561),
.A2(n_303),
.B(n_212),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_615),
.A2(n_425),
.B(n_440),
.C(n_444),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_612),
.B(n_525),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_SL g722 ( 
.A1(n_619),
.A2(n_258),
.B(n_273),
.C(n_292),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_644),
.B(n_208),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_594),
.B(n_456),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_642),
.A2(n_299),
.B(n_212),
.Y(n_725)
);

NOR2xp67_ASAP7_75t_L g726 ( 
.A(n_562),
.B(n_208),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_566),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_630),
.B(n_531),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_644),
.B(n_255),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_622),
.B(n_656),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_596),
.A2(n_521),
.B(n_303),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_647),
.B(n_255),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_611),
.A2(n_531),
.B1(n_301),
.B2(n_299),
.Y(n_733)
);

AND2x2_ASAP7_75t_SL g734 ( 
.A(n_598),
.B(n_258),
.Y(n_734)
);

OAI21xp33_ASAP7_75t_L g735 ( 
.A1(n_599),
.A2(n_301),
.B(n_457),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_611),
.A2(n_471),
.B1(n_258),
.B2(n_273),
.Y(n_736)
);

AND2x6_ASAP7_75t_SL g737 ( 
.A(n_654),
.B(n_273),
.Y(n_737)
);

AO22x1_ASAP7_75t_L g738 ( 
.A1(n_625),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_566),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_597),
.A2(n_521),
.B(n_89),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_648),
.A2(n_521),
.B(n_91),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_565),
.B(n_11),
.Y(n_742)
);

AO22x1_ASAP7_75t_L g743 ( 
.A1(n_594),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_567),
.A2(n_93),
.B(n_192),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_651),
.A2(n_84),
.B(n_190),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_567),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_586),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_626),
.A2(n_83),
.B(n_178),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_609),
.B(n_13),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_569),
.B(n_576),
.C(n_600),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_598),
.B(n_602),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_586),
.A2(n_81),
.B(n_175),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_626),
.A2(n_195),
.B(n_80),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_613),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_613),
.B(n_14),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_650),
.A2(n_94),
.B(n_172),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_739),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_700),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_730),
.B(n_565),
.Y(n_759)
);

NAND2x1p5_ASAP7_75t_L g760 ( 
.A(n_685),
.B(n_627),
.Y(n_760)
);

OAI21x1_ASAP7_75t_L g761 ( 
.A1(n_676),
.A2(n_617),
.B(n_638),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_702),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_667),
.A2(n_751),
.B1(n_663),
.B2(n_678),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_683),
.A2(n_668),
.B(n_681),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_702),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_660),
.A2(n_616),
.B(n_650),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_693),
.A2(n_617),
.B(n_614),
.Y(n_767)
);

AOI21xp33_ASAP7_75t_L g768 ( 
.A1(n_666),
.A2(n_659),
.B(n_627),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_665),
.A2(n_707),
.B(n_696),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_670),
.A2(n_588),
.B(n_614),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_681),
.A2(n_638),
.B(n_631),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_700),
.B(n_590),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_682),
.A2(n_631),
.B(n_636),
.Y(n_773)
);

BUFx12f_ASAP7_75t_L g774 ( 
.A(n_737),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_682),
.A2(n_636),
.B(n_639),
.Y(n_775)
);

INVx4_ASAP7_75t_L g776 ( 
.A(n_702),
.Y(n_776)
);

OAI21x1_ASAP7_75t_SL g777 ( 
.A1(n_744),
.A2(n_752),
.B(n_756),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_667),
.A2(n_588),
.B1(n_659),
.B2(n_633),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_677),
.A2(n_620),
.B(n_634),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_703),
.B(n_646),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_715),
.B(n_649),
.C(n_582),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_680),
.B(n_673),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_661),
.B(n_582),
.Y(n_783)
);

OA21x2_ASAP7_75t_L g784 ( 
.A1(n_679),
.A2(n_645),
.B(n_643),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_739),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_694),
.B(n_671),
.Y(n_786)
);

OA21x2_ASAP7_75t_L g787 ( 
.A1(n_748),
.A2(n_641),
.B(n_637),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_713),
.B(n_633),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_723),
.B(n_729),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_666),
.B(n_623),
.Y(n_790)
);

OAI21x1_ASAP7_75t_L g791 ( 
.A1(n_688),
.A2(n_635),
.B(n_632),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_716),
.A2(n_754),
.B1(n_685),
.B2(n_674),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_742),
.A2(n_628),
.B(n_629),
.C(n_608),
.Y(n_793)
);

OAI22x1_ASAP7_75t_L g794 ( 
.A1(n_742),
.A2(n_572),
.B1(n_595),
.B2(n_17),
.Y(n_794)
);

OAI21x1_ASAP7_75t_L g795 ( 
.A1(n_692),
.A2(n_96),
.B(n_173),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_734),
.A2(n_595),
.B1(n_16),
.B2(n_18),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_669),
.A2(n_97),
.B(n_168),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_734),
.A2(n_595),
.B1(n_77),
.B2(n_101),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_716),
.Y(n_799)
);

A2O1A1Ixp33_ASAP7_75t_L g800 ( 
.A1(n_706),
.A2(n_15),
.B(n_19),
.C(n_20),
.Y(n_800)
);

OAI21x1_ASAP7_75t_L g801 ( 
.A1(n_662),
.A2(n_76),
.B(n_164),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_698),
.B(n_15),
.Y(n_802)
);

OAI21x1_ASAP7_75t_L g803 ( 
.A1(n_701),
.A2(n_74),
.B(n_159),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_702),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_685),
.A2(n_73),
.B(n_156),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_754),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_732),
.B(n_20),
.Y(n_807)
);

O2A1O1Ixp5_ASAP7_75t_L g808 ( 
.A1(n_725),
.A2(n_104),
.B(n_155),
.C(n_154),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_672),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_704),
.A2(n_66),
.B(n_153),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_685),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_675),
.A2(n_62),
.B(n_152),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_753),
.A2(n_61),
.B(n_151),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_691),
.A2(n_58),
.B(n_144),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_711),
.B(n_21),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_697),
.A2(n_721),
.B(n_747),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_689),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_684),
.B(n_22),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_684),
.B(n_22),
.Y(n_819)
);

AOI21x1_ASAP7_75t_L g820 ( 
.A1(n_709),
.A2(n_71),
.B(n_143),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_717),
.B(n_57),
.Y(n_821)
);

AO31x2_ASAP7_75t_L g822 ( 
.A1(n_699),
.A2(n_24),
.A3(n_25),
.B(n_26),
.Y(n_822)
);

BUFx12f_ASAP7_75t_L g823 ( 
.A(n_774),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_786),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_759),
.B(n_695),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_811),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_811),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_789),
.B(n_735),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_SL g829 ( 
.A(n_821),
.B(n_724),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_757),
.B(n_705),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_757),
.B(n_727),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_785),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_782),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_786),
.B(n_694),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_788),
.B(n_719),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_758),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_765),
.Y(n_837)
);

NAND2x1p5_ASAP7_75t_L g838 ( 
.A(n_765),
.B(n_687),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_758),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_777),
.A2(n_671),
.B(n_741),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_800),
.A2(n_750),
.B(n_736),
.C(n_720),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_785),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_790),
.B(n_750),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_807),
.B(n_726),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_815),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_772),
.B(n_728),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_809),
.B(n_746),
.Y(n_847)
);

BUFx10_ASAP7_75t_L g848 ( 
.A(n_772),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_770),
.A2(n_740),
.B(n_731),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_SL g850 ( 
.A(n_774),
.B(n_749),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_802),
.Y(n_851)
);

AND2x4_ASAP7_75t_SL g852 ( 
.A(n_776),
.B(n_687),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_817),
.B(n_747),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_776),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_799),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_760),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_806),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_783),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_768),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_760),
.B(n_743),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_780),
.B(n_728),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_781),
.B(n_733),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_762),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_763),
.B(n_699),
.Y(n_864)
);

CKINVDCx11_ASAP7_75t_R g865 ( 
.A(n_778),
.Y(n_865)
);

BUFx4_ASAP7_75t_SL g866 ( 
.A(n_794),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_798),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_790),
.B(n_714),
.Y(n_869)
);

INVx3_ASAP7_75t_SL g870 ( 
.A(n_804),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_804),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_818),
.B(n_755),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_796),
.B(n_714),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_SL g874 ( 
.A(n_800),
.B(n_745),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_797),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_771),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_796),
.B(n_690),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_770),
.B(n_664),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_L g879 ( 
.A(n_819),
.B(n_686),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_832),
.Y(n_880)
);

OA21x2_ASAP7_75t_L g881 ( 
.A1(n_849),
.A2(n_764),
.B(n_808),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_836),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_832),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_868),
.A2(n_829),
.B1(n_877),
.B2(n_859),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_842),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_840),
.A2(n_769),
.B(n_767),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_862),
.A2(n_812),
.B1(n_814),
.B2(n_767),
.Y(n_887)
);

NAND2x1p5_ASAP7_75t_L g888 ( 
.A(n_843),
.B(n_801),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_878),
.A2(n_820),
.B(n_816),
.Y(n_889)
);

OA21x2_ASAP7_75t_L g890 ( 
.A1(n_876),
.A2(n_808),
.B(n_761),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_826),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_830),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_876),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_826),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_825),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_836),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_834),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_868),
.A2(n_814),
.B1(n_792),
.B2(n_784),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_825),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_839),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_874),
.A2(n_766),
.B(n_793),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_864),
.A2(n_816),
.B(n_766),
.Y(n_902)
);

INVx8_ASAP7_75t_L g903 ( 
.A(n_826),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_859),
.A2(n_793),
.B1(n_784),
.B2(n_805),
.Y(n_904)
);

AOI21x1_ASAP7_75t_L g905 ( 
.A1(n_869),
.A2(n_779),
.B(n_787),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_830),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_843),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_853),
.B(n_822),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_831),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_831),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_853),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_865),
.A2(n_784),
.B1(n_805),
.B2(n_787),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_847),
.Y(n_913)
);

BUFx2_ASAP7_75t_SL g914 ( 
.A(n_834),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_855),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_847),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_846),
.A2(n_718),
.B1(n_787),
.B2(n_708),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_824),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_857),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_834),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_865),
.A2(n_791),
.B1(n_795),
.B2(n_810),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_826),
.Y(n_922)
);

BUFx2_ASAP7_75t_L g923 ( 
.A(n_824),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_861),
.A2(n_803),
.B(n_722),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_870),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_845),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_833),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_870),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_875),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_858),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_875),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_872),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_872),
.A2(n_813),
.B(n_775),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_867),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_823),
.Y(n_935)
);

CKINVDCx6p67_ASAP7_75t_R g936 ( 
.A(n_823),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_841),
.A2(n_773),
.B(n_712),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_826),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_871),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_863),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_863),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_856),
.B(n_822),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_856),
.B(n_827),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_827),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_879),
.Y(n_945)
);

INVx5_ASAP7_75t_SL g946 ( 
.A(n_942),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_893),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_893),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_929),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_929),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_942),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_931),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_SL g953 ( 
.A1(n_904),
.A2(n_873),
.B1(n_851),
.B2(n_828),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_931),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_905),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_905),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_882),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_908),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_902),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_908),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_907),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_907),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_890),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_901),
.A2(n_844),
.B(n_722),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_942),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_887),
.A2(n_835),
.B(n_860),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_885),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_885),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_915),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_915),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_882),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_919),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_886),
.A2(n_937),
.B(n_889),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_925),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_945),
.A2(n_860),
.B(n_710),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_919),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_895),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_945),
.A2(n_860),
.B(n_827),
.Y(n_978)
);

BUFx2_ASAP7_75t_SL g979 ( 
.A(n_928),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_886),
.A2(n_838),
.B(n_837),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_890),
.Y(n_981)
);

NOR2x1_ASAP7_75t_SL g982 ( 
.A(n_932),
.B(n_860),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_895),
.B(n_822),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_932),
.B(n_822),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_899),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_899),
.Y(n_986)
);

AOI221xp5_ASAP7_75t_L g987 ( 
.A1(n_966),
.A2(n_738),
.B1(n_884),
.B2(n_926),
.C(n_930),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_963),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_958),
.B(n_881),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_969),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_961),
.B(n_927),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_965),
.B(n_937),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_971),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_963),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_961),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_953),
.A2(n_851),
.B1(n_898),
.B2(n_927),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_969),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_962),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_965),
.B(n_933),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_962),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_950),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_958),
.B(n_881),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_951),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_950),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_963),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_960),
.B(n_881),
.Y(n_1006)
);

OAI211xp5_ASAP7_75t_L g1007 ( 
.A1(n_978),
.A2(n_866),
.B(n_912),
.C(n_900),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_960),
.B(n_881),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_970),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_978),
.A2(n_848),
.B1(n_897),
.B2(n_918),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_974),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_950),
.Y(n_1012)
);

AO21x2_ASAP7_75t_L g1013 ( 
.A1(n_973),
.A2(n_889),
.B(n_924),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_984),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_977),
.B(n_913),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_951),
.B(n_933),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_974),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_970),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_972),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_972),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_983),
.B(n_888),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_976),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_983),
.B(n_888),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_984),
.B(n_888),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_981),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_976),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_949),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_949),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_959),
.A2(n_921),
.B(n_917),
.Y(n_1029)
);

NAND4xp25_ASAP7_75t_L g1030 ( 
.A(n_987),
.B(n_896),
.C(n_957),
.D(n_975),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1021),
.B(n_946),
.Y(n_1031)
);

AOI21x1_ASAP7_75t_L g1032 ( 
.A1(n_1029),
.A2(n_955),
.B(n_956),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_SL g1033 ( 
.A1(n_996),
.A2(n_975),
.B(n_957),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_987),
.B(n_913),
.C(n_916),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_996),
.B(n_848),
.Y(n_1035)
);

AND2x2_ASAP7_75t_SL g1036 ( 
.A(n_1003),
.B(n_946),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1021),
.B(n_946),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_991),
.B(n_967),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_991),
.B(n_967),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1021),
.B(n_946),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1023),
.B(n_946),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1010),
.B(n_968),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1023),
.B(n_952),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_993),
.B(n_1015),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1023),
.B(n_952),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1001),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_1007),
.B(n_1029),
.C(n_1024),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_1007),
.B(n_954),
.C(n_968),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1015),
.B(n_977),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_SL g1050 ( 
.A1(n_1003),
.A2(n_982),
.B1(n_979),
.B2(n_914),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1001),
.B(n_954),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1027),
.B(n_985),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1027),
.B(n_985),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_1014),
.B(n_959),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1028),
.B(n_986),
.Y(n_1055)
);

AND2x2_ASAP7_75t_SL g1056 ( 
.A(n_1016),
.B(n_982),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_1036),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1054),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1043),
.B(n_989),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1054),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1043),
.B(n_989),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1051),
.B(n_989),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_1044),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1046),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1046),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1045),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_1051),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_1049),
.B(n_988),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1052),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1045),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1056),
.B(n_1002),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1053),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1055),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1056),
.B(n_1002),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1032),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1038),
.Y(n_1076)
);

NOR2xp67_ASAP7_75t_L g1077 ( 
.A(n_1047),
.B(n_1012),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1031),
.B(n_999),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_1048),
.B(n_1033),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1064),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1064),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1065),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1062),
.B(n_1024),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1077),
.B(n_1056),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1065),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1069),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1069),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1072),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1067),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1063),
.B(n_848),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1084),
.B(n_1071),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_1086),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1084),
.B(n_1071),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1080),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1081),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1079),
.B(n_1076),
.Y(n_1096)
);

OAI21xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1090),
.A2(n_1074),
.B(n_1071),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1087),
.B(n_1076),
.Y(n_1098)
);

INVxp67_ASAP7_75t_SL g1099 ( 
.A(n_1096),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_1091),
.B(n_1090),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1095),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1091),
.B(n_1088),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_1101),
.Y(n_1103)
);

OAI21xp33_ASAP7_75t_SL g1104 ( 
.A1(n_1100),
.A2(n_1093),
.B(n_1098),
.Y(n_1104)
);

OAI21xp33_ASAP7_75t_L g1105 ( 
.A1(n_1099),
.A2(n_1097),
.B(n_1093),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1102),
.B(n_1092),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_1102),
.B(n_1094),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1101),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1099),
.A2(n_1030),
.B1(n_1057),
.B2(n_1035),
.Y(n_1109)
);

AO32x1_ASAP7_75t_L g1110 ( 
.A1(n_1101),
.A2(n_1095),
.A3(n_1089),
.B1(n_1085),
.B2(n_1082),
.Y(n_1110)
);

OAI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1099),
.A2(n_1057),
.B1(n_1063),
.B2(n_1034),
.C(n_1050),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1099),
.B(n_1074),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1099),
.B(n_936),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_1103),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1108),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1113),
.B(n_936),
.Y(n_1116)
);

NOR2x1_ASAP7_75t_L g1117 ( 
.A(n_1107),
.B(n_935),
.Y(n_1117)
);

OAI31xp33_ASAP7_75t_SL g1118 ( 
.A1(n_1105),
.A2(n_1034),
.A3(n_1089),
.B(n_1074),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1106),
.B(n_1083),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_1112),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1110),
.Y(n_1121)
);

OAI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1104),
.A2(n_1057),
.B1(n_1042),
.B2(n_850),
.C(n_1072),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1111),
.B(n_1073),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1110),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1109),
.B(n_1073),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1107),
.B(n_1058),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_1103),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1108),
.Y(n_1128)
);

NAND2x1_ASAP7_75t_SL g1129 ( 
.A(n_1109),
.B(n_1078),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1114),
.B(n_1067),
.Y(n_1130)
);

AOI31xp33_ASAP7_75t_L g1131 ( 
.A1(n_1117),
.A2(n_1127),
.A3(n_1120),
.B(n_1116),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1121),
.A2(n_979),
.B1(n_1075),
.B2(n_1062),
.C(n_1070),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1118),
.A2(n_1078),
.B(n_1031),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_1124),
.A2(n_1075),
.B(n_1058),
.Y(n_1134)
);

AOI211xp5_ASAP7_75t_L g1135 ( 
.A1(n_1122),
.A2(n_925),
.B(n_1078),
.C(n_1075),
.Y(n_1135)
);

AOI322xp5_ASAP7_75t_L g1136 ( 
.A1(n_1123),
.A2(n_1067),
.A3(n_1061),
.B1(n_1059),
.B2(n_1070),
.C1(n_1066),
.C2(n_1036),
.Y(n_1136)
);

OAI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1124),
.A2(n_1066),
.B1(n_1070),
.B2(n_1011),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1123),
.A2(n_1036),
.B(n_1078),
.Y(n_1138)
);

NAND4xp25_ASAP7_75t_L g1139 ( 
.A(n_1115),
.B(n_1128),
.C(n_1125),
.D(n_1119),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1127),
.B(n_1058),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1126),
.B(n_1060),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1129),
.A2(n_1078),
.B1(n_1066),
.B2(n_1068),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_L g1143 ( 
.A(n_1121),
.B(n_928),
.C(n_940),
.Y(n_1143)
);

AOI31xp33_ASAP7_75t_L g1144 ( 
.A1(n_1117),
.A2(n_1037),
.A3(n_1040),
.B(n_1041),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1120),
.B(n_1060),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1117),
.A2(n_1037),
.B(n_1040),
.Y(n_1146)
);

NAND4xp75_ASAP7_75t_L g1147 ( 
.A(n_1117),
.B(n_1041),
.C(n_27),
.D(n_29),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_SL g1148 ( 
.A1(n_1121),
.A2(n_1060),
.B(n_1068),
.C(n_31),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1134),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1134),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_1131),
.B(n_934),
.C(n_939),
.Y(n_1151)
);

NOR2x1_ASAP7_75t_L g1152 ( 
.A(n_1147),
.B(n_25),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1145),
.Y(n_1153)
);

NOR3x1_ASAP7_75t_L g1154 ( 
.A(n_1139),
.B(n_923),
.C(n_918),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_L g1155 ( 
.A(n_1146),
.B(n_891),
.C(n_922),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1148),
.B(n_1059),
.Y(n_1156)
);

NOR3x1_ASAP7_75t_L g1157 ( 
.A(n_1143),
.B(n_923),
.C(n_1068),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_1144),
.B(n_891),
.C(n_894),
.Y(n_1158)
);

NAND2x1_ASAP7_75t_SL g1159 ( 
.A(n_1141),
.B(n_1059),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1140),
.Y(n_1160)
);

NOR2x1_ASAP7_75t_L g1161 ( 
.A(n_1130),
.B(n_1137),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1133),
.B(n_30),
.Y(n_1162)
);

NOR3x1_ASAP7_75t_L g1163 ( 
.A(n_1138),
.B(n_897),
.C(n_1039),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_SL g1164 ( 
.A(n_1135),
.B(n_891),
.C(n_31),
.Y(n_1164)
);

OAI211xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1136),
.A2(n_30),
.B(n_32),
.C(n_34),
.Y(n_1165)
);

AOI211xp5_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_1142),
.B(n_1132),
.C(n_37),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1162),
.A2(n_1011),
.B1(n_1017),
.B2(n_1016),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_1164),
.B(n_922),
.C(n_894),
.Y(n_1168)
);

OAI211xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1161),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_1152),
.B(n_939),
.C(n_934),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1153),
.B(n_1160),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1149),
.B(n_938),
.C(n_922),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1151),
.A2(n_1156),
.B1(n_1150),
.B2(n_1155),
.C(n_1158),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1156),
.B(n_35),
.C(n_36),
.Y(n_1174)
);

NAND4xp25_ASAP7_75t_L g1175 ( 
.A(n_1154),
.B(n_1011),
.C(n_1017),
.D(n_894),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_SL g1176 ( 
.A(n_1159),
.B(n_39),
.C(n_40),
.Y(n_1176)
);

NOR4xp25_ASAP7_75t_L g1177 ( 
.A(n_1157),
.B(n_39),
.C(n_43),
.D(n_44),
.Y(n_1177)
);

NOR2x1_ASAP7_75t_L g1178 ( 
.A(n_1163),
.B(n_43),
.Y(n_1178)
);

OAI211xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1161),
.A2(n_938),
.B(n_916),
.C(n_941),
.Y(n_1179)
);

XNOR2xp5_ASAP7_75t_L g1180 ( 
.A(n_1152),
.B(n_943),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1152),
.B(n_1061),
.Y(n_1181)
);

OAI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1165),
.A2(n_1017),
.B1(n_914),
.B2(n_1032),
.C(n_938),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_SL g1183 ( 
.A(n_1162),
.B(n_838),
.C(n_1061),
.Y(n_1183)
);

NAND5xp2_ASAP7_75t_L g1184 ( 
.A(n_1160),
.B(n_911),
.C(n_986),
.D(n_1028),
.E(n_910),
.Y(n_1184)
);

OAI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_1165),
.A2(n_911),
.B1(n_1026),
.B2(n_1022),
.C(n_1020),
.Y(n_1185)
);

OAI211xp5_ASAP7_75t_L g1186 ( 
.A1(n_1165),
.A2(n_903),
.B(n_854),
.C(n_837),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1162),
.B(n_941),
.C(n_943),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_L g1188 ( 
.A(n_1162),
.B(n_854),
.C(n_837),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1149),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1166),
.B(n_990),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1189),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1169),
.A2(n_1016),
.B1(n_943),
.B2(n_999),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1181),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1186),
.A2(n_1016),
.B1(n_999),
.B2(n_992),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1171),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1180),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1176),
.A2(n_1016),
.B1(n_999),
.B2(n_992),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1170),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1174),
.Y(n_1199)
);

NOR2x1_ASAP7_75t_L g1200 ( 
.A(n_1179),
.B(n_854),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1178),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1187),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_L g1203 ( 
.A(n_1182),
.B(n_964),
.Y(n_1203)
);

NOR2xp67_ASAP7_75t_L g1204 ( 
.A(n_1172),
.B(n_48),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1173),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1185),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1184),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1168),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1183),
.A2(n_999),
.B1(n_992),
.B2(n_964),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1177),
.A2(n_964),
.B1(n_903),
.B2(n_1013),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1188),
.Y(n_1211)
);

NOR3xp33_ASAP7_75t_L g1212 ( 
.A(n_1175),
.B(n_944),
.C(n_910),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1167),
.A2(n_1026),
.B1(n_990),
.B2(n_1022),
.Y(n_1213)
);

NAND4xp75_ASAP7_75t_L g1214 ( 
.A(n_1205),
.B(n_51),
.C(n_53),
.D(n_54),
.Y(n_1214)
);

AND3x4_ASAP7_75t_L g1215 ( 
.A(n_1196),
.B(n_1204),
.C(n_1212),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1201),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1193),
.B(n_1014),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1199),
.B(n_997),
.Y(n_1218)
);

NOR2x1_ASAP7_75t_L g1219 ( 
.A(n_1191),
.B(n_964),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_L g1220 ( 
.A(n_1195),
.B(n_997),
.C(n_1020),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1198),
.Y(n_1221)
);

NOR4xp75_ASAP7_75t_SL g1222 ( 
.A(n_1190),
.B(n_903),
.C(n_920),
.D(n_109),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1211),
.B(n_944),
.Y(n_1223)
);

NAND4xp75_ASAP7_75t_L g1224 ( 
.A(n_1206),
.B(n_1002),
.C(n_1008),
.D(n_1006),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1208),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_L g1226 ( 
.A(n_1197),
.B(n_107),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1202),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1207),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1200),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1210),
.A2(n_1203),
.B(n_1213),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1210),
.B(n_1019),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1192),
.B(n_1009),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1209),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1194),
.B(n_1019),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1201),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1216),
.B(n_1000),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1235),
.B(n_903),
.Y(n_1237)
);

NOR3xp33_ASAP7_75t_L g1238 ( 
.A(n_1228),
.B(n_944),
.C(n_992),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1227),
.B(n_998),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1227),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1215),
.A2(n_992),
.B1(n_1018),
.B2(n_1009),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1225),
.B(n_1018),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1221),
.B(n_1000),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1226),
.A2(n_980),
.B(n_973),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1217),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1229),
.A2(n_995),
.B1(n_998),
.B2(n_1004),
.Y(n_1246)
);

XOR2xp5_ASAP7_75t_L g1247 ( 
.A(n_1214),
.B(n_108),
.Y(n_1247)
);

NOR3xp33_ASAP7_75t_L g1248 ( 
.A(n_1233),
.B(n_909),
.C(n_112),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1214),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1223),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1245),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1240),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1249),
.A2(n_1224),
.B1(n_1218),
.B2(n_1230),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1239),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1247),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1243),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1236),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1242),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1250),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1241),
.A2(n_1232),
.B1(n_1231),
.B2(n_1220),
.Y(n_1260)
);

AO22x2_ASAP7_75t_L g1261 ( 
.A1(n_1248),
.A2(n_1222),
.B1(n_1234),
.B2(n_1219),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1237),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1237),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1244),
.A2(n_995),
.B1(n_909),
.B2(n_1004),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1246),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1251),
.B(n_1238),
.Y(n_1266)
);

NOR3x2_ASAP7_75t_L g1267 ( 
.A(n_1255),
.B(n_111),
.C(n_117),
.Y(n_1267)
);

NAND4xp25_ASAP7_75t_L g1268 ( 
.A(n_1253),
.B(n_120),
.C(n_121),
.D(n_124),
.Y(n_1268)
);

AOI221xp5_ASAP7_75t_L g1269 ( 
.A1(n_1259),
.A2(n_852),
.B1(n_1012),
.B2(n_947),
.C(n_948),
.Y(n_1269)
);

NOR2x1_ASAP7_75t_L g1270 ( 
.A(n_1252),
.B(n_128),
.Y(n_1270)
);

XOR2x2_ASAP7_75t_L g1271 ( 
.A(n_1258),
.B(n_129),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1265),
.A2(n_1263),
.B1(n_1262),
.B2(n_1261),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1256),
.B(n_130),
.C(n_131),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1254),
.A2(n_906),
.B1(n_892),
.B2(n_883),
.Y(n_1274)
);

OAI211xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1257),
.A2(n_132),
.B(n_134),
.C(n_135),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1272),
.A2(n_1260),
.B(n_1264),
.Y(n_1276)
);

AO22x2_ASAP7_75t_L g1277 ( 
.A1(n_1266),
.A2(n_1025),
.B1(n_988),
.B2(n_994),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1270),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1267),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1268),
.A2(n_852),
.B1(n_1008),
.B2(n_1006),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1271),
.A2(n_1275),
.B1(n_1273),
.B2(n_1274),
.Y(n_1281)
);

OA21x2_ASAP7_75t_L g1282 ( 
.A1(n_1278),
.A2(n_1279),
.B(n_1281),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1276),
.A2(n_1269),
.B1(n_1008),
.B2(n_1006),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1280),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1277),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1282),
.A2(n_138),
.B(n_140),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1286),
.A2(n_1283),
.B1(n_1284),
.B2(n_1285),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1287),
.A2(n_1013),
.B1(n_920),
.B2(n_1005),
.Y(n_1288)
);

AOI221xp5_ASAP7_75t_L g1289 ( 
.A1(n_1288),
.A2(n_142),
.B1(n_166),
.B2(n_948),
.C(n_947),
.Y(n_1289)
);

AOI211xp5_ASAP7_75t_L g1290 ( 
.A1(n_1289),
.A2(n_980),
.B(n_883),
.C(n_880),
.Y(n_1290)
);


endmodule