module fake_jpeg_11011_n_402 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_402);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_402;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_10),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_68),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_22),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_47),
.A2(n_71),
.B1(n_42),
.B2(n_32),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_12),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_64),
.B(n_39),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_79),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_36),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_28),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_90),
.B(n_102),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_95),
.A2(n_114),
.B1(n_42),
.B2(n_32),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_100),
.B(n_111),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_37),
.B1(n_30),
.B2(n_31),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_103),
.A2(n_31),
.B1(n_99),
.B2(n_94),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_104),
.B(n_105),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_29),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_79),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2x1_ASAP7_75t_SL g126 ( 
.A(n_57),
.B(n_37),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_37),
.B(n_42),
.C(n_32),
.Y(n_143)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_25),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_21),
.B1(n_43),
.B2(n_59),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_48),
.B1(n_43),
.B2(n_76),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_150),
.Y(n_176)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_45),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_137),
.B(n_152),
.Y(n_208)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_51),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_171),
.Y(n_200)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_145),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_146),
.A2(n_153),
.B1(n_160),
.B2(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_45),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_43),
.B1(n_23),
.B2(n_26),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_169),
.Y(n_192)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_126),
.B1(n_116),
.B2(n_113),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_163),
.B1(n_107),
.B2(n_122),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_26),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_172),
.C(n_174),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_161),
.B1(n_166),
.B2(n_167),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_77),
.B1(n_74),
.B2(n_48),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_72),
.B1(n_65),
.B2(n_60),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_40),
.B1(n_31),
.B2(n_71),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_99),
.A2(n_31),
.B1(n_79),
.B2(n_3),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_98),
.A2(n_91),
.B1(n_122),
.B2(n_119),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_86),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_87),
.B(n_0),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_92),
.B(n_0),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_154),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_119),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_206),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_191),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_136),
.B1(n_143),
.B2(n_140),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_186),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_134),
.A2(n_93),
.B(n_97),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_189),
.B(n_172),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_97),
.B(n_132),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_91),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_164),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_196),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_157),
.A2(n_174),
.B1(n_172),
.B2(n_141),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_201),
.A2(n_202),
.B1(n_163),
.B2(n_106),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_127),
.B1(n_108),
.B2(n_106),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_149),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_0),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_127),
.C(n_108),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_218),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_150),
.B1(n_171),
.B2(n_169),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_148),
.B1(n_155),
.B2(n_162),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_213),
.A2(n_217),
.B(n_237),
.Y(n_261)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_185),
.B1(n_188),
.B2(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_216),
.B(n_231),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_200),
.A2(n_135),
.B(n_156),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_196),
.B1(n_202),
.B2(n_208),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_151),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_221),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_170),
.B(n_145),
.C(n_139),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_178),
.A2(n_138),
.B1(n_142),
.B2(n_144),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_224),
.A2(n_227),
.B1(n_238),
.B2(n_195),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_233),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_192),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_1),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_183),
.C(n_177),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_1),
.B(n_5),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_240),
.B1(n_248),
.B2(n_220),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_185),
.B1(n_206),
.B2(n_204),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_241),
.B(n_254),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_218),
.A2(n_178),
.B1(n_176),
.B2(n_194),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_249),
.B(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_176),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_264),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_236),
.B1(n_227),
.B2(n_223),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_225),
.A2(n_176),
.B1(n_194),
.B2(n_182),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_217),
.B(n_237),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_192),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_259),
.Y(n_270)
);

AND2x6_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_207),
.Y(n_251)
);

AOI32xp33_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_190),
.A3(n_192),
.B1(n_198),
.B2(n_183),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_190),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_198),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_212),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_230),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_235),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_182),
.B(n_209),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_243),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_210),
.B1(n_234),
.B2(n_232),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_268),
.B1(n_285),
.B2(n_240),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_273),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_262),
.A2(n_256),
.B1(n_261),
.B2(n_242),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_269),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_247),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_274),
.A2(n_288),
.B1(n_228),
.B2(n_226),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_243),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_290),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_239),
.A2(n_211),
.B1(n_221),
.B2(n_220),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_235),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_248),
.C(n_257),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_292),
.A2(n_302),
.B1(n_305),
.B2(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_250),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_300),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_297),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_275),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_249),
.B1(n_251),
.B2(n_221),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_272),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_307),
.C(n_311),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_268),
.A2(n_261),
.B1(n_252),
.B2(n_259),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_264),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_260),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_263),
.Y(n_310)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_263),
.C(n_226),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_11),
.B1(n_15),
.B2(n_13),
.Y(n_332)
);

OAI31xp33_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_236),
.A3(n_179),
.B(n_227),
.Y(n_313)
);

FAx1_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_266),
.CI(n_275),
.CON(n_318),
.SN(n_318)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_295),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_316),
.B(n_317),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_219),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_305),
.B(n_302),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_319),
.A2(n_299),
.B1(n_296),
.B2(n_310),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_271),
.Y(n_320)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_287),
.B1(n_279),
.B2(n_280),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_323),
.A2(n_330),
.B1(n_332),
.B2(n_296),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_282),
.C(n_283),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_314),
.C(n_315),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_281),
.Y(n_327)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_327),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_236),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_328),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_179),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_292),
.B1(n_301),
.B2(n_304),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_299),
.A2(n_277),
.B1(n_209),
.B2(n_13),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_333),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_334),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_346),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_319),
.A2(n_322),
.B1(n_320),
.B2(n_326),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_323),
.A2(n_294),
.B1(n_308),
.B2(n_304),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_321),
.A2(n_331),
.B1(n_332),
.B2(n_330),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_326),
.A2(n_298),
.B1(n_306),
.B2(n_313),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_318),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_307),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_331),
.A2(n_298),
.B(n_306),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_318),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_11),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_325),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_325),
.C(n_327),
.Y(n_358)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_347),
.Y(n_351)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_344),
.Y(n_352)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_352),
.Y(n_373)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_356),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_358),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_345),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_361),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_360),
.A2(n_357),
.B1(n_336),
.B2(n_334),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_349),
.C(n_346),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_16),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_363),
.B1(n_357),
.B2(n_338),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_366),
.A2(n_372),
.B1(n_6),
.B2(n_7),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_6),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_338),
.B(n_333),
.Y(n_369)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_369),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_350),
.A2(n_342),
.B1(n_341),
.B2(n_335),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_348),
.Y(n_374)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_373),
.A2(n_363),
.B1(n_13),
.B2(n_15),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_376),
.B(n_379),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_380),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_370),
.Y(n_378)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_6),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_382),
.B(n_383),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_9),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_366),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_369),
.C(n_8),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_L g386 ( 
.A1(n_378),
.A2(n_371),
.B(n_365),
.C(n_364),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_386),
.B(n_387),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_381),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_383),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_393),
.B(n_394),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_375),
.C(n_380),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_382),
.C(n_8),
.Y(n_395)
);

NOR3xp33_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_390),
.C(n_389),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_397),
.A2(n_396),
.B(n_389),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_L g399 ( 
.A(n_398),
.B(n_392),
.C(n_8),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_399),
.B(n_7),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_400),
.A2(n_7),
.B1(n_9),
.B2(n_331),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_7),
.Y(n_402)
);


endmodule