module fake_jpeg_31261_n_549 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_549);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_549;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_60),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_59),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_17),
.B(n_0),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_61),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_54),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_67),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_72),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_73),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_81),
.Y(n_137)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_89),
.Y(n_177)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_100),
.Y(n_168)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_112),
.Y(n_119)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_50),
.B1(n_36),
.B2(n_43),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_48),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_124),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_48),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_23),
.B1(n_53),
.B2(n_52),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_129),
.A2(n_132),
.B1(n_32),
.B2(n_27),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_63),
.B(n_54),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_130),
.B(n_149),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_58),
.A2(n_35),
.B1(n_30),
.B2(n_53),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_55),
.A2(n_47),
.B(n_36),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_37),
.C(n_29),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_36),
.B1(n_52),
.B2(n_49),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_142),
.A2(n_178),
.B1(n_31),
.B2(n_25),
.Y(n_226)
);

BUFx12_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_76),
.B(n_30),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_165),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_79),
.A2(n_49),
.B(n_27),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_81),
.B(n_35),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_36),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_62),
.A2(n_73),
.B1(n_70),
.B2(n_64),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_179),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_191),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_181),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_182),
.B(n_186),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_32),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_187),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_185),
.B(n_204),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_122),
.B(n_23),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_37),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_129),
.A2(n_71),
.B1(n_29),
.B2(n_75),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_194),
.B(n_144),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_122),
.A2(n_93),
.B(n_47),
.C(n_89),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_198),
.A2(n_226),
.B1(n_126),
.B2(n_116),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_199),
.B(n_224),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_139),
.A2(n_145),
.B1(n_166),
.B2(n_158),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_200),
.A2(n_159),
.B1(n_151),
.B2(n_123),
.Y(n_267)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_113),
.A2(n_111),
.B1(n_110),
.B2(n_94),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_203),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_137),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_74),
.B1(n_99),
.B2(n_95),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_213),
.Y(n_272)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_215),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_228),
.B1(n_168),
.B2(n_123),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_142),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_229),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_115),
.A2(n_105),
.B1(n_84),
.B2(n_82),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_115),
.B(n_47),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_127),
.A2(n_31),
.B1(n_25),
.B2(n_47),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_150),
.A2(n_31),
.B1(n_25),
.B2(n_47),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_1),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_138),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_225),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_145),
.A2(n_56),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_227),
.A2(n_159),
.B1(n_151),
.B2(n_133),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_117),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_231),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_138),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_233),
.Y(n_271)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_236),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_153),
.B(n_4),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_154),
.Y(n_262)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_167),
.C(n_143),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_8),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_192),
.A2(n_128),
.B1(n_170),
.B2(n_163),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_240),
.A2(n_267),
.B1(n_276),
.B2(n_221),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_168),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_243),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_279),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_264),
.A2(n_219),
.B(n_202),
.Y(n_312)
);

AO22x2_ASAP7_75t_L g265 ( 
.A1(n_198),
.A2(n_170),
.B1(n_163),
.B2(n_154),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g298 ( 
.A1(n_265),
.A2(n_280),
.B1(n_213),
.B2(n_236),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_192),
.A2(n_176),
.B1(n_125),
.B2(n_140),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_205),
.B1(n_179),
.B2(n_208),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_7),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_281),
.A2(n_298),
.B1(n_301),
.B2(n_265),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_261),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_280),
.B1(n_251),
.B2(n_265),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_299),
.B1(n_305),
.B2(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_220),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_287),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_187),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_184),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_289),
.B(n_295),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_302),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_237),
.A2(n_210),
.B1(n_204),
.B2(n_218),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_291),
.A2(n_293),
.B1(n_268),
.B2(n_239),
.Y(n_316)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_237),
.A2(n_222),
.B1(n_194),
.B2(n_191),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_277),
.B1(n_274),
.B2(n_250),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_246),
.B(n_207),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_235),
.B1(n_181),
.B2(n_215),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_243),
.A2(n_212),
.B1(n_189),
.B2(n_233),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_238),
.B(n_193),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_308),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_190),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_304),
.B(n_312),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_280),
.A2(n_229),
.B1(n_225),
.B2(n_234),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_265),
.A2(n_230),
.B1(n_216),
.B2(n_206),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_263),
.A2(n_201),
.B(n_116),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_307),
.A2(n_257),
.B(n_260),
.Y(n_342)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_219),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_314),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_249),
.B(n_7),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_315),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_242),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_322),
.B1(n_328),
.B2(n_332),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_311),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_319),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_321),
.A2(n_342),
.B(n_297),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_293),
.A2(n_268),
.B1(n_265),
.B2(n_252),
.Y(n_322)
);

BUFx12_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_257),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_244),
.C(n_249),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_283),
.C(n_315),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_327),
.A2(n_330),
.B1(n_334),
.B2(n_320),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_291),
.A2(n_252),
.B1(n_244),
.B2(n_240),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_285),
.A2(n_244),
.B1(n_276),
.B2(n_259),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_281),
.A2(n_259),
.B1(n_272),
.B2(n_245),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_299),
.A2(n_272),
.B1(n_245),
.B2(n_271),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_284),
.A2(n_255),
.B1(n_270),
.B2(n_258),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_337),
.A2(n_306),
.B1(n_305),
.B2(n_328),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_338),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_307),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_340),
.B(n_298),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_258),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_344),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_289),
.B(n_260),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_296),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_342),
.A2(n_288),
.B(n_312),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_347),
.A2(n_349),
.B(n_340),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_350),
.A2(n_359),
.B1(n_332),
.B2(n_337),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_351),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_336),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_358),
.Y(n_379)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_367),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_357),
.B(n_368),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_320),
.A2(n_298),
.B1(n_303),
.B2(n_287),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_360),
.Y(n_399)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_313),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_364),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_326),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_317),
.B(n_295),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_365),
.B(n_366),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_242),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_310),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_309),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_324),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_370),
.Y(n_385)
);

BUFx24_ASAP7_75t_SL g371 ( 
.A(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_371),
.B(n_373),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_329),
.B(n_302),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_326),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_L g373 ( 
.A(n_324),
.B(n_308),
.C(n_300),
.Y(n_373)
);

INVx8_ASAP7_75t_L g374 ( 
.A(n_318),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_339),
.Y(n_375)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_375),
.Y(n_382)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_376),
.Y(n_383)
);

INVx5_ASAP7_75t_SL g384 ( 
.A(n_348),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_331),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_338),
.Y(n_386)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_352),
.A2(n_330),
.B1(n_334),
.B2(n_316),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_387),
.A2(n_372),
.B1(n_368),
.B2(n_298),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_347),
.A2(n_342),
.B(n_322),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_388),
.B(n_349),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_351),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_394),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_352),
.B1(n_358),
.B2(n_359),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_361),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_364),
.B(n_335),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_397),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_350),
.A2(n_369),
.B1(n_375),
.B2(n_362),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_335),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_398),
.A2(n_331),
.B(n_343),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_404),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_361),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_407),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_411),
.A2(n_425),
.B1(n_426),
.B2(n_298),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g460 ( 
.A(n_412),
.B(n_435),
.Y(n_460)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_344),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_415),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_399),
.B(n_319),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_436),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_406),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_418),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_355),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_386),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_420),
.A2(n_423),
.B(n_428),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_389),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_424),
.A2(n_398),
.B(n_379),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_298),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_346),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_427),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_393),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_381),
.B(n_370),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_432),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_343),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_402),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_433),
.A2(n_434),
.B1(n_420),
.B2(n_414),
.Y(n_437)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_382),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_345),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_385),
.B(n_345),
.Y(n_436)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_409),
.A2(n_391),
.B1(n_379),
.B2(n_380),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_438),
.A2(n_459),
.B1(n_434),
.B2(n_410),
.Y(n_461)
);

FAx1_ASAP7_75t_SL g441 ( 
.A(n_418),
.B(n_395),
.CI(n_397),
.CON(n_441),
.SN(n_441)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_392),
.C(n_400),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_447),
.C(n_448),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_446),
.B(n_454),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_408),
.B(n_392),
.C(n_400),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_357),
.C(n_403),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_415),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_387),
.C(n_388),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_453),
.C(n_425),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_417),
.C(n_416),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_412),
.B(n_380),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_405),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_458),
.Y(n_470)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_423),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_457),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_432),
.B(n_377),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_468),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_428),
.C(n_422),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_462),
.B(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_419),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_422),
.C(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_472),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_450),
.A2(n_425),
.B1(n_435),
.B2(n_427),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_469),
.A2(n_456),
.B1(n_444),
.B2(n_459),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_424),
.C(n_436),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g484 ( 
.A(n_471),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_430),
.C(n_421),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_442),
.Y(n_473)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_421),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_478),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_430),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_460),
.B(n_383),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_479),
.B(n_455),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_383),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_439),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_482),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_455),
.C(n_444),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_466),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_467),
.B(n_440),
.C(n_441),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_492),
.Y(n_508)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_476),
.Y(n_491)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_491),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_441),
.C(n_451),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_452),
.B1(n_449),
.B2(n_407),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_495),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_323),
.Y(n_504)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_475),
.B(n_458),
.C(n_378),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_498),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_470),
.B(n_478),
.C(n_466),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_484),
.B(n_470),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_504),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_485),
.A2(n_477),
.B1(n_471),
.B2(n_479),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_500),
.A2(n_248),
.B1(n_11),
.B2(n_12),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_501),
.B(n_512),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_486),
.B(n_318),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_506),
.B(n_509),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_489),
.B(n_374),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_483),
.B(n_378),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_513),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_488),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_256),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_323),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_323),
.Y(n_513)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_497),
.B(n_250),
.CI(n_253),
.CON(n_514),
.SN(n_514)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_277),
.C(n_256),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_508),
.A2(n_492),
.B(n_498),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_515),
.A2(n_523),
.B(n_10),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_490),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_516),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_502),
.A2(n_483),
.B1(n_487),
.B2(n_253),
.Y(n_517)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_517),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_519),
.A2(n_526),
.B(n_248),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_522),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_511),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_505),
.C(n_501),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_527),
.B(n_531),
.C(n_533),
.Y(n_538)
);

NAND4xp25_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_514),
.C(n_503),
.D(n_504),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_528),
.A2(n_533),
.B(n_527),
.Y(n_537)
);

XNOR2x1_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_521),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_518),
.C(n_525),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_535),
.B(n_532),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_529),
.A2(n_526),
.B(n_12),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_536),
.A2(n_537),
.B(n_539),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_534),
.A2(n_11),
.B(n_13),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_540),
.A2(n_542),
.B(n_14),
.Y(n_544)
);

AOI21x1_ASAP7_75t_L g542 ( 
.A1(n_538),
.A2(n_11),
.B(n_13),
.Y(n_542)
);

OAI31xp33_ASAP7_75t_SL g543 ( 
.A1(n_541),
.A2(n_11),
.A3(n_13),
.B(n_14),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_543),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_544),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_14),
.B(n_15),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_15),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_15),
.Y(n_549)
);


endmodule