module fake_netlist_1_5129_n_533 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_533);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_533;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_29), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_23), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_45), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_63), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_56), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_73), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_10), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_67), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_57), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_70), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_19), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_69), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_3), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_24), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_50), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_11), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_39), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_16), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_36), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_9), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_18), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_52), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_44), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_8), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_33), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_75), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_0), .B(n_47), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_13), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_48), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_12), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_41), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_17), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_43), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_46), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_99), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_81), .Y(n_115) );
NAND2x1_ASAP7_75t_L g116 ( .A(n_90), .B(n_0), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_99), .Y(n_117) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_79), .B(n_31), .Y(n_118) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_100), .A2(n_30), .B(n_74), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_100), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_84), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_85), .A2(n_28), .B(n_72), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_104), .B(n_1), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_102), .B(n_1), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_102), .B(n_2), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_121), .B(n_94), .Y(n_136) );
INVx4_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_115), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_121), .B(n_78), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_122), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_119), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_122), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_119), .Y(n_143) );
BUFx4f_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_122), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_120), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_123), .B(n_98), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_123), .B(n_83), .Y(n_148) );
INVxp67_ASAP7_75t_L g149 ( .A(n_129), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
INVx3_ASAP7_75t_R g151 ( .A(n_135), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_124), .B(n_103), .Y(n_152) );
INVx2_ASAP7_75t_SL g153 ( .A(n_124), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_125), .B(n_95), .Y(n_154) );
INVx5_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_125), .B(n_109), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_126), .B(n_97), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_126), .B(n_97), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_114), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_160), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_138), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_154), .B(n_127), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_154), .B(n_149), .Y(n_168) );
NOR2xp33_ASAP7_75t_SL g169 ( .A(n_137), .B(n_82), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_139), .B(n_127), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_153), .B(n_132), .Y(n_171) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_153), .B(n_132), .Y(n_176) );
INVx1_ASAP7_75t_SL g177 ( .A(n_156), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
NOR2xp67_ASAP7_75t_L g181 ( .A(n_137), .B(n_158), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_159), .B(n_134), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_146), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_157), .B(n_134), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_144), .B(n_130), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_137), .A2(n_116), .B1(n_131), .B2(n_107), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_157), .B(n_135), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_137), .A2(n_116), .B1(n_90), .B2(n_114), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_157), .B(n_114), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
OR2x6_ASAP7_75t_L g192 ( .A(n_158), .B(n_128), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_179), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_173), .B(n_158), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_183), .Y(n_196) );
AOI221xp5_ASAP7_75t_L g197 ( .A1(n_168), .A2(n_158), .B1(n_144), .B2(n_159), .C(n_157), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_172), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
BUFx12f_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_184), .A2(n_144), .B1(n_160), .B2(n_147), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_182), .B(n_144), .Y(n_204) );
BUFx2_ASAP7_75t_SL g205 ( .A(n_173), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_172), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_172), .B(n_160), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_162), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_177), .B(n_136), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_165), .B(n_160), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_180), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_SL g212 ( .A1(n_185), .A2(n_141), .B(n_143), .C(n_136), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_191), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_170), .A2(n_147), .B(n_148), .C(n_117), .Y(n_214) );
AOI21x1_ASAP7_75t_L g215 ( .A1(n_192), .A2(n_143), .B(n_141), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_161), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_171), .A2(n_141), .B(n_143), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_191), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_165), .B(n_93), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
AOI221xp5_ASAP7_75t_L g222 ( .A1(n_174), .A2(n_148), .B1(n_133), .B2(n_117), .C(n_120), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_188), .B(n_148), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_176), .A2(n_128), .B(n_89), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_196), .Y(n_225) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_215), .A2(n_112), .B(n_96), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_196), .Y(n_227) );
OAI21x1_ASAP7_75t_L g228 ( .A1(n_215), .A2(n_181), .B(n_167), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_198), .Y(n_229) );
INVx6_ASAP7_75t_L g230 ( .A(n_206), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_198), .Y(n_231) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_224), .A2(n_112), .B(n_101), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_213), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_213), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_219), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_194), .Y(n_237) );
NOR3xp33_ASAP7_75t_SL g238 ( .A(n_220), .B(n_187), .C(n_190), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_193), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_204), .A2(n_164), .B1(n_178), .B2(n_167), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_218), .A2(n_164), .B(n_178), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_209), .B(n_186), .Y(n_242) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_212), .A2(n_91), .B(n_108), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_203), .A2(n_180), .B(n_166), .Y(n_244) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_193), .A2(n_108), .B(n_103), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_214), .A2(n_163), .B(n_166), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_202), .A2(n_175), .B(n_91), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_202), .A2(n_192), .B1(n_175), .B2(n_189), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_221), .A2(n_96), .B(n_101), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_242), .B(n_209), .Y(n_251) );
INVx5_ASAP7_75t_SL g252 ( .A(n_225), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_246), .A2(n_197), .B(n_223), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_248), .A2(n_200), .B1(n_208), .B2(n_201), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_242), .A2(n_204), .B1(n_208), .B2(n_195), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_238), .B(n_201), .Y(n_257) );
BUFx8_ASAP7_75t_L g258 ( .A(n_237), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_225), .Y(n_259) );
CKINVDCx6p67_ASAP7_75t_R g260 ( .A(n_227), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_248), .A2(n_192), .B(n_221), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_228), .A2(n_192), .B(n_221), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_238), .B(n_210), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_249), .Y(n_264) );
AOI22xp33_ASAP7_75t_SL g265 ( .A1(n_237), .A2(n_205), .B1(n_194), .B2(n_207), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_249), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_237), .A2(n_222), .B1(n_194), .B2(n_152), .Y(n_267) );
OAI21xp33_ASAP7_75t_SL g268 ( .A1(n_233), .A2(n_194), .B(n_216), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_240), .A2(n_152), .B1(n_205), .B2(n_217), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_228), .A2(n_189), .B(n_216), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_240), .A2(n_217), .B1(n_207), .B2(n_206), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_239), .A2(n_207), .B1(n_206), .B2(n_199), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_251), .B(n_233), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_264), .B(n_239), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_268), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_266), .Y(n_276) );
INVx8_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_259), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_259), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_254), .B(n_235), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_252), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_260), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_252), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_258), .Y(n_284) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_261), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_252), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_253), .B(n_225), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_258), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_270), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_261), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_256), .B(n_229), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_270), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_263), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_262), .Y(n_294) );
AO31x2_ASAP7_75t_L g295 ( .A1(n_289), .A2(n_262), .A3(n_272), .B(n_239), .Y(n_295) );
OAI33xp33_ASAP7_75t_L g296 ( .A1(n_276), .A2(n_255), .A3(n_111), .B1(n_86), .B2(n_271), .B3(n_235), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_287), .B(n_229), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_293), .A2(n_257), .B1(n_133), .B2(n_106), .C(n_111), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_282), .B(n_113), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_273), .B(n_236), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_273), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_289), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
INVxp67_ASAP7_75t_SL g306 ( .A(n_280), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_292), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_287), .B(n_229), .Y(n_308) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_292), .A2(n_228), .B(n_243), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g310 ( .A1(n_293), .A2(n_133), .B1(n_236), .B2(n_267), .C(n_155), .Y(n_310) );
OAI33xp33_ASAP7_75t_L g311 ( .A1(n_293), .A2(n_2), .A3(n_3), .B1(n_4), .B2(n_5), .B3(n_6), .Y(n_311) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_282), .A2(n_265), .B1(n_269), .B2(n_245), .C(n_231), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_291), .B(n_231), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_291), .B(n_231), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_291), .B(n_234), .Y(n_316) );
NAND3xp33_ASAP7_75t_L g317 ( .A(n_294), .B(n_245), .C(n_232), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_275), .B(n_234), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_278), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_277), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_274), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_303), .B(n_274), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_301), .Y(n_325) );
OAI322xp33_ASAP7_75t_L g326 ( .A1(n_301), .A2(n_290), .A3(n_285), .B1(n_288), .B2(n_294), .C1(n_283), .C2(n_281), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_319), .B(n_282), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_302), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_306), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_322), .Y(n_331) );
BUFx2_ASAP7_75t_SL g332 ( .A(n_321), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_322), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_313), .B(n_288), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_296), .B(n_288), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_313), .B(n_285), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_298), .B(n_284), .Y(n_338) );
AND2x4_ASAP7_75t_SL g339 ( .A(n_321), .B(n_286), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_298), .B(n_284), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_308), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
AND2x4_ASAP7_75t_SL g344 ( .A(n_321), .B(n_286), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_284), .Y(n_345) );
NAND5xp2_ASAP7_75t_L g346 ( .A(n_299), .B(n_290), .C(n_279), .D(n_286), .E(n_7), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_318), .B(n_279), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_297), .B(n_283), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_315), .B(n_283), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_316), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_314), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_318), .B(n_278), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_307), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_307), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_318), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_297), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_321), .B(n_286), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_295), .B(n_281), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_317), .Y(n_364) );
AND2x2_ASAP7_75t_SL g365 ( .A(n_305), .B(n_281), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g366 ( .A(n_300), .B(n_245), .C(n_232), .Y(n_366) );
AOI211xp5_ASAP7_75t_SL g367 ( .A1(n_326), .A2(n_312), .B(n_310), .C(n_305), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_328), .B(n_309), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g369 ( .A(n_362), .B(n_278), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_331), .B(n_309), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_333), .B(n_309), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_327), .B(n_305), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_364), .B(n_317), .C(n_245), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_325), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_324), .B(n_295), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_350), .B(n_320), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_342), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_338), .B(n_295), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_354), .B(n_295), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_356), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_337), .B(n_295), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_340), .B(n_320), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_341), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_347), .B(n_320), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_337), .B(n_323), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_352), .B(n_323), .Y(n_390) );
AND3x2_ASAP7_75t_L g391 ( .A(n_336), .B(n_311), .C(n_234), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_353), .B(n_277), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_357), .Y(n_394) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_349), .B(n_4), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_360), .B(n_245), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_330), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_330), .B(n_277), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_336), .A2(n_332), .B1(n_344), .B2(n_339), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_334), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_348), .B(n_278), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_334), .B(n_243), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_358), .B(n_278), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_348), .B(n_5), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_365), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_348), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_339), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_344), .A2(n_243), .B1(n_232), .B2(n_277), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_359), .B(n_6), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g410 ( .A1(n_346), .A2(n_250), .B(n_92), .C(n_105), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_351), .B(n_232), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_365), .B(n_7), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_351), .Y(n_413) );
NOR3xp33_ASAP7_75t_L g414 ( .A(n_366), .B(n_250), .C(n_247), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_349), .B(n_277), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_363), .B(n_277), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_361), .B(n_243), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_361), .Y(n_418) );
NAND4xp75_ASAP7_75t_L g419 ( .A(n_399), .B(n_232), .C(n_226), .D(n_355), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_418), .B(n_343), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_375), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_383), .B(n_343), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_395), .A2(n_355), .B(n_343), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_381), .B(n_343), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_394), .B(n_355), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_378), .B(n_226), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_373), .A2(n_226), .B(n_247), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_412), .A2(n_8), .B(n_9), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_404), .A2(n_10), .B(n_11), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_407), .B(n_12), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_392), .Y(n_433) );
AOI32xp33_ASAP7_75t_L g434 ( .A1(n_410), .A2(n_250), .A3(n_247), .B1(n_246), .B2(n_244), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_370), .B(n_226), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_374), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_379), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_385), .A2(n_155), .B1(n_13), .B2(n_14), .C1(n_246), .C2(n_244), .Y(n_438) );
NOR2x1_ASAP7_75t_L g439 ( .A(n_415), .B(n_226), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_385), .A2(n_110), .B1(n_87), .B2(n_155), .C(n_14), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_406), .B(n_244), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_367), .A2(n_241), .B(n_152), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_405), .B(n_241), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_382), .B(n_241), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_372), .B(n_15), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_384), .Y(n_446) );
NOR4xp25_ASAP7_75t_SL g447 ( .A(n_391), .B(n_20), .C(n_21), .D(n_22), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_367), .B(n_155), .C(n_151), .D(n_27), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_386), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_390), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_380), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_388), .B(n_155), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_397), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_376), .A2(n_230), .B1(n_152), .B2(n_155), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_390), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_368), .Y(n_456) );
O2A1O1Ixp5_ASAP7_75t_L g457 ( .A1(n_370), .A2(n_25), .B(n_26), .C(n_32), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_389), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_405), .B(n_199), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_409), .B(n_151), .C(n_35), .D(n_37), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_389), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_401), .B(n_34), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_450), .B(n_371), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_431), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_437), .B(n_393), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_429), .A2(n_414), .B(n_417), .C(n_371), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_442), .A2(n_416), .B(n_408), .C(n_396), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_455), .B(n_413), .Y(n_468) );
INVxp33_ASAP7_75t_L g469 ( .A(n_449), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_458), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_461), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_446), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_436), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_421), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_448), .A2(n_403), .B1(n_400), .B2(n_396), .Y(n_475) );
INVxp67_ASAP7_75t_L g476 ( .A(n_456), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_428), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_453), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_425), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_425), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_441), .A2(n_403), .B1(n_398), .B2(n_402), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_433), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_434), .A2(n_411), .B(n_369), .C(n_199), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_451), .Y(n_486) );
XNOR2xp5_ASAP7_75t_L g487 ( .A(n_445), .B(n_419), .Y(n_487) );
AOI321xp33_ASAP7_75t_L g488 ( .A1(n_429), .A2(n_411), .A3(n_369), .B1(n_42), .B2(n_49), .C(n_51), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_452), .B(n_38), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_430), .A2(n_40), .B(n_54), .C(n_55), .Y(n_491) );
AOI211x1_ASAP7_75t_SL g492 ( .A1(n_430), .A2(n_58), .B(n_60), .C(n_62), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_477), .Y(n_493) );
AOI211xp5_ASAP7_75t_L g494 ( .A1(n_487), .A2(n_460), .B(n_423), .C(n_444), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_464), .A2(n_438), .B1(n_440), .B2(n_443), .Y(n_495) );
OAI321xp33_ASAP7_75t_L g496 ( .A1(n_488), .A2(n_422), .A3(n_426), .B1(n_420), .B2(n_424), .C(n_454), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_480), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_464), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_476), .A2(n_457), .B(n_439), .Y(n_499) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_491), .B(n_462), .Y(n_500) );
AOI21xp33_ASAP7_75t_SL g501 ( .A1(n_476), .A2(n_459), .B(n_462), .Y(n_501) );
XOR2xp5_ASAP7_75t_L g502 ( .A(n_490), .B(n_422), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_481), .Y(n_503) );
INVxp67_ASAP7_75t_L g504 ( .A(n_489), .Y(n_504) );
XNOR2x1_ASAP7_75t_L g505 ( .A(n_486), .B(n_447), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_468), .Y(n_506) );
AOI211xp5_ASAP7_75t_L g507 ( .A1(n_469), .A2(n_427), .B(n_435), .C(n_199), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_479), .Y(n_508) );
AOI32xp33_ASAP7_75t_L g509 ( .A1(n_465), .A2(n_435), .A3(n_230), .B1(n_66), .B2(n_68), .Y(n_509) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_500), .B(n_466), .Y(n_510) );
AOI21xp33_ASAP7_75t_L g511 ( .A1(n_505), .A2(n_467), .B(n_472), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_496), .A2(n_485), .B(n_475), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_SL g513 ( .A1(n_499), .A2(n_494), .B(n_509), .C(n_495), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_506), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_495), .A2(n_483), .B1(n_473), .B2(n_474), .C(n_471), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_498), .A2(n_483), .B1(n_482), .B2(n_463), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_493), .Y(n_517) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_498), .A2(n_470), .B1(n_478), .B2(n_484), .C(n_492), .Y(n_518) );
OR5x1_ASAP7_75t_L g519 ( .A(n_513), .B(n_510), .C(n_511), .D(n_512), .E(n_515), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_518), .B(n_514), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_517), .Y(n_521) );
NAND3x1_ASAP7_75t_L g522 ( .A(n_516), .B(n_497), .C(n_503), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_515), .B(n_504), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_520), .B(n_501), .C(n_507), .Y(n_524) );
NOR2x1_ASAP7_75t_L g525 ( .A(n_523), .B(n_519), .Y(n_525) );
NOR2x1p5_ASAP7_75t_L g526 ( .A(n_521), .B(n_508), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_526), .B(n_504), .Y(n_527) );
OR3x1_ASAP7_75t_L g528 ( .A(n_525), .B(n_522), .C(n_524), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_527), .Y(n_529) );
AOI21xp33_ASAP7_75t_SL g530 ( .A1(n_529), .A2(n_528), .B(n_502), .Y(n_530) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_530), .A2(n_152), .B1(n_230), .B2(n_199), .C1(n_76), .C2(n_64), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_531), .A2(n_152), .B(n_230), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_532), .A2(n_65), .B(n_71), .Y(n_533) );
endmodule