module fake_jpeg_988_n_477 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_477);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_477;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_94),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_58),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_52),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_96),
.Y(n_129)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_97),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_20),
.B(n_14),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_20),
.B(n_14),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_14),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_31),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_104),
.Y(n_154)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_23),
.B1(n_29),
.B2(n_33),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_108),
.A2(n_139),
.B1(n_23),
.B2(n_21),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_118),
.B(n_144),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_122),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_24),
.B(n_51),
.C(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_135),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_54),
.B(n_39),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_56),
.B(n_39),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_140),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_59),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_60),
.B(n_42),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_61),
.B(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_64),
.B(n_30),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_158),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_58),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_160),
.B1(n_32),
.B2(n_92),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_73),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_78),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_34),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_55),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_166),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_174),
.A2(n_176),
.B1(n_202),
.B2(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_32),
.B1(n_25),
.B2(n_28),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_107),
.A2(n_95),
.B1(n_91),
.B2(n_89),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_179),
.A2(n_209),
.B1(n_210),
.B2(n_119),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_182),
.Y(n_244)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_122),
.A2(n_88),
.B1(n_84),
.B2(n_83),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_208),
.B1(n_119),
.B2(n_110),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_R g189 ( 
.A(n_137),
.B(n_34),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_192),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_45),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_25),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

BUFx4f_ASAP7_75t_SL g197 ( 
.A(n_117),
.Y(n_197)
);

INVx4_ASAP7_75t_SL g198 ( 
.A(n_131),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_199),
.Y(n_243)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_131),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_200),
.B(n_207),
.Y(n_239)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_204),
.Y(n_245)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_113),
.B(n_49),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_206),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_115),
.B(n_42),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_148),
.A2(n_160),
.B1(n_77),
.B2(n_113),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_155),
.A2(n_24),
.B1(n_51),
.B2(n_50),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_37),
.B1(n_38),
.B2(n_48),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_112),
.B(n_49),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_213),
.B(n_143),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_172),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_225),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_38),
.B(n_37),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_217),
.A2(n_234),
.B(n_218),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_249),
.B1(n_243),
.B2(n_225),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_162),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_145),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_249),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_180),
.A2(n_21),
.B(n_48),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_159),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_251),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_212),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_267),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_188),
.B1(n_174),
.B2(n_198),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_255),
.A2(n_259),
.B1(n_278),
.B2(n_281),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_223),
.A2(n_192),
.B1(n_168),
.B2(n_184),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_270),
.B(n_272),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_205),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_268),
.C(n_228),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_176),
.B1(n_127),
.B2(n_151),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

BUFx24_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

INVx4_ASAP7_75t_SL g287 ( 
.A(n_263),
.Y(n_287)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_280),
.B1(n_235),
.B2(n_221),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_178),
.B(n_173),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_227),
.B(n_219),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_217),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_187),
.C(n_213),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_229),
.B(n_189),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_273),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_242),
.A2(n_197),
.B(n_207),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_169),
.B(n_190),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_197),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_194),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_236),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_248),
.A2(n_127),
.B1(n_151),
.B2(n_110),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_235),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_126),
.B1(n_146),
.B2(n_153),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_232),
.A2(n_116),
.B1(n_134),
.B2(n_153),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_290),
.B1(n_307),
.B2(n_278),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_286),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_289),
.B(n_299),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_265),
.A2(n_203),
.B1(n_134),
.B2(n_116),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_267),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_292),
.A2(n_294),
.B(n_296),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_255),
.A2(n_170),
.B1(n_228),
.B2(n_221),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_293),
.A2(n_264),
.B1(n_260),
.B2(n_275),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_254),
.A2(n_227),
.B(n_231),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_247),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_252),
.B(n_247),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_268),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_251),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_302),
.B(n_306),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_214),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_262),
.A2(n_276),
.B(n_256),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_270),
.B(n_272),
.C(n_274),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_276),
.B(n_240),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_257),
.A2(n_269),
.B1(n_259),
.B2(n_280),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_312),
.A2(n_305),
.B1(n_297),
.B2(n_290),
.Y(n_362)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_314),
.A2(n_317),
.B1(n_318),
.B2(n_322),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_321),
.C(n_326),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_258),
.B1(n_266),
.B2(n_273),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_285),
.A2(n_253),
.B1(n_261),
.B2(n_271),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_320),
.B(n_323),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_240),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_284),
.A2(n_271),
.B1(n_281),
.B2(n_261),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_230),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_271),
.B1(n_231),
.B2(n_222),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_324),
.A2(n_305),
.B1(n_302),
.B2(n_298),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_289),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_325),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_220),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_222),
.C(n_214),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_286),
.C(n_283),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_296),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_330),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_300),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_308),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_334),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_336),
.Y(n_338)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_292),
.A2(n_226),
.B1(n_220),
.B2(n_263),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_335),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_295),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_345),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_310),
.A2(n_288),
.B1(n_293),
.B2(n_303),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_341),
.A2(n_362),
.B1(n_322),
.B2(n_342),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_328),
.A2(n_283),
.B(n_294),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_344),
.A2(n_310),
.B(n_312),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_315),
.B(n_295),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_359),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_309),
.C(n_299),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_358),
.C(n_360),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_230),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_351),
.B(n_353),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_363),
.B1(n_336),
.B2(n_125),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_330),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_328),
.A2(n_286),
.B(n_293),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_324),
.B(n_319),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_298),
.C(n_297),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_317),
.B(n_288),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_316),
.C(n_329),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_314),
.A2(n_291),
.B1(n_287),
.B2(n_244),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_356),
.Y(n_364)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_366),
.A2(n_367),
.B(n_263),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_349),
.Y(n_369)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_369),
.Y(n_392)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_346),
.Y(n_371)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_311),
.C(n_334),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_377),
.C(n_379),
.Y(n_395)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_374),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_375),
.A2(n_380),
.B1(n_341),
.B2(n_363),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_332),
.C(n_313),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_226),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_345),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_291),
.C(n_185),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_361),
.A2(n_355),
.B1(n_357),
.B2(n_349),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_338),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_383),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_186),
.C(n_287),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_350),
.C(n_130),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_287),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_358),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_263),
.Y(n_406)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_387),
.A2(n_142),
.B1(n_128),
.B2(n_125),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_244),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_146),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_389),
.A2(n_391),
.B1(n_408),
.B2(n_387),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_407),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_364),
.A2(n_362),
.B1(n_359),
.B2(n_350),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_370),
.B(n_344),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_376),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_397),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_406),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_404),
.Y(n_422)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_126),
.C(n_263),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_163),
.B1(n_142),
.B2(n_128),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_401),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_373),
.B1(n_367),
.B2(n_366),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_414),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_395),
.B(n_377),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_385),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_417),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_365),
.C(n_370),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_419),
.C(n_402),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_393),
.B(n_376),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_392),
.A2(n_369),
.B(n_380),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_418),
.A2(n_396),
.B(n_399),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_365),
.C(n_379),
.Y(n_419)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_420),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_394),
.Y(n_423)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_423),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_382),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_403),
.Y(n_437)
);

XOR2x1_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_394),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_427),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_426),
.B(n_429),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_397),
.C(n_388),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_383),
.C(n_399),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_436),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_433),
.A2(n_435),
.B(n_422),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_418),
.A2(n_405),
.B(n_384),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_400),
.C(n_374),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_438),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_404),
.C(n_182),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_413),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_428),
.A2(n_421),
.B1(n_422),
.B2(n_417),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_442),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_441),
.A2(n_166),
.B(n_13),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_427),
.C(n_431),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_443),
.B(n_451),
.Y(n_455)
);

NOR2x1_ASAP7_75t_R g447 ( 
.A(n_432),
.B(n_411),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_447),
.A2(n_2),
.B(n_3),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_449),
.B(n_450),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_434),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_413),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_428),
.A2(n_424),
.B1(n_163),
.B2(n_166),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_13),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_453),
.A2(n_456),
.B(n_458),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_457),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_444),
.A2(n_47),
.B(n_40),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_0),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_450),
.A2(n_47),
.B(n_40),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_447),
.C(n_449),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_445),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_462),
.A2(n_464),
.B(n_466),
.Y(n_468)
);

AO21x1_ASAP7_75t_L g464 ( 
.A1(n_459),
.A2(n_446),
.B(n_448),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_52),
.C(n_5),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_461),
.B(n_3),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_467),
.A2(n_461),
.B(n_47),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_469),
.B(n_470),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_463),
.A2(n_52),
.B(n_5),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_3),
.C(n_6),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_472),
.B(n_468),
.C(n_6),
.Y(n_474)
);

OAI321xp33_ASAP7_75t_L g475 ( 
.A1(n_474),
.A2(n_473),
.A3(n_8),
.B1(n_11),
.B2(n_12),
.C(n_3),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_8),
.C(n_12),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_476),
.A2(n_8),
.B(n_12),
.Y(n_477)
);


endmodule