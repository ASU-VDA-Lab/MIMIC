module real_jpeg_13686_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_41),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_45),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_45),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_20),
.B(n_21),
.C(n_26),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_10),
.B(n_73),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_10),
.B(n_34),
.C(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_10),
.B(n_59),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_10),
.A2(n_79),
.B(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_52),
.Y(n_110)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_93),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_63),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_17),
.B(n_63),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_42),
.C(n_54),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_18),
.B(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_29),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_29),
.Y(n_84)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_20),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_58)
);

AO22x1_ASAP7_75t_SL g59 ( 
.A1(n_20),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_24),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_23),
.B(n_50),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_23),
.B(n_30),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_25),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_25),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_26),
.A2(n_27),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B(n_38),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_30),
.A2(n_32),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_30),
.A2(n_38),
.B(n_116),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_31),
.B(n_40),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_31),
.A2(n_39),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_33),
.B(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_42),
.A2(n_54),
.B1(n_55),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_42),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_44),
.A2(n_50),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_46),
.B(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_82),
.B2(n_83),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_77),
.B2(n_78),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_88),
.B(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_131),
.B(n_136),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_112),
.B(n_130),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_100),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_107),
.C(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_120),
.B(n_129),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_114),
.B(n_118),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_124),
.B(n_128),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);


endmodule