module real_aes_9844_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_0), .A2(n_188), .B1(n_704), .B2(n_706), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_0), .A2(n_3), .B1(n_454), .B2(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1), .Y(n_1109) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_2), .A2(n_66), .B1(n_751), .B2(n_910), .Y(n_916) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_2), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_3), .A2(n_152), .B1(n_645), .B2(n_701), .C(n_702), .Y(n_700) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_4), .Y(n_247) );
AND2x2_ASAP7_75t_L g267 ( .A(n_4), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g300 ( .A(n_4), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_4), .B(n_176), .Y(n_309) );
INVxp67_ASAP7_75t_L g848 ( .A(n_5), .Y(n_848) );
OAI222xp33_ASAP7_75t_L g863 ( .A1(n_5), .A2(n_36), .B1(n_225), .B2(n_864), .C1(n_865), .C2(n_867), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_6), .A2(n_313), .B1(n_315), .B2(n_323), .C(n_334), .Y(n_312) );
INVx1_ASAP7_75t_L g404 ( .A(n_6), .Y(n_404) );
XNOR2x2_ASAP7_75t_L g609 ( .A(n_7), .B(n_610), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_8), .A2(n_154), .B1(n_521), .B2(n_565), .C(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g590 ( .A(n_8), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_9), .A2(n_47), .B1(n_292), .B2(n_295), .C(n_296), .Y(n_291) );
INVx1_ASAP7_75t_L g425 ( .A(n_9), .Y(n_425) );
INVx1_ASAP7_75t_L g274 ( .A(n_10), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_10), .A2(n_49), .B1(n_396), .B2(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g1221 ( .A(n_11), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_12), .A2(n_75), .B1(n_575), .B2(n_1321), .Y(n_1320) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_12), .A2(n_27), .B1(n_266), .B2(n_307), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_13), .A2(n_215), .B1(n_575), .B2(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g600 ( .A(n_13), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_14), .A2(n_32), .B1(n_521), .B2(n_691), .Y(n_690) );
INVxp33_ASAP7_75t_SL g735 ( .A(n_14), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_15), .A2(n_223), .B1(n_772), .B2(n_880), .C(n_881), .Y(n_948) );
INVx1_ASAP7_75t_L g968 ( .A(n_15), .Y(n_968) );
AO221x2_ASAP7_75t_L g1130 ( .A1(n_16), .A2(n_52), .B1(n_1107), .B2(n_1129), .C(n_1131), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_17), .Y(n_328) );
INVx1_ASAP7_75t_L g1148 ( .A(n_18), .Y(n_1148) );
AOI221xp5_ASAP7_75t_L g1345 ( .A1(n_19), .A2(n_127), .B1(n_296), .B2(n_1346), .C(n_1347), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_19), .A2(n_198), .B1(n_429), .B2(n_675), .Y(n_1354) );
INVx2_ASAP7_75t_L g350 ( .A(n_20), .Y(n_350) );
OR2x2_ASAP7_75t_L g420 ( .A(n_20), .B(n_348), .Y(n_420) );
AO22x1_ASAP7_75t_L g259 ( .A1(n_21), .A2(n_260), .B1(n_431), .B2(n_432), .Y(n_259) );
INVx1_ASAP7_75t_L g432 ( .A(n_21), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g1011 ( .A1(n_22), .A2(n_168), .B1(n_287), .B2(n_617), .C(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1019 ( .A(n_22), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_23), .A2(n_210), .B1(n_517), .B2(n_786), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g801 ( .A1(n_23), .A2(n_210), .B1(n_456), .B2(n_461), .C(n_802), .Y(n_801) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_24), .A2(n_91), .B1(n_456), .B2(n_461), .C(n_464), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_24), .A2(n_91), .B1(n_514), .B2(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g851 ( .A(n_25), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_26), .A2(n_58), .B1(n_1317), .B2(n_1318), .Y(n_1316) );
INVx1_ASAP7_75t_L g1342 ( .A(n_26), .Y(n_1342) );
OAI222xp33_ASAP7_75t_L g1353 ( .A1(n_27), .A2(n_127), .B1(n_131), .B2(n_554), .C1(n_1088), .C2(n_1089), .Y(n_1353) );
BUFx2_ASAP7_75t_L g339 ( .A(n_28), .Y(n_339) );
BUFx2_ASAP7_75t_L g344 ( .A(n_28), .Y(n_344) );
INVx1_ASAP7_75t_L g372 ( .A(n_28), .Y(n_372) );
OR2x2_ASAP7_75t_L g460 ( .A(n_28), .B(n_309), .Y(n_460) );
INVx1_ASAP7_75t_L g1219 ( .A(n_29), .Y(n_1219) );
INVx1_ASAP7_75t_L g995 ( .A(n_30), .Y(n_995) );
INVx1_ASAP7_75t_L g1042 ( .A(n_31), .Y(n_1042) );
INVxp33_ASAP7_75t_SL g730 ( .A(n_32), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g909 ( .A1(n_33), .A2(n_164), .B1(n_751), .B2(n_910), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g933 ( .A1(n_33), .A2(n_220), .B1(n_655), .B2(n_934), .C(n_935), .Y(n_933) );
INVx1_ASAP7_75t_L g837 ( .A(n_34), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g1365 ( .A1(n_35), .A2(n_1312), .B1(n_1366), .B2(n_1367), .Y(n_1365) );
CKINVDCx5p33_ASAP7_75t_R g1366 ( .A(n_35), .Y(n_1366) );
INVxp67_ASAP7_75t_L g846 ( .A(n_36), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_37), .A2(n_180), .B1(n_575), .B2(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g807 ( .A(n_37), .Y(n_807) );
CKINVDCx16_ASAP7_75t_R g1145 ( .A(n_38), .Y(n_1145) );
INVx1_ASAP7_75t_L g322 ( .A(n_39), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_39), .A2(n_123), .B1(n_394), .B2(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g1215 ( .A(n_40), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_41), .A2(n_132), .B1(n_302), .B2(n_310), .Y(n_301) );
OAI22xp5_ASAP7_75t_SL g364 ( .A1(n_41), .A2(n_132), .B1(n_365), .B2(n_373), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_42), .A2(n_45), .B1(n_615), .B2(n_617), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_42), .A2(n_59), .B1(n_429), .B2(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g1003 ( .A(n_43), .Y(n_1003) );
INVx1_ASAP7_75t_L g1330 ( .A(n_44), .Y(n_1330) );
OAI221xp5_ASAP7_75t_L g1349 ( .A1(n_44), .A2(n_76), .B1(n_302), .B2(n_310), .C(n_1350), .Y(n_1349) );
INVxp67_ASAP7_75t_SL g672 ( .A(n_45), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_46), .A2(n_81), .B1(n_912), .B2(n_913), .Y(n_915) );
INVxp33_ASAP7_75t_SL g942 ( .A(n_46), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_47), .A2(n_96), .B1(n_427), .B2(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g635 ( .A(n_48), .Y(n_635) );
INVx1_ASAP7_75t_L g280 ( .A(n_49), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_50), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_51), .A2(n_173), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
INVxp67_ASAP7_75t_SL g1079 ( .A(n_51), .Y(n_1079) );
INVx1_ASAP7_75t_L g498 ( .A(n_53), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g1084 ( .A(n_54), .Y(n_1084) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_55), .A2(n_61), .B1(n_572), .B2(n_772), .C(n_774), .Y(n_771) );
INVxp67_ASAP7_75t_SL g810 ( .A(n_55), .Y(n_810) );
INVx1_ASAP7_75t_L g1157 ( .A(n_56), .Y(n_1157) );
CKINVDCx16_ASAP7_75t_R g1162 ( .A(n_57), .Y(n_1162) );
INVx1_ASAP7_75t_L g1340 ( .A(n_58), .Y(n_1340) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_59), .A2(n_166), .B1(n_296), .B2(n_620), .C(n_622), .Y(n_619) );
INVxp33_ASAP7_75t_SL g475 ( .A(n_60), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_60), .A2(n_86), .B1(n_530), .B2(n_531), .C(n_533), .Y(n_529) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_61), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g998 ( .A1(n_62), .A2(n_114), .B1(n_485), .B2(n_999), .C(n_1000), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_62), .A2(n_79), .B1(n_536), .B2(n_539), .Y(n_1022) );
INVxp33_ASAP7_75t_SL g715 ( .A(n_63), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g750 ( .A1(n_63), .A2(n_101), .B1(n_743), .B2(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g1115 ( .A(n_64), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_65), .A2(n_207), .B1(n_521), .B2(n_662), .Y(n_949) );
INVx1_ASAP7_75t_L g969 ( .A(n_65), .Y(n_969) );
INVxp33_ASAP7_75t_L g941 ( .A(n_66), .Y(n_941) );
INVx1_ASAP7_75t_L g1002 ( .A(n_67), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1021 ( .A1(n_67), .A2(n_114), .B1(n_520), .B2(n_531), .C(n_533), .Y(n_1021) );
INVxp33_ASAP7_75t_L g442 ( .A(n_68), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_68), .A2(n_233), .B1(n_520), .B2(n_521), .C(n_522), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_69), .A2(n_124), .B1(n_878), .B2(n_880), .C(n_881), .Y(n_877) );
OAI221xp5_ASAP7_75t_L g885 ( .A1(n_69), .A2(n_136), .B1(n_886), .B2(n_887), .C(n_889), .Y(n_885) );
CKINVDCx16_ASAP7_75t_R g1164 ( .A(n_70), .Y(n_1164) );
AOI22xp5_ASAP7_75t_L g1122 ( .A1(n_71), .A2(n_119), .B1(n_1123), .B2(n_1126), .Y(n_1122) );
INVx1_ASAP7_75t_L g348 ( .A(n_72), .Y(n_348) );
INVx1_ASAP7_75t_L g381 ( .A(n_72), .Y(n_381) );
INVxp33_ASAP7_75t_L g716 ( .A(n_73), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_73), .A2(n_184), .B1(n_454), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g766 ( .A(n_74), .Y(n_766) );
INVx1_ASAP7_75t_L g1348 ( .A(n_75), .Y(n_1348) );
INVx1_ASAP7_75t_L g1328 ( .A(n_76), .Y(n_1328) );
INVx1_ASAP7_75t_L g1013 ( .A(n_77), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_77), .A2(n_168), .B1(n_540), .B2(n_865), .C(n_1018), .Y(n_1017) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_78), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g922 ( .A1(n_78), .A2(n_192), .B1(n_923), .B2(n_924), .Y(n_922) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_79), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_80), .A2(n_115), .B1(n_521), .B2(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_80), .A2(n_115), .B1(n_1081), .B2(n_1082), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g921 ( .A(n_81), .Y(n_921) );
INVx1_ASAP7_75t_L g1008 ( .A(n_82), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1024 ( .A1(n_82), .A2(n_120), .B1(n_649), .B2(n_1025), .C(n_1026), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_83), .A2(n_217), .B1(n_695), .B2(n_697), .Y(n_694) );
INVxp67_ASAP7_75t_SL g722 ( .A(n_83), .Y(n_722) );
INVx1_ASAP7_75t_L g637 ( .A(n_84), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_84), .A2(n_227), .B1(n_645), .B2(n_648), .C(n_650), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g827 ( .A(n_85), .B(n_828), .Y(n_827) );
INVxp67_ASAP7_75t_SL g479 ( .A(n_86), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_87), .Y(n_959) );
INVxp67_ASAP7_75t_L g835 ( .A(n_88), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g869 ( .A1(n_88), .A2(n_139), .B1(n_572), .B2(n_774), .C(n_870), .Y(n_869) );
OAI21xp33_ASAP7_75t_L g991 ( .A1(n_89), .A2(n_992), .B(n_1015), .Y(n_991) );
INVx1_ASAP7_75t_L g1031 ( .A(n_89), .Y(n_1031) );
INVx1_ASAP7_75t_L g1147 ( .A(n_89), .Y(n_1147) );
AOI22xp33_ASAP7_75t_SL g1319 ( .A1(n_90), .A2(n_135), .B1(n_657), .B2(n_880), .Y(n_1319) );
AOI21xp33_ASAP7_75t_L g1338 ( .A1(n_90), .A2(n_361), .B(n_468), .Y(n_1338) );
INVx1_ASAP7_75t_L g1014 ( .A(n_92), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_93), .A2(n_194), .B1(n_530), .B2(n_772), .C(n_937), .Y(n_954) );
INVx1_ASAP7_75t_L g978 ( .A(n_93), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_94), .A2(n_202), .B1(n_783), .B2(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g799 ( .A(n_94), .Y(n_799) );
AO221x2_ASAP7_75t_L g1100 ( .A1(n_95), .A2(n_158), .B1(n_1101), .B2(n_1107), .C(n_1108), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_96), .A2(n_107), .B1(n_287), .B2(n_288), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_97), .A2(n_187), .B1(n_423), .B2(n_772), .C(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g798 ( .A(n_97), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_98), .A2(n_211), .B1(n_373), .B2(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1071 ( .A(n_98), .Y(n_1071) );
INVx1_ASAP7_75t_L g239 ( .A(n_99), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_100), .Y(n_581) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_101), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g961 ( .A(n_102), .Y(n_961) );
XOR2x2_ASAP7_75t_L g1033 ( .A(n_103), .B(n_1034), .Y(n_1033) );
OA22x2_ASAP7_75t_L g943 ( .A1(n_104), .A2(n_944), .B1(n_985), .B2(n_986), .Y(n_943) );
INVx1_ASAP7_75t_L g986 ( .A(n_104), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_105), .Y(n_681) );
INVx1_ASAP7_75t_L g1049 ( .A(n_106), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1073 ( .A1(n_106), .A2(n_313), .B1(n_639), .B2(n_1074), .C(n_1076), .Y(n_1073) );
INVx1_ASAP7_75t_L g421 ( .A(n_107), .Y(n_421) );
OAI221xp5_ASAP7_75t_SL g1006 ( .A1(n_108), .A2(n_208), .B1(n_489), .B2(n_634), .C(n_1007), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_108), .A2(n_208), .B1(n_394), .B2(n_708), .Y(n_1027) );
AOI22xp5_ASAP7_75t_L g1128 ( .A1(n_109), .A2(n_151), .B1(n_1107), .B2(n_1129), .Y(n_1128) );
AOI221xp5_ASAP7_75t_L g1064 ( .A1(n_110), .A2(n_170), .B1(n_1065), .B2(n_1066), .C(n_1067), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_110), .A2(n_147), .B1(n_429), .B2(n_675), .Y(n_1086) );
INVx1_ASAP7_75t_L g503 ( .A(n_111), .Y(n_503) );
INVx1_ASAP7_75t_L g642 ( .A(n_112), .Y(n_642) );
OAI222xp33_ASAP7_75t_L g830 ( .A1(n_113), .A2(n_138), .B1(n_228), .B2(n_553), .C1(n_831), .C2(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g858 ( .A(n_113), .Y(n_858) );
INVx1_ASAP7_75t_L g1132 ( .A(n_116), .Y(n_1132) );
INVx1_ASAP7_75t_L g1061 ( .A(n_117), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_117), .A2(n_170), .B1(n_1088), .B2(n_1089), .Y(n_1087) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_118), .Y(n_960) );
XNOR2xp5_ASAP7_75t_L g1311 ( .A(n_119), .B(n_1312), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_119), .A2(n_1360), .B1(n_1364), .B2(n_1368), .Y(n_1359) );
INVx1_ASAP7_75t_L g1009 ( .A(n_120), .Y(n_1009) );
INVx1_ASAP7_75t_L g491 ( .A(n_121), .Y(n_491) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_122), .A2(n_229), .B1(n_533), .B2(n_572), .C(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g599 ( .A(n_122), .Y(n_599) );
INVx1_ASAP7_75t_L g319 ( .A(n_123), .Y(n_319) );
OAI332xp33_ASAP7_75t_L g833 ( .A1(n_124), .A2(n_467), .A3(n_821), .B1(n_834), .B2(n_838), .B3(n_841), .C1(n_847), .C2(n_852), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_125), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_126), .A2(n_146), .B1(n_302), .B2(n_310), .Y(n_625) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_126), .A2(n_146), .B1(n_667), .B2(n_669), .C(n_670), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g918 ( .A(n_128), .Y(n_918) );
INVx1_ASAP7_75t_L g770 ( .A(n_129), .Y(n_770) );
XNOR2xp5_ASAP7_75t_L g556 ( .A(n_130), .B(n_557), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g1135 ( .A1(n_130), .A2(n_143), .B1(n_1123), .B2(n_1126), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_131), .A2(n_198), .B1(n_288), .B2(n_999), .Y(n_1344) );
AOI22xp33_ASAP7_75t_SL g1322 ( .A1(n_133), .A2(n_148), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
INVx1_ASAP7_75t_L g1333 ( .A(n_133), .Y(n_1333) );
XOR2x2_ASAP7_75t_L g893 ( .A(n_134), .B(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g1337 ( .A(n_135), .Y(n_1337) );
INVx1_ASAP7_75t_L g876 ( .A(n_136), .Y(n_876) );
INVxp33_ASAP7_75t_L g471 ( .A(n_137), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_137), .A2(n_172), .B1(n_536), .B2(n_539), .Y(n_535) );
INVx1_ASAP7_75t_L g874 ( .A(n_138), .Y(n_874) );
INVx1_ASAP7_75t_L g839 ( .A(n_139), .Y(n_839) );
INVx1_ASAP7_75t_L g550 ( .A(n_140), .Y(n_550) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_141), .Y(n_241) );
AND3x2_ASAP7_75t_L g1105 ( .A(n_141), .B(n_239), .C(n_1106), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_141), .B(n_239), .Y(n_1112) );
OAI22xp33_ASAP7_75t_SL g562 ( .A1(n_142), .A2(n_161), .B1(n_514), .B2(n_563), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_142), .A2(n_161), .B1(n_456), .B2(n_461), .C(n_464), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g1136 ( .A1(n_144), .A2(n_182), .B1(n_1101), .B2(n_1137), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_145), .A2(n_214), .B1(n_685), .B2(n_687), .C(n_688), .Y(n_684) );
INVxp33_ASAP7_75t_SL g732 ( .A(n_145), .Y(n_732) );
INVx1_ASAP7_75t_L g1063 ( .A(n_147), .Y(n_1063) );
INVx1_ASAP7_75t_L g1334 ( .A(n_148), .Y(n_1334) );
INVx2_ASAP7_75t_L g252 ( .A(n_149), .Y(n_252) );
INVx1_ASAP7_75t_L g788 ( .A(n_150), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_152), .A2(n_188), .B1(n_741), .B2(n_743), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_153), .A2(n_216), .B1(n_880), .B2(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g975 ( .A(n_153), .Y(n_975) );
INVx1_ASAP7_75t_L g587 ( .A(n_154), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_155), .Y(n_957) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_156), .Y(n_906) );
OAI211xp5_ASAP7_75t_L g262 ( .A1(n_157), .A2(n_263), .B(n_273), .C(n_285), .Y(n_262) );
INVx1_ASAP7_75t_L g405 ( .A(n_157), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_159), .A2(n_167), .B1(n_1107), .B2(n_1129), .Y(n_1174) );
INVx1_ASAP7_75t_L g994 ( .A(n_160), .Y(n_994) );
INVxp33_ASAP7_75t_SL g907 ( .A(n_162), .Y(n_907) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_162), .A2(n_201), .B1(n_926), .B2(n_928), .C(n_929), .Y(n_925) );
INVx1_ASAP7_75t_L g633 ( .A(n_163), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_164), .A2(n_186), .B1(n_708), .B2(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g1106 ( .A(n_165), .Y(n_1106) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_166), .Y(n_673) );
CKINVDCx16_ASAP7_75t_R g1143 ( .A(n_169), .Y(n_1143) );
INVx1_ASAP7_75t_L g1217 ( .A(n_171), .Y(n_1217) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_172), .Y(n_483) );
INVxp67_ASAP7_75t_SL g1077 ( .A(n_173), .Y(n_1077) );
OAI211xp5_ASAP7_75t_L g612 ( .A1(n_174), .A2(n_263), .B(n_613), .C(n_626), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_174), .A2(n_178), .B1(n_655), .B2(n_658), .C(n_659), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_175), .Y(n_677) );
INVx1_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
INVx2_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
INVx1_ASAP7_75t_L g627 ( .A(n_177), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_178), .A2(n_313), .B1(n_630), .B2(n_636), .C(n_639), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g1173 ( .A1(n_179), .A2(n_212), .B1(n_1123), .B2(n_1126), .Y(n_1173) );
INVx1_ASAP7_75t_L g815 ( .A(n_180), .Y(n_815) );
INVx1_ASAP7_75t_L g341 ( .A(n_181), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_183), .A2(n_761), .B1(n_822), .B2(n_823), .Y(n_760) );
INVx1_ASAP7_75t_L g823 ( .A(n_183), .Y(n_823) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_184), .Y(n_693) );
INVx1_ASAP7_75t_L g496 ( .A(n_185), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_186), .A2(n_220), .B1(n_912), .B2(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g795 ( .A(n_187), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_189), .Y(n_570) );
INVx1_ASAP7_75t_L g449 ( .A(n_190), .Y(n_449) );
INVx1_ASAP7_75t_L g1039 ( .A(n_191), .Y(n_1039) );
INVxp67_ASAP7_75t_SL g901 ( .A(n_192), .Y(n_901) );
INVx1_ASAP7_75t_L g437 ( .A(n_193), .Y(n_437) );
INVx1_ASAP7_75t_L g976 ( .A(n_194), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_195), .Y(n_950) );
INVx1_ASAP7_75t_L g904 ( .A(n_196), .Y(n_904) );
CKINVDCx5p33_ASAP7_75t_R g582 ( .A(n_197), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_199), .A2(n_205), .B1(n_517), .B2(n_952), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g970 ( .A1(n_199), .A2(n_205), .B1(n_461), .B2(n_802), .C(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g1158 ( .A(n_200), .Y(n_1158) );
INVxp33_ASAP7_75t_SL g903 ( .A(n_201), .Y(n_903) );
INVx1_ASAP7_75t_L g793 ( .A(n_202), .Y(n_793) );
INVx1_ASAP7_75t_L g1104 ( .A(n_203), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_203), .B(n_1114), .Y(n_1117) );
INVx1_ASAP7_75t_L g860 ( .A(n_204), .Y(n_860) );
INVx1_ASAP7_75t_L g779 ( .A(n_206), .Y(n_779) );
INVx1_ASAP7_75t_L g965 ( .A(n_207), .Y(n_965) );
INVx1_ASAP7_75t_L g840 ( .A(n_209), .Y(n_840) );
INVx1_ASAP7_75t_L g1069 ( .A(n_211), .Y(n_1069) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_213), .Y(n_567) );
INVxp33_ASAP7_75t_L g734 ( .A(n_214), .Y(n_734) );
INVx1_ASAP7_75t_L g595 ( .A(n_215), .Y(n_595) );
INVx1_ASAP7_75t_L g980 ( .A(n_216), .Y(n_980) );
INVxp67_ASAP7_75t_SL g726 ( .A(n_217), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_218), .Y(n_331) );
INVx2_ASAP7_75t_L g251 ( .A(n_219), .Y(n_251) );
INVx1_ASAP7_75t_L g1051 ( .A(n_221), .Y(n_1051) );
OAI211xp5_ASAP7_75t_SL g1058 ( .A1(n_221), .A2(n_263), .B(n_1059), .C(n_1068), .Y(n_1058) );
INVx1_ASAP7_75t_L g628 ( .A(n_222), .Y(n_628) );
INVx1_ASAP7_75t_L g966 ( .A(n_223), .Y(n_966) );
INVx1_ASAP7_75t_L g446 ( .A(n_224), .Y(n_446) );
INVxp67_ASAP7_75t_L g842 ( .A(n_225), .Y(n_842) );
INVx1_ASAP7_75t_L g583 ( .A(n_226), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g638 ( .A1(n_227), .A2(n_468), .B(n_620), .Y(n_638) );
INVx1_ASAP7_75t_L g861 ( .A(n_228), .Y(n_861) );
INVx1_ASAP7_75t_L g596 ( .A(n_229), .Y(n_596) );
BUFx3_ASAP7_75t_L g353 ( .A(n_230), .Y(n_353) );
INVx1_ASAP7_75t_L g387 ( .A(n_230), .Y(n_387) );
BUFx3_ASAP7_75t_L g355 ( .A(n_231), .Y(n_355) );
INVx1_ASAP7_75t_L g389 ( .A(n_231), .Y(n_389) );
INVx1_ASAP7_75t_L g765 ( .A(n_232), .Y(n_765) );
INVxp33_ASAP7_75t_L g452 ( .A(n_233), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_255), .B(n_1092), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_242), .Y(n_236) );
AND2x4_ASAP7_75t_L g1358 ( .A(n_237), .B(n_243), .Y(n_1358) );
NOR2xp33_ASAP7_75t_SL g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx1_ASAP7_75t_SL g1363 ( .A(n_238), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_238), .B(n_240), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_240), .B(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g333 ( .A(n_246), .B(n_254), .Y(n_333) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g468 ( .A(n_247), .B(n_469), .Y(n_468) );
OR2x6_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
INVx2_ASAP7_75t_SL g330 ( .A(n_249), .Y(n_330) );
BUFx2_ASAP7_75t_L g474 ( .A(n_249), .Y(n_474) );
OR2x2_ASAP7_75t_L g553 ( .A(n_249), .B(n_460), .Y(n_553) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_249), .Y(n_606) );
INVx2_ASAP7_75t_SL g806 ( .A(n_249), .Y(n_806) );
INVx1_ASAP7_75t_L g850 ( .A(n_249), .Y(n_850) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_249), .A2(n_501), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
OAI22xp33_ASAP7_75t_L g1012 ( .A1(n_249), .A2(n_501), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g271 ( .A(n_251), .Y(n_271) );
INVx2_ASAP7_75t_L g277 ( .A(n_251), .Y(n_277) );
AND2x4_ASAP7_75t_L g284 ( .A(n_251), .B(n_272), .Y(n_284) );
AND2x2_ASAP7_75t_L g294 ( .A(n_251), .B(n_252), .Y(n_294) );
INVx1_ASAP7_75t_L g327 ( .A(n_251), .Y(n_327) );
INVx2_ASAP7_75t_L g272 ( .A(n_252), .Y(n_272) );
INVx1_ASAP7_75t_L g279 ( .A(n_252), .Y(n_279) );
INVx1_ASAP7_75t_L g305 ( .A(n_252), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_252), .B(n_277), .Y(n_318) );
INVx1_ASAP7_75t_L g326 ( .A(n_252), .Y(n_326) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_755), .B1(n_756), .B2(n_1091), .Y(n_255) );
INVx1_ASAP7_75t_L g1091 ( .A(n_256), .Y(n_1091) );
XNOR2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_433), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g431 ( .A(n_260), .Y(n_431) );
NAND4xp25_ASAP7_75t_L g260 ( .A(n_261), .B(n_340), .C(n_363), .D(n_414), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_312), .B(n_336), .Y(n_261) );
INVx8_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI221xp5_ASAP7_75t_SL g1343 ( .A1(n_264), .A2(n_1344), .B1(n_1345), .B2(n_1348), .C(n_1349), .Y(n_1343) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
AND2x4_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g275 ( .A(n_267), .B(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g314 ( .A(n_267), .B(n_293), .Y(n_314) );
AND2x4_ASAP7_75t_L g445 ( .A(n_267), .B(n_372), .Y(n_445) );
INVx1_ASAP7_75t_L g299 ( .A(n_268), .Y(n_299) );
INVx1_ASAP7_75t_L g469 ( .A(n_268), .Y(n_469) );
BUFx6f_ASAP7_75t_L g1347 ( .A(n_269), .Y(n_1347) );
BUFx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx3_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_270), .Y(n_624) );
BUFx2_ASAP7_75t_L g728 ( .A(n_270), .Y(n_728) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_270), .Y(n_745) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_275), .B1(n_280), .B2(n_281), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_275), .A2(n_281), .B1(n_627), .B2(n_628), .Y(n_626) );
INVx3_ASAP7_75t_L g1081 ( .A(n_275), .Y(n_1081) );
AOI221x1_ASAP7_75t_L g1332 ( .A1(n_275), .A2(n_281), .B1(n_1333), .B2(n_1334), .C(n_1335), .Y(n_1332) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_276), .Y(n_287) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_276), .Y(n_454) );
INVx1_ASAP7_75t_L g616 ( .A(n_276), .Y(n_616) );
BUFx6f_ASAP7_75t_L g999 ( .A(n_276), .Y(n_999) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g311 ( .A(n_277), .Y(n_311) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g1082 ( .A(n_281), .Y(n_1082) );
INVx1_ASAP7_75t_L g1341 ( .A(n_282), .Y(n_1341) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g818 ( .A(n_283), .Y(n_818) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g290 ( .A(n_284), .Y(n_290) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_284), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_291), .B(n_301), .Y(n_285) );
BUFx3_ASAP7_75t_L g912 ( .A(n_287), .Y(n_912) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g485 ( .A(n_289), .Y(n_485) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx3_ASAP7_75t_L g321 ( .A(n_290), .Y(n_321) );
INVx3_ASAP7_75t_L g495 ( .A(n_290), .Y(n_495) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g742 ( .A(n_293), .Y(n_742) );
BUFx2_ASAP7_75t_L g1346 ( .A(n_293), .Y(n_1346) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g362 ( .A(n_294), .Y(n_362) );
AND2x6_ASAP7_75t_L g447 ( .A(n_295), .B(n_445), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g465 ( .A(n_295), .B(n_459), .Y(n_465) );
INVx2_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_297), .B(n_358), .Y(n_1010) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x6_ASAP7_75t_L g506 ( .A(n_298), .B(n_371), .Y(n_506) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_298), .Y(n_1067) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NAND2x1_ASAP7_75t_SL g458 ( .A(n_303), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_305), .Y(n_721) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x6_ASAP7_75t_L g310 ( .A(n_307), .B(n_311), .Y(n_310) );
OR2x6_ASAP7_75t_L g334 ( .A(n_307), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
OR2x2_ASAP7_75t_L g639 ( .A(n_307), .B(n_335), .Y(n_639) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
CKINVDCx11_ASAP7_75t_R g1072 ( .A(n_310), .Y(n_1072) );
INVx1_ASAP7_75t_L g463 ( .A(n_311), .Y(n_463) );
CKINVDCx6p67_ASAP7_75t_R g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B1(n_320), .B2(n_322), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g844 ( .A(n_317), .Y(n_844) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g482 ( .A(n_318), .Y(n_482) );
INVx1_ASAP7_75t_L g490 ( .A(n_318), .Y(n_490) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g444 ( .A(n_321), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g634 ( .A(n_321), .Y(n_634) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_328), .B1(n_329), .B2(n_331), .C(n_332), .Y(n_323) );
OAI21xp5_ASAP7_75t_SL g1336 ( .A1(n_324), .A2(n_1337), .B(n_1338), .Y(n_1336) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g335 ( .A(n_325), .Y(n_335) );
BUFx2_ASAP7_75t_L g477 ( .A(n_325), .Y(n_477) );
INVx2_ASAP7_75t_L g607 ( .A(n_325), .Y(n_607) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_326), .B(n_327), .Y(n_502) );
INVx1_ASAP7_75t_L g725 ( .A(n_327), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_328), .A2(n_331), .B1(n_383), .B2(n_390), .C(n_393), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_329), .A2(n_335), .B1(n_839), .B2(n_840), .Y(n_838) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_332), .A2(n_805), .B1(n_1039), .B2(n_1042), .C(n_1075), .Y(n_1074) );
BUFx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g739 ( .A(n_333), .B(n_358), .Y(n_739) );
AND2x4_ASAP7_75t_L g997 ( .A(n_333), .B(n_358), .Y(n_997) );
OAI21xp5_ASAP7_75t_L g1335 ( .A1(n_334), .A2(n_1336), .B(n_1339), .Y(n_1335) );
INVx1_ASAP7_75t_L g809 ( .A(n_335), .Y(n_809) );
BUFx8_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g508 ( .A(n_337), .Y(n_508) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g884 ( .A(n_338), .Y(n_884) );
BUFx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g358 ( .A(n_339), .Y(n_358) );
OR2x6_ASAP7_75t_L g467 ( .A(n_339), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_342), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_342), .B(n_1084), .Y(n_1083) );
OR2x6_ASAP7_75t_L g342 ( .A(n_343), .B(n_356), .Y(n_342) );
INVx2_ASAP7_75t_L g554 ( .A(n_343), .Y(n_554) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x4_ASAP7_75t_L g399 ( .A(n_344), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g1325 ( .A(n_344), .B(n_400), .Y(n_1325) );
INVx2_ASAP7_75t_L g857 ( .A(n_345), .Y(n_857) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_351), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_346), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g515 ( .A(n_346), .B(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g518 ( .A(n_346), .B(n_375), .Y(n_518) );
BUFx2_ASAP7_75t_L g543 ( .A(n_346), .Y(n_543) );
AND2x4_ASAP7_75t_L g696 ( .A(n_346), .B(n_516), .Y(n_696) );
AND2x2_ASAP7_75t_L g698 ( .A(n_346), .B(n_375), .Y(n_698) );
INVx1_ASAP7_75t_L g713 ( .A(n_346), .Y(n_713) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g400 ( .A(n_349), .B(n_381), .Y(n_400) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g380 ( .A(n_350), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g424 ( .A(n_351), .Y(n_424) );
INVx6_ASAP7_75t_L g538 ( .A(n_351), .Y(n_538) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g376 ( .A(n_352), .Y(n_376) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g395 ( .A(n_353), .B(n_389), .Y(n_395) );
AND2x2_ASAP7_75t_L g412 ( .A(n_353), .B(n_355), .Y(n_412) );
INVx1_ASAP7_75t_L g368 ( .A(n_354), .Y(n_368) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g397 ( .A(n_355), .B(n_387), .Y(n_397) );
NOR2xp67_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_357), .A2(n_551), .B1(n_559), .B2(n_583), .Y(n_558) );
INVx2_ASAP7_75t_L g717 ( .A(n_357), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g945 ( .A1(n_357), .A2(n_789), .B1(n_946), .B2(n_961), .Y(n_945) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g378 ( .A(n_358), .B(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g640 ( .A(n_358), .Y(n_640) );
OR2x6_ASAP7_75t_L g652 ( .A(n_358), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_360), .B(n_721), .Y(n_1070) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_361), .Y(n_1065) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g451 ( .A(n_362), .Y(n_451) );
INVx2_ASAP7_75t_L g1352 ( .A(n_362), .Y(n_1352) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_377), .C(n_408), .Y(n_363) );
INVx2_ASAP7_75t_L g668 ( .A(n_365), .Y(n_668) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_365), .Y(n_1056) );
INVx2_ASAP7_75t_L g1327 ( .A(n_365), .Y(n_1327) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_366), .B(n_369), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g516 ( .A(n_367), .Y(n_516) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
OR2x6_ASAP7_75t_L g373 ( .A(n_370), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
OR2x2_ASAP7_75t_L g669 ( .A(n_370), .B(n_374), .Y(n_669) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g419 ( .A(n_372), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g1329 ( .A(n_373), .Y(n_1329) );
OR2x2_ASAP7_75t_L g924 ( .A(n_374), .B(n_713), .Y(n_924) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI22xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_382), .B1(n_398), .B2(n_401), .Y(n_377) );
INVx3_ASAP7_75t_L g1315 ( .A(n_378), .Y(n_1315) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g534 ( .A(n_380), .Y(n_534) );
INVx2_ASAP7_75t_L g653 ( .A(n_380), .Y(n_653) );
INVx1_ASAP7_75t_L g702 ( .A(n_380), .Y(n_702) );
INVx2_ASAP7_75t_SL g937 ( .A(n_380), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g929 ( .A1(n_383), .A2(n_430), .B1(n_904), .B2(n_906), .C(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g524 ( .A(n_384), .Y(n_524) );
INVx2_ASAP7_75t_L g1048 ( .A(n_384), .Y(n_1048) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g403 ( .A(n_385), .Y(n_403) );
OR2x2_ASAP7_75t_L g546 ( .A(n_385), .B(n_420), .Y(n_546) );
INVx1_ASAP7_75t_L g866 ( .A(n_385), .Y(n_866) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
AND2x2_ASAP7_75t_L g392 ( .A(n_386), .B(n_388), .Y(n_392) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_390), .A2(n_402), .B1(n_404), .B2(n_405), .C(n_406), .Y(n_401) );
INVx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g1041 ( .A(n_391), .Y(n_1041) );
INVx1_ASAP7_75t_L g1050 ( .A(n_391), .Y(n_1050) );
BUFx4f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
INVx1_ASAP7_75t_L g523 ( .A(n_392), .Y(n_523) );
BUFx2_ASAP7_75t_L g701 ( .A(n_394), .Y(n_701) );
INVx1_ASAP7_75t_L g927 ( .A(n_394), .Y(n_927) );
BUFx3_ASAP7_75t_L g934 ( .A(n_394), .Y(n_934) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_395), .Y(n_407) );
INVx2_ASAP7_75t_SL g417 ( .A(n_395), .Y(n_417) );
BUFx2_ASAP7_75t_L g530 ( .A(n_395), .Y(n_530) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_395), .Y(n_565) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_395), .Y(n_572) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_395), .Y(n_662) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_395), .Y(n_783) );
BUFx3_ASAP7_75t_L g1323 ( .A(n_395), .Y(n_1323) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_396), .Y(n_521) );
BUFx3_ASAP7_75t_L g928 ( .A(n_396), .Y(n_928) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_397), .Y(n_541) );
INVx2_ASAP7_75t_L g549 ( .A(n_397), .Y(n_549) );
INVx1_ASAP7_75t_L g1046 ( .A(n_397), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_398), .A2(n_652), .B1(n_1037), .B2(n_1047), .Y(n_1036) );
INVx4_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_399), .A2(n_644), .B1(n_651), .B2(n_654), .C(n_666), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_400), .A2(n_446), .B1(n_449), .B2(n_523), .C(n_524), .Y(n_522) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_400), .A2(n_523), .B1(n_524), .B2(n_567), .C(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g689 ( .A(n_400), .Y(n_689) );
INVx2_ASAP7_75t_SL g781 ( .A(n_400), .Y(n_781) );
INVx1_ASAP7_75t_L g881 ( .A(n_400), .Y(n_881) );
HB1xp67_ASAP7_75t_L g930 ( .A(n_400), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_400), .Y(n_1026) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g511 ( .A(n_407), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_SL g692 ( .A(n_407), .Y(n_692) );
BUFx3_ASAP7_75t_L g1053 ( .A(n_407), .Y(n_1053) );
BUFx2_ASAP7_75t_L g1054 ( .A(n_408), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1326 ( .A1(n_408), .A2(n_1327), .B1(n_1328), .B2(n_1329), .C(n_1330), .Y(n_1326) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_411), .Y(n_647) );
INVx2_ASAP7_75t_L g773 ( .A(n_411), .Y(n_773) );
BUFx6f_ASAP7_75t_L g1025 ( .A(n_411), .Y(n_1025) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_412), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_413), .B(n_657), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_421), .B1(n_422), .B2(n_425), .C(n_426), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_415), .A2(n_422), .B1(n_672), .B2(n_673), .C(n_674), .Y(n_671) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g520 ( .A(n_417), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_417), .A2(n_540), .B1(n_633), .B2(n_635), .Y(n_650) );
INVx2_ASAP7_75t_SL g1317 ( .A(n_417), .Y(n_1317) );
AND2x2_ASAP7_75t_L g422 ( .A(n_418), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OR2x6_ASAP7_75t_L g427 ( .A(n_419), .B(n_428), .Y(n_427) );
OR2x6_ASAP7_75t_L g429 ( .A(n_419), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g675 ( .A(n_419), .B(n_428), .Y(n_675) );
OR2x2_ASAP7_75t_L g1088 ( .A(n_419), .B(n_524), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_419), .B(n_864), .Y(n_1089) );
INVx2_ASAP7_75t_L g512 ( .A(n_420), .Y(n_512) );
OR2x2_ASAP7_75t_L g548 ( .A(n_420), .B(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g658 ( .A(n_423), .Y(n_658) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g939 ( .A(n_424), .Y(n_939) );
INVx2_ASAP7_75t_L g1324 ( .A(n_428), .Y(n_1324) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_432), .A2(n_1111), .B1(n_1116), .B2(n_1132), .Y(n_1131) );
XNOR2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_608), .Y(n_433) );
AO22x2_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_555), .B2(n_556), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
XNOR2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_507), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_455), .C(n_466), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_448), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_446), .B2(n_447), .Y(n_441) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g588 ( .A(n_444), .Y(n_588) );
BUFx2_ASAP7_75t_L g731 ( .A(n_444), .Y(n_731) );
BUFx2_ASAP7_75t_L g888 ( .A(n_444), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_444), .A2(n_447), .B1(n_965), .B2(n_966), .Y(n_964) );
AND2x4_ASAP7_75t_L g450 ( .A(n_445), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g453 ( .A(n_445), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g591 ( .A(n_445), .B(n_454), .Y(n_591) );
AND2x2_ASAP7_75t_L g794 ( .A(n_445), .B(n_495), .Y(n_794) );
AND2x2_ASAP7_75t_L g796 ( .A(n_445), .B(n_745), .Y(n_796) );
AND2x2_ASAP7_75t_L g800 ( .A(n_445), .B(n_454), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g1005 ( .A1(n_445), .A2(n_1006), .B1(n_1010), .B2(n_1011), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_447), .A2(n_567), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_447), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_447), .A2(n_588), .B1(n_903), .B2(n_904), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B1(n_452), .B2(n_453), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_450), .A2(n_568), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_450), .A2(n_453), .B1(n_734), .B2(n_735), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_450), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_797) );
INVx1_ASAP7_75t_L g886 ( .A(n_450), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_450), .A2(n_591), .B1(n_906), .B2(n_907), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_450), .A2(n_591), .B1(n_968), .B2(n_969), .Y(n_967) );
INVx1_ASAP7_75t_L g621 ( .A(n_451), .Y(n_621) );
BUFx3_ASAP7_75t_L g751 ( .A(n_451), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_451), .A2(n_728), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_458), .Y(n_971) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_459), .B(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g720 ( .A(n_459), .B(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g723 ( .A(n_459), .B(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g727 ( .A(n_459), .B(n_728), .Y(n_727) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx4f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx4f_ASAP7_75t_L g832 ( .A(n_462), .Y(n_832) );
BUFx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g802 ( .A(n_465), .Y(n_802) );
OAI33xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_470), .A3(n_478), .B1(n_486), .B2(n_497), .B3(n_504), .Y(n_466) );
OAI33xp33_ASAP7_75t_L g593 ( .A1(n_467), .A2(n_504), .A3(n_594), .B1(n_598), .B2(n_601), .B3(n_605), .Y(n_593) );
OAI33xp33_ASAP7_75t_L g803 ( .A1(n_467), .A2(n_804), .A3(n_811), .B1(n_816), .B2(n_819), .B3(n_821), .Y(n_803) );
OAI33xp33_ASAP7_75t_L g972 ( .A1(n_467), .A2(n_504), .A3(n_973), .B1(n_977), .B2(n_981), .B3(n_984), .Y(n_972) );
OAI22xp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_475), .B2(n_476), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_472), .A2(n_498), .B1(n_499), .B2(n_503), .Y(n_497) );
OAI22xp33_ASAP7_75t_L g594 ( .A1(n_472), .A2(n_595), .B1(n_596), .B2(n_597), .Y(n_594) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_SL g974 ( .A(n_473), .Y(n_974) );
INVx2_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g1075 ( .A(n_477), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_483), .B2(n_484), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_480), .A2(n_484), .B1(n_599), .B2(n_600), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_480), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_480), .A2(n_950), .B1(n_960), .B2(n_982), .Y(n_981) );
BUFx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_482), .Y(n_632) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_491), .B1(n_492), .B2(n_496), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g602 ( .A(n_488), .Y(n_602) );
INVx1_ASAP7_75t_L g1060 ( .A(n_488), .Y(n_1060) );
INVx2_ASAP7_75t_L g1078 ( .A(n_488), .Y(n_1078) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_489), .A2(n_1340), .B1(n_1341), .B2(n_1342), .Y(n_1339) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx3_ASAP7_75t_L g813 ( .A(n_490), .Y(n_813) );
AOI211xp5_ASAP7_75t_SL g510 ( .A1(n_491), .A2(n_511), .B(n_513), .C(n_519), .Y(n_510) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g983 ( .A(n_494), .Y(n_983) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g618 ( .A(n_495), .Y(n_618) );
INVx1_ASAP7_75t_L g845 ( .A(n_495), .Y(n_845) );
INVx2_ASAP7_75t_L g979 ( .A(n_495), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_496), .A2(n_498), .B1(n_545), .B2(n_547), .Y(n_544) );
OAI22xp5_ASAP7_75t_SL g847 ( .A1(n_499), .A2(n_848), .B1(n_849), .B2(n_851), .Y(n_847) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g597 ( .A(n_501), .Y(n_597) );
BUFx3_ASAP7_75t_L g820 ( .A(n_501), .Y(n_820) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_503), .A2(n_526), .B1(n_529), .B2(n_535), .C(n_542), .Y(n_525) );
CKINVDCx8_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
INVx5_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx6_ASAP7_75t_L g752 ( .A(n_506), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_550), .B2(n_551), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_525), .C(n_544), .Y(n_509) );
AOI211xp5_ASAP7_75t_SL g560 ( .A1(n_511), .A2(n_561), .B(n_562), .C(n_564), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_511), .A2(n_684), .B1(n_690), .B2(n_693), .C(n_694), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g920 ( .A1(n_511), .A2(n_921), .B(n_922), .C(n_925), .Y(n_920) );
AND2x4_ASAP7_75t_L g527 ( .A(n_512), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g778 ( .A(n_512), .B(n_662), .Y(n_778) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_512), .A2(n_527), .B1(n_542), .B2(n_851), .C(n_863), .Y(n_862) );
AOI222xp33_ASAP7_75t_L g1016 ( .A1(n_512), .A2(n_515), .B1(n_518), .B2(n_994), .C1(n_995), .C2(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g859 ( .A(n_514), .Y(n_859) );
INVx4_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_SL g786 ( .A(n_515), .Y(n_786) );
INVx2_ASAP7_75t_L g952 ( .A(n_515), .Y(n_952) );
INVx2_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g563 ( .A(n_518), .Y(n_563) );
AOI222xp33_ASAP7_75t_SL g855 ( .A1(n_518), .A2(n_856), .B1(n_858), .B2(n_859), .C1(n_860), .C2(n_861), .Y(n_855) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_527), .A2(n_542), .B1(n_570), .B2(n_571), .C(n_574), .Y(n_569) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_527), .Y(n_709) );
INVx2_ASAP7_75t_SL g769 ( .A(n_527), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_527), .A2(n_542), .B1(n_954), .B2(n_955), .C(n_957), .Y(n_953) );
INVx2_ASAP7_75t_SL g532 ( .A(n_528), .Y(n_532) );
AND2x4_ASAP7_75t_L g542 ( .A(n_528), .B(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_528), .Y(n_657) );
BUFx4f_ASAP7_75t_L g870 ( .A(n_528), .Y(n_870) );
INVx1_ASAP7_75t_L g879 ( .A(n_528), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_528), .A2(n_662), .B1(n_1014), .B2(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g573 ( .A(n_532), .Y(n_573) );
INVxp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx3_ASAP7_75t_L g774 ( .A(n_534), .Y(n_774) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g705 ( .A(n_537), .Y(n_705) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_538), .Y(n_576) );
INVx2_ASAP7_75t_L g649 ( .A(n_538), .Y(n_649) );
INVx1_ASAP7_75t_L g880 ( .A(n_538), .Y(n_880) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g784 ( .A(n_540), .Y(n_784) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g665 ( .A(n_541), .Y(n_665) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_541), .Y(n_708) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_541), .Y(n_776) );
INVx2_ASAP7_75t_L g867 ( .A(n_541), .Y(n_867) );
BUFx6f_ASAP7_75t_L g1318 ( .A(n_541), .Y(n_1318) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_542), .A2(n_768), .B1(n_770), .B2(n_771), .C(n_775), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g1020 ( .A1(n_542), .A2(n_1021), .B(n_1022), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_545), .A2(n_547), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_545), .A2(n_547), .B1(n_715), .B2(n_716), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_545), .A2(n_547), .B1(n_765), .B2(n_766), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_545), .A2(n_547), .B1(n_941), .B2(n_942), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_545), .A2(n_547), .B1(n_959), .B2(n_960), .Y(n_958) );
INVx6_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g579 ( .A(n_549), .Y(n_579) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx5_ASAP7_75t_L g680 ( .A(n_552), .Y(n_680) );
INVx2_ASAP7_75t_SL g789 ( .A(n_552), .Y(n_789) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx2_ASAP7_75t_L g1004 ( .A(n_553), .Y(n_1004) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_584), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_569), .C(n_580), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_561), .A2(n_582), .B1(n_602), .B2(n_603), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_570), .A2(n_581), .B1(n_606), .B2(n_607), .Y(n_605) );
BUFx3_ASAP7_75t_L g873 ( .A(n_572), .Y(n_873) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx4_ASAP7_75t_L g687 ( .A(n_576), .Y(n_687) );
INVx1_ASAP7_75t_L g875 ( .A(n_577), .Y(n_875) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g956 ( .A(n_578), .Y(n_956) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NOR3xp33_ASAP7_75t_SL g584 ( .A(n_585), .B(n_592), .C(n_593), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
OAI22xp33_ASAP7_75t_L g973 ( .A1(n_597), .A2(n_974), .B1(n_975), .B2(n_976), .Y(n_973) );
INVx2_ASAP7_75t_SL g749 ( .A(n_603), .Y(n_749) );
OAI22xp33_ASAP7_75t_L g834 ( .A1(n_603), .A2(n_835), .B1(n_836), .B2(n_837), .Y(n_834) );
INVx4_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx3_ASAP7_75t_L g747 ( .A(n_604), .Y(n_747) );
INVx2_ASAP7_75t_SL g914 ( .A(n_604), .Y(n_914) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_606), .A2(n_765), .B1(n_770), .B2(n_820), .Y(n_819) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_607), .A2(n_637), .B(n_638), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_676), .B1(n_753), .B2(n_754), .Y(n_608) );
INVx1_ASAP7_75t_L g753 ( .A(n_609), .Y(n_753) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_641), .C(n_643), .D(n_671), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_629), .B(n_640), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_619), .B(n_625), .Y(n_613) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g1062 ( .A(n_617), .Y(n_1062) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g1066 ( .A(n_624), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_627), .A2(n_628), .B1(n_660), .B2(n_663), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_633), .B1(n_634), .B2(n_635), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_631), .A2(n_766), .B1(n_779), .B2(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_634), .A2(n_812), .B1(n_814), .B2(n_815), .Y(n_811) );
CKINVDCx8_ASAP7_75t_R g787 ( .A(n_640), .Y(n_787) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g686 ( .A(n_647), .Y(n_686) );
AND2x4_ASAP7_75t_L g711 ( .A(n_647), .B(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx4f_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g864 ( .A(n_662), .Y(n_864) );
BUFx2_ASAP7_75t_L g1044 ( .A(n_662), .Y(n_1044) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI221xp5_ASAP7_75t_SL g868 ( .A1(n_665), .A2(n_837), .B1(n_840), .B2(n_865), .C(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_676), .Y(n_754) );
XNOR2x1_ASAP7_75t_SL g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_718), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B(n_682), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g917 ( .A1(n_680), .A2(n_918), .B(n_919), .Y(n_917) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_699), .A3(n_714), .B(n_717), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g923 ( .A(n_696), .Y(n_923) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B1(n_709), .B2(n_710), .C(n_711), .Y(n_699) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_709), .A2(n_711), .B1(n_932), .B2(n_933), .C(n_938), .Y(n_931) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
AOI31xp33_ASAP7_75t_SL g1015 ( .A1(n_717), .A2(n_1016), .A3(n_1020), .B(n_1023), .Y(n_1015) );
OAI31xp33_ASAP7_75t_L g1057 ( .A1(n_717), .A2(n_1058), .A3(n_1073), .B(n_1080), .Y(n_1057) );
AND4x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_729), .C(n_733), .D(n_736), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_722), .B1(n_723), .B2(n_726), .C(n_727), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g889 ( .A1(n_720), .A2(n_727), .B(n_860), .Y(n_889) );
INVx1_ASAP7_75t_L g900 ( .A(n_720), .Y(n_900) );
AOI221xp5_ASAP7_75t_L g993 ( .A1(n_720), .A2(n_723), .B1(n_727), .B2(n_994), .C(n_995), .Y(n_993) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_723), .Y(n_897) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_727), .A2(n_897), .B1(n_898), .B2(n_899), .C(n_901), .Y(n_896) );
AOI33xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_740), .A3(n_746), .B1(n_748), .B2(n_750), .B3(n_752), .Y(n_736) );
AOI33xp33_ASAP7_75t_L g908 ( .A1(n_737), .A2(n_752), .A3(n_909), .B1(n_911), .B2(n_915), .B3(n_916), .Y(n_908) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g910 ( .A(n_744), .Y(n_910) );
INVx2_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g821 ( .A(n_752), .Y(n_821) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
XNOR2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_890), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_824), .B2(n_825), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g822 ( .A(n_761), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_790), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .C(n_777), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g1321 ( .A(n_773), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_779), .B1(n_780), .B2(n_782), .C(n_785), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_778), .A2(n_948), .B1(n_949), .B2(n_950), .C(n_951), .Y(n_947) );
NOR3xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_801), .C(n_803), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_792), .B(n_797), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_792) );
INVxp67_ASAP7_75t_L g852 ( .A(n_796), .Y(n_852) );
INVx1_ASAP7_75t_L g831 ( .A(n_800), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_807), .B1(n_808), .B2(n_810), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_808), .A2(n_957), .B1(n_959), .B2(n_974), .Y(n_984) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g836 ( .A(n_813), .Y(n_836) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_853), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_833), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_845), .B2(n_846), .Y(n_841) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AOI21xp5_ASAP7_75t_SL g853 ( .A1(n_854), .A2(n_882), .B(n_885), .Y(n_853) );
NAND4xp25_ASAP7_75t_SL g854 ( .A(n_855), .B(n_862), .C(n_868), .D(n_871), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g1023 ( .A1(n_856), .A2(n_1003), .B1(n_1024), .B2(n_1027), .Y(n_1023) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_865), .Y(n_1038) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_874), .B1(n_875), .B2(n_876), .C(n_877), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
AOI31xp33_ASAP7_75t_L g919 ( .A1(n_883), .A2(n_920), .A3(n_931), .B(n_940), .Y(n_919) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AOI21x1_ASAP7_75t_L g1331 ( .A1(n_884), .A2(n_1332), .B(n_1343), .Y(n_1331) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
XNOR2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_988), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_892), .A2(n_893), .B1(n_943), .B2(n_987), .Y(n_891) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_895), .B(n_917), .Y(n_894) );
AND4x1_ASAP7_75t_L g895 ( .A(n_896), .B(n_902), .C(n_905), .D(n_908), .Y(n_895) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_SL g1076 ( .A1(n_914), .A2(n_1077), .B1(n_1078), .B2(n_1079), .Y(n_1076) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx3_ASAP7_75t_L g987 ( .A(n_943), .Y(n_987) );
INVx1_ASAP7_75t_L g985 ( .A(n_944), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_962), .Y(n_944) );
NAND3xp33_ASAP7_75t_L g946 ( .A(n_947), .B(n_953), .C(n_958), .Y(n_946) );
NOR3xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_970), .C(n_972), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_967), .Y(n_963) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_1032), .B1(n_1033), .B2(n_1090), .Y(n_988) );
INVx1_ASAP7_75t_L g1090 ( .A(n_989), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
NAND2xp5_ASAP7_75t_SL g990 ( .A(n_991), .B(n_1028), .Y(n_990) );
INVx1_ASAP7_75t_L g1030 ( .A(n_992), .Y(n_1030) );
NAND3xp33_ASAP7_75t_SL g992 ( .A(n_993), .B(n_996), .C(n_1005), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B1(n_1003), .B2(n_1004), .Y(n_996) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1015), .Y(n_1029) );
NAND3xp33_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1030), .C(n_1031), .Y(n_1028) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
AND4x1_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1057), .C(n_1083), .D(n_1085), .Y(n_1034) );
NOR3xp33_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1054), .C(n_1055), .Y(n_1035) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1039), .B1(n_1040), .B2(n_1042), .C(n_1043), .Y(n_1037) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
OAI221xp5_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1050), .B2(n_1051), .C(n_1052), .Y(n_1047) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_1060), .A2(n_1061), .B1(n_1062), .B2(n_1063), .C(n_1064), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1070), .B1(n_1071), .B2(n_1072), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1087), .Y(n_1085) );
OAI221xp5_ASAP7_75t_L g1092 ( .A1(n_1093), .A2(n_1306), .B1(n_1308), .B2(n_1355), .C(n_1359), .Y(n_1092) );
NOR2x1_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1272), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1223), .Y(n_1094) );
NOR4xp25_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1165), .C(n_1185), .D(n_1201), .Y(n_1095) );
AOI21xp33_ASAP7_75t_L g1096 ( .A1(n_1097), .A2(n_1149), .B(n_1153), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1118), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1098), .B(n_1150), .Y(n_1229) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1098), .Y(n_1267) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1099), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1099), .B(n_1231), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1099), .B(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1099), .Y(n_1297) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1100), .B(n_1172), .Y(n_1171) );
INVx2_ASAP7_75t_SL g1184 ( .A(n_1100), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1199 ( .A(n_1100), .B(n_1172), .Y(n_1199) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1101), .Y(n_1163) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1101), .Y(n_1216) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1105), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1102), .B(n_1105), .Y(n_1129) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_1103), .B(n_1105), .Y(n_1107) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1104), .B(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1106), .Y(n_1114) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1107), .Y(n_1138) );
INVx1_ASAP7_75t_SL g1144 ( .A(n_1107), .Y(n_1144) );
OAI22xp33_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1110), .B1(n_1115), .B2(n_1116), .Y(n_1108) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_1110), .A2(n_1116), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
OAI22xp33_ASAP7_75t_L g1156 ( .A1(n_1110), .A2(n_1157), .B1(n_1158), .B2(n_1159), .Y(n_1156) );
BUFx3_ASAP7_75t_L g1220 ( .A(n_1110), .Y(n_1220) );
BUFx6f_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1113), .Y(n_1111) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1112), .B(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1112), .Y(n_1125) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1113), .Y(n_1124) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1116), .Y(n_1160) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1117), .Y(n_1127) );
A2O1A1Ixp33_ASAP7_75t_L g1165 ( .A1(n_1118), .A2(n_1166), .B(n_1170), .C(n_1175), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1133), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1119), .B(n_1169), .Y(n_1168) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_1119), .A2(n_1195), .B(n_1196), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1249 ( .A(n_1119), .B(n_1207), .C(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1256 ( .A(n_1120), .B(n_1134), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1120), .B(n_1140), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1130), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1121), .B(n_1130), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1121), .B(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1121), .Y(n_1189) );
O2A1O1Ixp33_ASAP7_75t_SL g1201 ( .A1(n_1121), .A2(n_1202), .B(n_1205), .C(n_1212), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1121), .B(n_1140), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1128), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1125), .Y(n_1123) );
OAI21xp33_ASAP7_75t_SL g1369 ( .A1(n_1124), .A2(n_1363), .B(n_1370), .Y(n_1369) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1125), .B(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1129), .Y(n_1142) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1130), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1130), .B(n_1139), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1130), .B(n_1189), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1130), .B(n_1133), .Y(n_1228) );
AOI32xp33_ASAP7_75t_L g1259 ( .A1(n_1130), .A2(n_1191), .A3(n_1243), .B1(n_1260), .B2(n_1261), .Y(n_1259) );
A2O1A1Ixp33_ASAP7_75t_L g1263 ( .A1(n_1130), .A2(n_1134), .B(n_1198), .C(n_1233), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1133), .B(n_1152), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1139), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1134), .B(n_1152), .Y(n_1151) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_1134), .B(n_1139), .Y(n_1169) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1134), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1134), .B(n_1155), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1134), .B(n_1204), .Y(n_1203) );
INVx4_ASAP7_75t_L g1241 ( .A(n_1134), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1134), .B(n_1245), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1134), .B(n_1246), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1300 ( .A(n_1134), .B(n_1277), .Y(n_1300) );
AND2x6_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_1138), .A2(n_1215), .B1(n_1216), .B2(n_1217), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1150 ( .A(n_1139), .B(n_1151), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1139), .B(n_1177), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1139), .B(n_1178), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1139), .B(n_1211), .Y(n_1269) );
CKINVDCx6p67_ASAP7_75t_R g1139 ( .A(n_1140), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1140), .B(n_1189), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1140), .B(n_1189), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1140), .B(n_1177), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1140), .B(n_1211), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1140), .B(n_1152), .Y(n_1254) );
OAI211xp5_ASAP7_75t_SL g1258 ( .A1(n_1140), .A2(n_1186), .B(n_1259), .C(n_1263), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1140), .B(n_1266), .Y(n_1265) );
OR2x6_ASAP7_75t_SL g1140 ( .A(n_1141), .B(n_1146), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1143), .B1(n_1144), .B2(n_1145), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g1161 ( .A1(n_1144), .A2(n_1162), .B1(n_1163), .B2(n_1164), .Y(n_1161) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1152), .B(n_1241), .Y(n_1266) );
INVx1_ASAP7_75t_SL g1243 ( .A(n_1153), .Y(n_1243) );
INVx3_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1154), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1154), .B(n_1172), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1154), .B(n_1213), .Y(n_1212) );
OAI211xp5_ASAP7_75t_L g1224 ( .A1(n_1154), .A2(n_1225), .B(n_1229), .C(n_1230), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1154), .B(n_1171), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1154), .B(n_1184), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1154), .B(n_1207), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1154), .B(n_1246), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1154), .B(n_1172), .Y(n_1301) );
INVx3_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1155), .B(n_1172), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1155), .B(n_1199), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1161), .Y(n_1155) );
HB1xp67_ASAP7_75t_L g1222 ( .A(n_1159), .Y(n_1222) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_1168), .B(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g1238 ( .A1(n_1171), .A2(n_1239), .B1(n_1242), .B2(n_1247), .C(n_1248), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1171), .B(n_1240), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1273 ( .A1(n_1171), .A2(n_1274), .B1(n_1280), .B2(n_1283), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1172), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1172), .B(n_1184), .Y(n_1204) );
INVx2_ASAP7_75t_L g1207 ( .A(n_1172), .Y(n_1207) );
AND2x4_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1174), .Y(n_1172) );
OAI21xp5_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1179), .B(n_1182), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_1176), .A2(n_1232), .B1(n_1241), .B2(n_1269), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1176), .B(n_1241), .Y(n_1294) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1177), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1177), .B(n_1240), .Y(n_1239) );
O2A1O1Ixp33_ASAP7_75t_L g1295 ( .A1(n_1179), .A2(n_1226), .B(n_1287), .C(n_1296), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1181), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1180), .B(n_1192), .Y(n_1191) );
NOR2xp33_ASAP7_75t_L g1206 ( .A(n_1180), .B(n_1207), .Y(n_1206) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1180), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1182), .B(n_1187), .Y(n_1186) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1246 ( .A(n_1184), .Y(n_1246) );
OAI221xp5_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1188), .B1(n_1190), .B2(n_1193), .C(n_1194), .Y(n_1185) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1188), .Y(n_1192) );
OAI211xp5_ASAP7_75t_SL g1248 ( .A1(n_1188), .A2(n_1193), .B(n_1249), .C(n_1252), .Y(n_1248) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1200), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1198), .B(n_1241), .Y(n_1283) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_1199), .A2(n_1226), .B1(n_1227), .B2(n_1228), .Y(n_1225) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1204), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1207), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .Y(n_1208) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g1252 ( .A(n_1213), .Y(n_1252) );
OR2x6_ASAP7_75t_SL g1213 ( .A(n_1214), .B(n_1218), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1220), .B1(n_1221), .B2(n_1222), .Y(n_1218) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1220), .Y(n_1307) );
OAI32xp33_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1234), .A3(n_1252), .B1(n_1258), .B2(n_1264), .Y(n_1223) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1226), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1233), .Y(n_1231) );
OAI211xp5_ASAP7_75t_SL g1234 ( .A1(n_1235), .A2(n_1236), .B(n_1238), .C(n_1253), .Y(n_1234) );
OAI21xp33_ASAP7_75t_L g1299 ( .A1(n_1235), .A2(n_1241), .B(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1237), .B(n_1254), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_1240), .B(n_1247), .Y(n_1303) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1244), .Y(n_1242) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1244), .Y(n_1288) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
A2O1A1Ixp33_ASAP7_75t_SL g1272 ( .A1(n_1252), .A2(n_1273), .B(n_1284), .C(n_1298), .Y(n_1272) );
OAI21xp5_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1255), .B(n_1257), .Y(n_1253) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
A2O1A1Ixp33_ASAP7_75t_L g1302 ( .A1(n_1256), .A2(n_1303), .B(n_1304), .C(n_1305), .Y(n_1302) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
O2A1O1Ixp33_ASAP7_75t_SL g1264 ( .A1(n_1265), .A2(n_1267), .B(n_1268), .C(n_1270), .Y(n_1264) );
O2A1O1Ixp33_ASAP7_75t_L g1284 ( .A1(n_1269), .A2(n_1285), .B(n_1288), .C(n_1289), .Y(n_1284) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
NOR2xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1278), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
A2O1A1Ixp33_ASAP7_75t_L g1289 ( .A1(n_1290), .A2(n_1291), .B(n_1293), .C(n_1295), .Y(n_1289) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
AOI21xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1301), .B(n_1302), .Y(n_1298) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
HB1xp67_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVxp67_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1312), .Y(n_1367) );
NOR4xp75_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1331), .C(n_1353), .D(n_1354), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1326), .Y(n_1313) );
AOI33xp33_ASAP7_75t_L g1314 ( .A1(n_1315), .A2(n_1316), .A3(n_1319), .B1(n_1320), .B2(n_1322), .B3(n_1325), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1351), .B(n_1352), .Y(n_1350) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
CKINVDCx5p33_ASAP7_75t_R g1361 ( .A(n_1362), .Y(n_1361) );
INVxp33_ASAP7_75t_SL g1364 ( .A(n_1365), .Y(n_1364) );
HB1xp67_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
endmodule