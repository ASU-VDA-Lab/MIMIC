module fake_jpeg_10813_n_595 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_595);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_595;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_12),
.B(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g201 ( 
.A(n_60),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_67),
.Y(n_138)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_21),
.B(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_70),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g164 ( 
.A(n_75),
.Y(n_164)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_30),
.B(n_15),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_81),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_21),
.B(n_41),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_25),
.Y(n_144)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_16),
.Y(n_95)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_43),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_31),
.B(n_10),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_103),
.B(n_111),
.Y(n_194)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_49),
.B(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_113),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_39),
.Y(n_114)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_115),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_118),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx5_ASAP7_75t_SL g186 ( 
.A(n_120),
.Y(n_186)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_42),
.Y(n_130)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_57),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_130),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_37),
.B1(n_20),
.B2(n_48),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_131),
.A2(n_170),
.B(n_171),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_139),
.B(n_177),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_144),
.B(n_148),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_67),
.A2(n_25),
.B(n_23),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_145),
.A2(n_15),
.B(n_9),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_56),
.B1(n_54),
.B2(n_34),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_147),
.A2(n_38),
.B1(n_51),
.B2(n_112),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_46),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_188),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_81),
.A2(n_34),
.B1(n_56),
.B2(n_54),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_80),
.B1(n_109),
.B2(n_106),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_60),
.B(n_31),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_162),
.B(n_173),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_59),
.A2(n_48),
.B1(n_42),
.B2(n_20),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_84),
.A2(n_56),
.B1(n_57),
.B2(n_53),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_75),
.B(n_46),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_72),
.A2(n_57),
.B1(n_53),
.B2(n_32),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_164),
.B1(n_146),
.B2(n_157),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_100),
.B(n_45),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_89),
.B(n_45),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_33),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_33),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_0),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_71),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_23),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

BUFx2_ASAP7_75t_SL g277 ( 
.A(n_202),
.Y(n_277)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_203),
.Y(n_301)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_194),
.A2(n_51),
.B(n_41),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_206),
.B(n_6),
.Y(n_312)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_208),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_209),
.A2(n_211),
.B1(n_258),
.B2(n_270),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_138),
.A2(n_119),
.B1(n_117),
.B2(n_116),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_216),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_218),
.B(n_242),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_221),
.Y(n_323)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_222),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_146),
.A2(n_64),
.B1(n_105),
.B2(n_102),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_223),
.A2(n_260),
.B1(n_261),
.B2(n_266),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_133),
.Y(n_227)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_227),
.Y(n_300)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_161),
.A2(n_88),
.B1(n_74),
.B2(n_82),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_230),
.A2(n_243),
.B1(n_250),
.B2(n_254),
.Y(n_317)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_164),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_155),
.Y(n_234)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_234),
.Y(n_310)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_235),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_130),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_237),
.Y(n_313)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_240),
.Y(n_328)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_125),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_245),
.Y(n_286)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_246),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_194),
.A2(n_9),
.B(n_38),
.Y(n_247)
);

NAND2x1_ASAP7_75t_SL g314 ( 
.A(n_247),
.B(n_6),
.Y(n_314)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_152),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_182),
.A2(n_90),
.B1(n_83),
.B2(n_65),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_145),
.A2(n_114),
.B1(n_113),
.B2(n_2),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_256),
.Y(n_319)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_183),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_257),
.B(n_267),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_135),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_186),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_259),
.B(n_262),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_129),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_263),
.A2(n_272),
.B1(n_185),
.B2(n_165),
.Y(n_321)
);

OA22x2_ASAP7_75t_SL g264 ( 
.A1(n_131),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_156),
.B(n_140),
.Y(n_283)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_190),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_265),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_152),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_268),
.Y(n_307)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_178),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_269),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_170),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_129),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_271),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_141),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_220),
.A2(n_176),
.B(n_184),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_280),
.A2(n_292),
.B(n_308),
.Y(n_371)
);

AOI32xp33_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_146),
.A3(n_137),
.B1(n_140),
.B2(n_153),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_282),
.A2(n_308),
.B(n_313),
.C(n_311),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_283),
.B(n_7),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_229),
.A2(n_153),
.B1(n_189),
.B2(n_180),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_287),
.A2(n_321),
.B1(n_329),
.B2(n_198),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_229),
.A2(n_165),
.B1(n_198),
.B2(n_185),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_290),
.A2(n_250),
.B1(n_203),
.B2(n_226),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_219),
.A2(n_142),
.B(n_168),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_150),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_295),
.B(n_296),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_150),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_253),
.A2(n_134),
.B(n_154),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_304),
.B(n_312),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_252),
.A2(n_180),
.B(n_189),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_218),
.B(n_205),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_253),
.B(n_200),
.C(n_151),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_223),
.C(n_271),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_230),
.A2(n_141),
.B1(n_200),
.B2(n_151),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_296),
.B(n_205),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_330),
.B(n_335),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_336),
.C(n_337),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_355),
.Y(n_392)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_280),
.A2(n_214),
.B(n_210),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_334),
.A2(n_347),
.B(n_352),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_213),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_202),
.C(n_262),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_247),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_264),
.C(n_266),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_349),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_207),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_340),
.B(n_342),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_279),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_357),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_235),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_344),
.A2(n_366),
.B1(n_278),
.B2(n_294),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_326),
.A2(n_264),
.B1(n_196),
.B2(n_224),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_345),
.A2(n_348),
.B1(n_356),
.B2(n_364),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_346),
.A2(n_294),
.B1(n_278),
.B2(n_289),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_305),
.A2(n_208),
.B(n_246),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_326),
.A2(n_196),
.B1(n_212),
.B2(n_217),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g349 ( 
.A(n_305),
.B(n_237),
.C(n_268),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_314),
.A2(n_221),
.B(n_260),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_350),
.A2(n_365),
.B(n_372),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_7),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_354),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_273),
.A2(n_7),
.B(n_261),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_353),
.A2(n_360),
.B(n_325),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_281),
.B(n_312),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_276),
.B(n_293),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_273),
.A2(n_292),
.B1(n_317),
.B2(n_285),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_297),
.Y(n_357)
);

AND2x2_ASAP7_75t_SL g358 ( 
.A(n_283),
.B(n_282),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_367),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_276),
.B(n_293),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_361),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_286),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_299),
.Y(n_362)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_362),
.Y(n_375)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_302),
.A2(n_284),
.B1(n_322),
.B2(n_318),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_319),
.B(n_284),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_298),
.Y(n_366)
);

BUFx2_ASAP7_75t_SL g367 ( 
.A(n_298),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_368),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_302),
.B(n_275),
.Y(n_369)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_369),
.Y(n_391)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_301),
.B(n_275),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_358),
.A2(n_329),
.B1(n_311),
.B2(n_313),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_377),
.A2(n_380),
.B1(n_386),
.B2(n_401),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_370),
.Y(n_381)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

AOI32xp33_ASAP7_75t_L g382 ( 
.A1(n_334),
.A2(n_315),
.A3(n_307),
.B1(n_318),
.B2(n_328),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_382),
.A2(n_400),
.B(n_404),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_383),
.A2(n_344),
.B1(n_341),
.B2(n_367),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_372),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_384),
.B(n_373),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_338),
.A2(n_294),
.A3(n_310),
.B1(n_328),
.B2(n_324),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_390),
.B(n_369),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_359),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_355),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_360),
.A2(n_307),
.B(n_301),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_358),
.A2(n_288),
.B1(n_291),
.B2(n_278),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_356),
.A2(n_323),
.B1(n_315),
.B2(n_291),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_403),
.A2(n_405),
.B1(n_346),
.B2(n_277),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_348),
.A2(n_324),
.B1(n_300),
.B2(n_303),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_407),
.Y(n_427)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_409),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_330),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_417),
.C(n_420),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_412),
.A2(n_416),
.B1(n_419),
.B2(n_422),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_335),
.C(n_343),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_435),
.Y(n_445)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_415),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_409),
.A2(n_339),
.B1(n_353),
.B2(n_360),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_354),
.Y(n_417)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_418),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_353),
.B1(n_371),
.B2(n_331),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_336),
.C(n_338),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_398),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_441),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_391),
.A2(n_371),
.B1(n_361),
.B2(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_423),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_349),
.C(n_354),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_392),
.Y(n_451)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_429),
.Y(n_469)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_385),
.Y(n_432)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_373),
.B(n_343),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_433),
.B(n_434),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_365),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_323),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_436),
.A2(n_402),
.B1(n_387),
.B2(n_352),
.Y(n_464)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_438),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_379),
.B(n_392),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_379),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_374),
.A2(n_377),
.B1(n_380),
.B2(n_401),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_440),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_395),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_374),
.A2(n_332),
.B1(n_340),
.B2(n_351),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_442),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_395),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_390),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_431),
.A2(n_399),
.B1(n_397),
.B2(n_393),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_446),
.A2(n_462),
.B1(n_464),
.B2(n_474),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_407),
.Y(n_449)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_451),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_411),
.B(n_392),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_457),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_406),
.Y(n_455)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_455),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_456),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_417),
.B(n_397),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_423),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_438),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_SL g461 ( 
.A1(n_437),
.A2(n_400),
.B(n_371),
.C(n_388),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_461),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_428),
.A2(n_397),
.B1(n_393),
.B2(n_404),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_387),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_465),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_420),
.B(n_388),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_470),
.C(n_419),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_428),
.Y(n_468)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_349),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_437),
.A2(n_422),
.B1(n_424),
.B2(n_416),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_451),
.Y(n_503)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_477),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_432),
.C(n_430),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_478),
.B(n_480),
.C(n_491),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_429),
.C(n_427),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_413),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_482),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_458),
.A2(n_413),
.B1(n_426),
.B2(n_425),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_484),
.A2(n_490),
.B1(n_473),
.B2(n_469),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_448),
.B(n_410),
.Y(n_485)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_444),
.Y(n_488)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_488),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_471),
.A2(n_427),
.B1(n_426),
.B2(n_425),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_396),
.C(n_410),
.Y(n_491)
);

XOR2x1_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_412),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_470),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_381),
.Y(n_494)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_494),
.Y(n_518)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_444),
.Y(n_497)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_497),
.Y(n_519)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_447),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_500),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_452),
.B(n_396),
.C(n_347),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_461),
.C(n_337),
.Y(n_522)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_504),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_479),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_495),
.A2(n_445),
.B1(n_453),
.B2(n_463),
.Y(n_507)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_507),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_460),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_510),
.B(n_512),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_475),
.B(n_457),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_520),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_485),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_489),
.A2(n_472),
.B1(n_453),
.B2(n_461),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_514),
.A2(n_493),
.B1(n_484),
.B2(n_491),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_481),
.A2(n_446),
.B1(n_464),
.B2(n_462),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_490),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_489),
.A2(n_461),
.B1(n_450),
.B2(n_473),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_517),
.A2(n_513),
.B1(n_508),
.B2(n_502),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_521),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_479),
.C(n_476),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_496),
.B(n_381),
.Y(n_523)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_523),
.Y(n_540)
);

OAI221xp5_ASAP7_75t_L g525 ( 
.A1(n_509),
.A2(n_486),
.B1(n_480),
.B2(n_483),
.C(n_487),
.Y(n_525)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_525),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_508),
.A2(n_483),
.B1(n_501),
.B2(n_494),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_526),
.B(n_539),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_542),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_529),
.B(n_537),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_514),
.A2(n_499),
.B(n_500),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_530),
.A2(n_517),
.B(n_522),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_492),
.Y(n_531)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_531),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_488),
.Y(n_534)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_534),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_513),
.A2(n_497),
.B1(n_498),
.B2(n_405),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g541 ( 
.A1(n_502),
.A2(n_274),
.B1(n_300),
.B2(n_303),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_541),
.B(n_515),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_518),
.A2(n_274),
.B1(n_521),
.B2(n_523),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_532),
.B(n_506),
.C(n_503),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_543),
.B(n_550),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_545),
.A2(n_530),
.B(n_538),
.Y(n_563)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_547),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_529),
.B(n_520),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_R g554 ( 
.A(n_540),
.B(n_518),
.C(n_515),
.Y(n_554)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_554),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_504),
.C(n_511),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_555),
.B(n_556),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_528),
.B(n_505),
.C(n_519),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_533),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_557),
.B(n_535),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_544),
.A2(n_536),
.B1(n_526),
.B2(n_538),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_559),
.A2(n_565),
.B1(n_568),
.B2(n_549),
.Y(n_578)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_560),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_546),
.B(n_527),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_561),
.B(n_567),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_563),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_556),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_546),
.B(n_542),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_554),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_505),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_569),
.A2(n_548),
.B(n_551),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_552),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_571),
.B(n_576),
.Y(n_583)
);

AO21x1_ASAP7_75t_L g572 ( 
.A1(n_566),
.A2(n_540),
.B(n_548),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_572),
.A2(n_539),
.B(n_519),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_574),
.A2(n_563),
.B(n_569),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_564),
.B(n_543),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_561),
.B(n_551),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_545),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_578),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_579),
.A2(n_583),
.B(n_580),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_570),
.B(n_562),
.Y(n_580)
);

AOI21xp33_ASAP7_75t_L g586 ( 
.A1(n_580),
.A2(n_573),
.B(n_572),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_550),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_582),
.B(n_584),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_585),
.A2(n_573),
.B(n_555),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_586),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_587),
.B(n_589),
.C(n_581),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_590),
.B(n_588),
.Y(n_592)
);

BUFx24_ASAP7_75t_SL g593 ( 
.A(n_592),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_591),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_594),
.B(n_535),
.Y(n_595)
);


endmodule