module fake_aes_11227_n_27 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NOR2xp33_ASAP7_75t_L g8 ( .A(n_6), .B(n_3), .Y(n_8) );
INVx1_ASAP7_75t_SL g9 ( .A(n_3), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_4), .Y(n_10) );
INVx2_ASAP7_75t_SL g11 ( .A(n_1), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_7), .B(n_5), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
AND2x6_ASAP7_75t_L g14 ( .A(n_4), .B(n_0), .Y(n_14) );
A2O1A1Ixp33_ASAP7_75t_L g15 ( .A1(n_10), .A2(n_1), .B(n_2), .C(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
OAI21x1_ASAP7_75t_L g17 ( .A1(n_12), .A2(n_2), .B(n_8), .Y(n_17) );
AOI21x1_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_14), .B(n_9), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_19), .B(n_9), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
OAI211xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_15), .B(n_20), .C(n_18), .Y(n_23) );
AOI221xp5_ASAP7_75t_SL g24 ( .A1(n_23), .A2(n_22), .B1(n_17), .B2(n_18), .C(n_14), .Y(n_24) );
INVx3_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_14), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_25), .B1(n_14), .B2(n_24), .Y(n_27) );
endmodule