module fake_jpeg_11517_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_42),
.B(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_3),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_55),
.B(n_64),
.Y(n_110)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_18),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

CKINVDCx9p33_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_61),
.Y(n_99)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_5),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_67),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_7),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_16),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_76),
.B(n_79),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_22),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_96),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_23),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_109),
.B1(n_50),
.B2(n_52),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_22),
.B1(n_39),
.B2(n_25),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_66),
.B1(n_71),
.B2(n_63),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_22),
.B1(n_39),
.B2(n_24),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_91),
.B1(n_104),
.B2(n_59),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_39),
.B1(n_27),
.B2(n_25),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_18),
.B(n_37),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_105),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_27),
.B1(n_37),
.B2(n_23),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_28),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_21),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_80),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_57),
.A2(n_28),
.B1(n_16),
.B2(n_11),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_53),
.B(n_16),
.C(n_9),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_110),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_9),
.Y(n_113)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_114),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_48),
.A2(n_10),
.B(n_16),
.C(n_62),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_103),
.B1(n_121),
.B2(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_140),
.B1(n_149),
.B2(n_103),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_52),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_95),
.C(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_10),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_127),
.Y(n_152)
);

NOR2x1_ASAP7_75t_R g125 ( 
.A(n_100),
.B(n_63),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_125),
.A2(n_143),
.B(n_131),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_10),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_139),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_79),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

BUFx4f_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_136),
.B1(n_116),
.B2(n_146),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_88),
.A2(n_93),
.B1(n_81),
.B2(n_102),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_107),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_109),
.B1(n_102),
.B2(n_84),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_148),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_94),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_81),
.B(n_84),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_82),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_86),
.A2(n_95),
.B1(n_90),
.B2(n_85),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_97),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_125),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_165),
.B1(n_170),
.B2(n_136),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_122),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_174),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_132),
.B1(n_164),
.B2(n_174),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_131),
.B1(n_139),
.B2(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_176),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_122),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_130),
.B(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_123),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_126),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_189),
.Y(n_211)
);

AOI221xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_201),
.B1(n_178),
.B2(n_171),
.C(n_166),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_186),
.B(n_177),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_131),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_194),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_143),
.B(n_129),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_188),
.A2(n_186),
.B(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_129),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_198),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_150),
.B1(n_119),
.B2(n_118),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_195),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_180),
.B1(n_167),
.B2(n_179),
.Y(n_205)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_132),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_199),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_168),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_159),
.A2(n_157),
.B1(n_155),
.B2(n_153),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_190),
.A2(n_158),
.B(n_179),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_212),
.B(n_216),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_210),
.B(n_188),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_209),
.B1(n_191),
.B2(n_199),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_184),
.A2(n_166),
.B1(n_171),
.B2(n_161),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_181),
.B(n_198),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_161),
.B(n_168),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_177),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_201),
.C(n_197),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_196),
.Y(n_218)
);

AO221x1_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_212),
.B1(n_216),
.B2(n_207),
.C(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_207),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_213),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_195),
.B1(n_187),
.B2(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_202),
.A2(n_188),
.B(n_200),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_227),
.B(n_230),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_204),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_222),
.B(n_182),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_218),
.C(n_211),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_215),
.C(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_227),
.C(n_215),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_228),
.A3(n_224),
.B1(n_230),
.B2(n_229),
.C1(n_219),
.C2(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_239),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_220),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_245),
.A2(n_232),
.B(n_221),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_203),
.B(n_213),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_246),
.A2(n_232),
.B(n_235),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_185),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_250),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_220),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_209),
.C(n_205),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_249),
.A2(n_242),
.B(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_256),
.C(n_250),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_260),
.C(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_197),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_259),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_225),
.B(n_193),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_262),
.Y(n_264)
);


endmodule