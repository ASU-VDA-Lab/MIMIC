module real_aes_7771_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g519 ( .A1(n_0), .A2(n_165), .B(n_520), .C(n_523), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_1), .B(n_515), .Y(n_524) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_93), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g463 ( .A(n_2), .Y(n_463) );
INVx1_ASAP7_75t_L g163 ( .A(n_3), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_4), .B(n_166), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_5), .A2(n_484), .B(n_559), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_6), .A2(n_768), .B1(n_771), .B2(n_772), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_6), .Y(n_772) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_7), .A2(n_173), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_8), .A2(n_38), .B1(n_153), .B2(n_201), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_9), .B(n_173), .Y(n_181) );
AND2x6_ASAP7_75t_L g168 ( .A(n_10), .B(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_11), .A2(n_168), .B(n_489), .C(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_12), .A2(n_42), .B1(n_769), .B2(n_770), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_12), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_13), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_13), .B(n_39), .Y(n_464) );
INVx1_ASAP7_75t_L g147 ( .A(n_14), .Y(n_147) );
INVx1_ASAP7_75t_L g144 ( .A(n_15), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_16), .B(n_149), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_17), .B(n_166), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_18), .B(n_140), .Y(n_247) );
AO32x2_ASAP7_75t_L g217 ( .A1(n_19), .A2(n_139), .A3(n_173), .B1(n_192), .B2(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_20), .B(n_153), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_21), .B(n_140), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_22), .A2(n_58), .B1(n_153), .B2(n_201), .Y(n_220) );
AOI22xp33_ASAP7_75t_SL g203 ( .A1(n_23), .A2(n_85), .B1(n_149), .B2(n_153), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_24), .B(n_153), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_25), .A2(n_192), .B(n_489), .C(n_507), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_26), .A2(n_192), .B(n_489), .C(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_27), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_28), .B(n_194), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_29), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_29), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_30), .A2(n_484), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_31), .B(n_194), .Y(n_235) );
INVx2_ASAP7_75t_L g151 ( .A(n_32), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_33), .A2(n_487), .B(n_491), .C(n_497), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_34), .B(n_153), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_35), .A2(n_106), .B1(n_114), .B2(n_782), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_36), .B(n_194), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_37), .B(n_212), .Y(n_542) );
INVx1_ASAP7_75t_L g109 ( .A(n_39), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_40), .B(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_41), .Y(n_536) );
INVx1_ASAP7_75t_L g770 ( .A(n_42), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_43), .B(n_166), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_44), .A2(n_451), .B1(n_454), .B2(n_455), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_44), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_45), .B(n_484), .Y(n_539) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_46), .A2(n_48), .B1(n_452), .B2(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_46), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_46), .A2(n_127), .B1(n_128), .B2(n_453), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_47), .A2(n_487), .B(n_497), .C(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_48), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_49), .B(n_153), .Y(n_176) );
INVx1_ASAP7_75t_L g521 ( .A(n_50), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_51), .A2(n_94), .B1(n_201), .B2(n_202), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_52), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_53), .B(n_153), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_54), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g552 ( .A(n_55), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_56), .B(n_484), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_57), .B(n_161), .Y(n_180) );
AOI22xp33_ASAP7_75t_SL g245 ( .A1(n_59), .A2(n_63), .B1(n_149), .B2(n_153), .Y(n_245) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_60), .A2(n_70), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_60), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_61), .B(n_153), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_62), .B(n_153), .Y(n_209) );
INVx1_ASAP7_75t_L g169 ( .A(n_64), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_65), .B(n_484), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_66), .B(n_515), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_67), .A2(n_155), .B(n_161), .C(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_68), .B(n_153), .Y(n_164) );
INVx1_ASAP7_75t_L g143 ( .A(n_69), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_70), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_71), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_72), .B(n_166), .Y(n_495) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_73), .A2(n_173), .A3(n_192), .B1(n_199), .B2(n_204), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_74), .B(n_167), .Y(n_533) );
INVx1_ASAP7_75t_L g188 ( .A(n_75), .Y(n_188) );
INVx1_ASAP7_75t_L g230 ( .A(n_76), .Y(n_230) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_77), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_78), .B(n_494), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_79), .A2(n_489), .B(n_497), .C(n_586), .Y(n_585) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_80), .A2(n_470), .B1(n_763), .B2(n_764), .C1(n_773), .C2(n_777), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_81), .B(n_149), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g560 ( .A(n_82), .Y(n_560) );
INVx1_ASAP7_75t_L g113 ( .A(n_83), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_84), .B(n_493), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_86), .B(n_201), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_87), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_88), .B(n_149), .Y(n_234) );
INVx2_ASAP7_75t_L g141 ( .A(n_89), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_90), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_91), .B(n_191), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_92), .B(n_149), .Y(n_177) );
OR2x2_ASAP7_75t_L g460 ( .A(n_93), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g474 ( .A(n_93), .B(n_462), .Y(n_474) );
INVx2_ASAP7_75t_L g762 ( .A(n_93), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_95), .A2(n_104), .B1(n_149), .B2(n_150), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_96), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g492 ( .A(n_97), .Y(n_492) );
INVxp67_ASAP7_75t_L g563 ( .A(n_98), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_99), .B(n_149), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g529 ( .A(n_101), .Y(n_529) );
INVx1_ASAP7_75t_L g587 ( .A(n_102), .Y(n_587) );
AND2x2_ASAP7_75t_L g554 ( .A(n_103), .B(n_194), .Y(n_554) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx6p67_ASAP7_75t_R g783 ( .A(n_107), .Y(n_783) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_468), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g781 ( .A(n_118), .Y(n_781) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_457), .B(n_465), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_126), .B2(n_456), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_122), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_123), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_128), .B1(n_449), .B2(n_450), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_415), .Y(n_128) );
NOR3xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_319), .C(n_403), .Y(n_129) );
NAND4xp25_ASAP7_75t_L g130 ( .A(n_131), .B(n_262), .C(n_284), .D(n_300), .Y(n_130) );
AOI221xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_195), .B1(n_221), .B2(n_240), .C(n_248), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_171), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_134), .B(n_240), .Y(n_274) );
NAND4xp25_ASAP7_75t_L g314 ( .A(n_134), .B(n_302), .C(n_315), .D(n_317), .Y(n_314) );
INVxp67_ASAP7_75t_L g431 ( .A(n_134), .Y(n_431) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g313 ( .A(n_135), .B(n_251), .Y(n_313) );
AND2x2_ASAP7_75t_L g337 ( .A(n_135), .B(n_171), .Y(n_337) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g304 ( .A(n_136), .B(n_239), .Y(n_304) );
AND2x2_ASAP7_75t_L g344 ( .A(n_136), .B(n_325), .Y(n_344) );
AND2x2_ASAP7_75t_L g361 ( .A(n_136), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_136), .B(n_172), .Y(n_385) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g238 ( .A(n_137), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g256 ( .A(n_137), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g268 ( .A(n_137), .B(n_172), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_137), .B(n_182), .Y(n_290) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_145), .B(n_170), .Y(n_137) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_138), .A2(n_183), .B(n_193), .Y(n_182) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_139), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_141), .B(n_142), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_159), .B(n_168), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_152), .C(n_155), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_148), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_148), .A2(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx1_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
INVx3_ASAP7_75t_L g229 ( .A(n_153), .Y(n_229) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_153), .Y(n_589) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g201 ( .A(n_154), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
AND2x6_ASAP7_75t_L g489 ( .A(n_154), .B(n_490), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_155), .A2(n_587), .B(n_588), .C(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_156), .A2(n_233), .B(n_234), .Y(n_232) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g494 ( .A(n_157), .Y(n_494) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx3_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx1_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
AND2x2_ASAP7_75t_L g485 ( .A(n_158), .B(n_162), .Y(n_485) );
INVx1_ASAP7_75t_L g490 ( .A(n_158), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_163), .B(n_164), .C(n_165), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_L g187 ( .A1(n_160), .A2(n_188), .B(n_189), .C(n_190), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_160), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_165), .A2(n_179), .B(n_180), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_191), .B1(n_219), .B2(n_220), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_165), .A2(n_191), .B1(n_244), .B2(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_166), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_166), .A2(n_185), .B(n_186), .Y(n_184) );
O2A1O1Ixp5_ASAP7_75t_SL g228 ( .A1(n_166), .A2(n_229), .B(n_230), .C(n_231), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_166), .B(n_563), .Y(n_562) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g199 ( .A1(n_167), .A2(n_191), .B1(n_200), .B2(n_203), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_168), .A2(n_175), .B(n_178), .Y(n_174) );
BUFx3_ASAP7_75t_L g192 ( .A(n_168), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_168), .A2(n_208), .B(n_213), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_168), .A2(n_228), .B(n_232), .Y(n_227) );
AND2x4_ASAP7_75t_L g484 ( .A(n_168), .B(n_485), .Y(n_484) );
INVx4_ASAP7_75t_SL g498 ( .A(n_168), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_168), .B(n_485), .Y(n_530) );
AND2x2_ASAP7_75t_L g271 ( .A(n_171), .B(n_272), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_171), .A2(n_321), .B1(n_324), .B2(n_326), .C(n_330), .Y(n_320) );
AND2x2_ASAP7_75t_L g379 ( .A(n_171), .B(n_344), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_171), .B(n_361), .Y(n_413) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_182), .Y(n_171) );
INVx3_ASAP7_75t_L g239 ( .A(n_172), .Y(n_239) );
AND2x2_ASAP7_75t_L g288 ( .A(n_172), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g342 ( .A(n_172), .B(n_257), .Y(n_342) );
AND2x2_ASAP7_75t_L g400 ( .A(n_172), .B(n_401), .Y(n_400) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_181), .Y(n_172) );
INVx4_ASAP7_75t_L g242 ( .A(n_173), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_173), .A2(n_539), .B(n_540), .Y(n_538) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_173), .Y(n_557) );
AND2x2_ASAP7_75t_L g240 ( .A(n_182), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g257 ( .A(n_182), .Y(n_257) );
INVx1_ASAP7_75t_L g312 ( .A(n_182), .Y(n_312) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_182), .Y(n_318) );
AND2x2_ASAP7_75t_L g363 ( .A(n_182), .B(n_239), .Y(n_363) );
OR2x2_ASAP7_75t_L g402 ( .A(n_182), .B(n_241), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_187), .B(n_192), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_190), .A2(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx4_ASAP7_75t_L g522 ( .A(n_191), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g261 ( .A(n_192), .B(n_242), .C(n_243), .Y(n_261) );
INVx2_ASAP7_75t_L g204 ( .A(n_194), .Y(n_204) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_194), .A2(n_207), .B(n_216), .Y(n_206) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_194), .A2(n_227), .B(n_235), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_194), .A2(n_483), .B(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g512 ( .A(n_194), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_194), .A2(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_195), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
AND2x2_ASAP7_75t_L g398 ( .A(n_196), .B(n_395), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_196), .B(n_380), .Y(n_430) );
BUFx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g329 ( .A(n_197), .B(n_253), .Y(n_329) );
AND2x2_ASAP7_75t_L g378 ( .A(n_197), .B(n_224), .Y(n_378) );
INVx1_ASAP7_75t_L g424 ( .A(n_197), .Y(n_424) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
AND2x2_ASAP7_75t_L g279 ( .A(n_198), .B(n_253), .Y(n_279) );
INVx1_ASAP7_75t_L g296 ( .A(n_198), .Y(n_296) );
AND2x2_ASAP7_75t_L g302 ( .A(n_198), .B(n_217), .Y(n_302) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_202), .Y(n_496) );
INVx2_ASAP7_75t_L g523 ( .A(n_202), .Y(n_523) );
INVx1_ASAP7_75t_L g510 ( .A(n_204), .Y(n_510) );
AND2x2_ASAP7_75t_L g370 ( .A(n_205), .B(n_278), .Y(n_370) );
INVx2_ASAP7_75t_L g435 ( .A(n_205), .Y(n_435) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_217), .Y(n_205) );
AND2x2_ASAP7_75t_L g252 ( .A(n_206), .B(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g265 ( .A(n_206), .B(n_225), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_206), .B(n_224), .Y(n_293) );
INVx1_ASAP7_75t_L g299 ( .A(n_206), .Y(n_299) );
INVx1_ASAP7_75t_L g316 ( .A(n_206), .Y(n_316) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_206), .Y(n_328) );
INVx2_ASAP7_75t_L g396 ( .A(n_206), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g253 ( .A(n_217), .Y(n_253) );
BUFx2_ASAP7_75t_L g350 ( .A(n_217), .Y(n_350) );
AND2x2_ASAP7_75t_L g395 ( .A(n_217), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_223), .B(n_332), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_223), .A2(n_394), .B(n_408), .Y(n_418) );
AND2x2_ASAP7_75t_L g443 ( .A(n_223), .B(n_329), .Y(n_443) );
BUFx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g365 ( .A(n_225), .Y(n_365) );
AND2x2_ASAP7_75t_L g394 ( .A(n_225), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_226), .Y(n_278) );
INVx2_ASAP7_75t_L g297 ( .A(n_226), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_226), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g251 ( .A(n_237), .Y(n_251) );
OR2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g332 ( .A(n_237), .B(n_328), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_237), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g433 ( .A(n_237), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_237), .B(n_370), .Y(n_445) );
AND2x2_ASAP7_75t_L g324 ( .A(n_238), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g347 ( .A(n_238), .B(n_240), .Y(n_347) );
INVx2_ASAP7_75t_L g259 ( .A(n_239), .Y(n_259) );
AND2x2_ASAP7_75t_L g287 ( .A(n_239), .B(n_260), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_239), .B(n_312), .Y(n_368) );
AND2x2_ASAP7_75t_L g282 ( .A(n_240), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g429 ( .A(n_240), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_240), .B(n_304), .Y(n_441) );
AND2x2_ASAP7_75t_L g267 ( .A(n_241), .B(n_257), .Y(n_267) );
INVx1_ASAP7_75t_L g362 ( .A(n_241), .Y(n_362) );
AO21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_246), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_242), .B(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g515 ( .A(n_242), .Y(n_515) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_242), .A2(n_528), .B(n_535), .Y(n_527) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_242), .A2(n_584), .B(n_591), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_242), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g260 ( .A(n_247), .B(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_251), .B(n_298), .Y(n_307) );
OR2x2_ASAP7_75t_L g439 ( .A(n_251), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g356 ( .A(n_252), .B(n_297), .Y(n_356) );
AND2x2_ASAP7_75t_L g364 ( .A(n_252), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g423 ( .A(n_252), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g447 ( .A(n_252), .B(n_294), .Y(n_447) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_253), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g434 ( .A(n_253), .B(n_297), .Y(n_434) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
AND2x2_ASAP7_75t_L g286 ( .A(n_256), .B(n_287), .Y(n_286) );
INVxp67_ASAP7_75t_L g448 ( .A(n_256), .Y(n_448) );
NOR2x1_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g283 ( .A(n_259), .Y(n_283) );
AND2x2_ASAP7_75t_L g334 ( .A(n_259), .B(n_267), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_259), .B(n_402), .Y(n_428) );
INVx2_ASAP7_75t_L g273 ( .A(n_260), .Y(n_273) );
INVx3_ASAP7_75t_L g325 ( .A(n_260), .Y(n_325) );
OR2x2_ASAP7_75t_L g353 ( .A(n_260), .B(n_354), .Y(n_353) );
AOI311xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .A3(n_268), .B(n_269), .C(n_280), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_263), .A2(n_301), .B(n_303), .C(n_305), .Y(n_300) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_SL g285 ( .A(n_265), .Y(n_285) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g303 ( .A(n_267), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_267), .B(n_283), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_267), .B(n_268), .Y(n_436) );
AND2x2_ASAP7_75t_L g358 ( .A(n_268), .B(n_272), .Y(n_358) );
AOI21xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .B(n_275), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g416 ( .A(n_272), .B(n_304), .Y(n_416) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_273), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g310 ( .A(n_273), .Y(n_310) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
AND2x2_ASAP7_75t_L g301 ( .A(n_277), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g346 ( .A(n_279), .Y(n_346) );
AND2x4_ASAP7_75t_L g408 ( .A(n_279), .B(n_377), .Y(n_408) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_282), .A2(n_348), .B1(n_360), .B2(n_364), .C1(n_366), .C2(n_370), .Y(n_359) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_288), .C(n_291), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_285), .B(n_329), .Y(n_352) );
INVx1_ASAP7_75t_L g374 ( .A(n_287), .Y(n_374) );
INVx1_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
OR2x2_ASAP7_75t_L g373 ( .A(n_290), .B(n_374), .Y(n_373) );
OAI21xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_294), .B(n_298), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_292), .B(n_310), .C(n_311), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_292), .A2(n_329), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_296), .Y(n_349) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_297), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g406 ( .A(n_297), .Y(n_406) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_297), .Y(n_422) );
INVx2_ASAP7_75t_L g380 ( .A(n_298), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_302), .B(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g354 ( .A(n_304), .Y(n_354) );
OAI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B1(n_309), .B2(n_313), .C(n_314), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_308), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g442 ( .A(n_308), .Y(n_442) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g323 ( .A(n_315), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_315), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g381 ( .A(n_315), .B(n_329), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_315), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g414 ( .A(n_315), .B(n_349), .Y(n_414) );
BUFx3_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND5xp2_ASAP7_75t_L g319 ( .A(n_320), .B(n_338), .C(n_359), .D(n_371), .E(n_386), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI32xp33_ASAP7_75t_L g411 ( .A1(n_323), .A2(n_350), .A3(n_366), .B1(n_412), .B2(n_414), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_325), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_SL g335 ( .A(n_329), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B1(n_335), .B2(n_336), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_345), .B1(n_347), .B2(n_348), .C(n_351), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g410 ( .A(n_342), .B(n_361), .Y(n_410) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_347), .A2(n_408), .B1(n_426), .B2(n_431), .C(n_432), .Y(n_425) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_L g391 ( .A(n_350), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_355), .B2(n_357), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g369 ( .A(n_361), .Y(n_369) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B1(n_379), .B2(n_380), .C1(n_381), .C2(n_382), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_380), .A2(n_427), .B1(n_429), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_397), .B(n_399), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g440 ( .A(n_395), .Y(n_440) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_407), .B(n_409), .C(n_411), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B(n_419), .C(n_444), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_416), .Y(n_420) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_425), .C(n_437), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B(n_436), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_451), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_460), .Y(n_467) );
NOR2x2_ASAP7_75t_L g779 ( .A(n_461), .B(n_762), .Y(n_779) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g761 ( .A(n_462), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_465), .B(n_469), .C(n_780), .Y(n_468) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_472), .B1(n_475), .B2(n_761), .Y(n_470) );
INVx1_ASAP7_75t_L g774 ( .A(n_471), .Y(n_774) );
OAI22x1_ASAP7_75t_SL g773 ( .A1(n_472), .A2(n_476), .B1(n_774), .B2(n_775), .Y(n_773) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR3x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_675), .C(n_718), .Y(n_476) );
NAND5xp2_ASAP7_75t_L g477 ( .A(n_478), .B(n_602), .C(n_632), .D(n_649), .E(n_664), .Y(n_477) );
AOI221xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_525), .B1(n_565), .B2(n_571), .C(n_575), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_501), .Y(n_479) );
OR2x2_ASAP7_75t_L g580 ( .A(n_480), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g619 ( .A(n_480), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g637 ( .A(n_480), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_480), .B(n_573), .Y(n_654) );
OR2x2_ASAP7_75t_L g666 ( .A(n_480), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_480), .B(n_625), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_480), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_480), .B(n_603), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_480), .B(n_611), .Y(n_717) );
AND2x2_ASAP7_75t_L g749 ( .A(n_480), .B(n_513), .Y(n_749) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_480), .Y(n_757) );
INVx5_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_481), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g577 ( .A(n_481), .B(n_555), .Y(n_577) );
BUFx2_ASAP7_75t_L g599 ( .A(n_481), .Y(n_599) );
AND2x2_ASAP7_75t_L g628 ( .A(n_481), .B(n_502), .Y(n_628) );
AND2x2_ASAP7_75t_L g683 ( .A(n_481), .B(n_581), .Y(n_683) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_499), .Y(n_481) );
BUFx2_ASAP7_75t_L g505 ( .A(n_484), .Y(n_505) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_488), .A2(n_498), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_488), .A2(n_498), .B(n_560), .C(n_561), .Y(n_559) );
INVx5_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_495), .C(n_496), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_493), .A2(n_496), .B(n_552), .C(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_501), .B(n_637), .Y(n_646) );
OAI32xp33_ASAP7_75t_L g660 ( .A1(n_501), .A2(n_596), .A3(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_501), .B(n_662), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_501), .B(n_580), .Y(n_703) );
INVx1_ASAP7_75t_SL g732 ( .A(n_501), .Y(n_732) );
NAND4xp25_ASAP7_75t_L g741 ( .A(n_501), .B(n_527), .C(n_683), .D(n_742), .Y(n_741) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_513), .Y(n_501) );
INVx5_ASAP7_75t_L g574 ( .A(n_502), .Y(n_574) );
AND2x2_ASAP7_75t_L g603 ( .A(n_502), .B(n_514), .Y(n_603) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_502), .Y(n_682) );
AND2x2_ASAP7_75t_L g752 ( .A(n_502), .B(n_699), .Y(n_752) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_511), .Y(n_502) );
AOI21xp5_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B(n_510), .Y(n_503) );
AND2x4_ASAP7_75t_L g625 ( .A(n_513), .B(n_574), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_513), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g659 ( .A(n_513), .B(n_581), .Y(n_659) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g573 ( .A(n_514), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g611 ( .A(n_514), .B(n_583), .Y(n_611) );
AND2x2_ASAP7_75t_L g620 ( .A(n_514), .B(n_582), .Y(n_620) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_524), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_525), .A2(n_689), .B1(n_691), .B2(n_693), .C1(n_696), .C2(n_697), .Y(n_688) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_544), .Y(n_525) );
AND2x2_ASAP7_75t_L g621 ( .A(n_526), .B(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_526), .B(n_599), .C(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
INVx5_ASAP7_75t_SL g570 ( .A(n_527), .Y(n_570) );
OAI322xp33_ASAP7_75t_L g575 ( .A1(n_527), .A2(n_576), .A3(n_578), .B1(n_579), .B2(n_593), .C1(n_596), .C2(n_598), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_527), .B(n_568), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_527), .B(n_556), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
INVx2_ASAP7_75t_L g568 ( .A(n_537), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_537), .B(n_546), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_544), .B(n_606), .Y(n_661) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g640 ( .A(n_545), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_555), .Y(n_545) );
OR2x2_ASAP7_75t_L g569 ( .A(n_546), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_546), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g608 ( .A(n_546), .B(n_556), .Y(n_608) );
AND2x2_ASAP7_75t_L g631 ( .A(n_546), .B(n_568), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_546), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_546), .B(n_606), .Y(n_647) );
AND2x2_ASAP7_75t_L g655 ( .A(n_546), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_546), .B(n_615), .Y(n_705) );
INVx5_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g595 ( .A(n_547), .B(n_570), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_547), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g622 ( .A(n_547), .B(n_556), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_547), .B(n_669), .Y(n_710) );
OR2x2_ASAP7_75t_L g726 ( .A(n_547), .B(n_670), .Y(n_726) );
AND2x2_ASAP7_75t_SL g733 ( .A(n_547), .B(n_687), .Y(n_733) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_547), .Y(n_740) );
OR2x6_ASAP7_75t_L g547 ( .A(n_548), .B(n_554), .Y(n_547) );
AND2x2_ASAP7_75t_L g594 ( .A(n_555), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g644 ( .A(n_555), .B(n_568), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_555), .B(n_570), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_555), .B(n_606), .Y(n_728) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_556), .B(n_570), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_556), .B(n_568), .Y(n_616) );
OR2x2_ASAP7_75t_L g670 ( .A(n_556), .B(n_568), .Y(n_670) );
AND2x2_ASAP7_75t_L g687 ( .A(n_556), .B(n_567), .Y(n_687) );
INVxp67_ASAP7_75t_L g709 ( .A(n_556), .Y(n_709) );
AND2x2_ASAP7_75t_L g736 ( .A(n_556), .B(n_606), .Y(n_736) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_556), .Y(n_743) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_564), .Y(n_556) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_567), .B(n_617), .Y(n_690) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g606 ( .A(n_568), .B(n_570), .Y(n_606) );
OR2x2_ASAP7_75t_L g673 ( .A(n_568), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g617 ( .A(n_569), .Y(n_617) );
OR2x2_ASAP7_75t_L g678 ( .A(n_569), .B(n_670), .Y(n_678) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g578 ( .A(n_573), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_573), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_574), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_574), .B(n_581), .Y(n_613) );
INVx2_ASAP7_75t_L g658 ( .A(n_574), .Y(n_658) );
AND2x2_ASAP7_75t_L g671 ( .A(n_574), .B(n_611), .Y(n_671) );
AND2x2_ASAP7_75t_L g696 ( .A(n_574), .B(n_620), .Y(n_696) );
INVx1_ASAP7_75t_L g648 ( .A(n_579), .Y(n_648) );
INVx2_ASAP7_75t_SL g635 ( .A(n_580), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_581), .Y(n_638) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_582), .Y(n_601) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g699 ( .A(n_583), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g668 ( .A(n_595), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g674 ( .A(n_595), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_595), .A2(n_677), .B1(n_679), .B2(n_684), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_595), .B(n_687), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_596), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g630 ( .A(n_597), .Y(n_630) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
OR2x2_ASAP7_75t_L g612 ( .A(n_599), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_599), .B(n_603), .Y(n_663) );
AND2x2_ASAP7_75t_L g686 ( .A(n_599), .B(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g662 ( .A(n_601), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_609), .C(n_623), .Y(n_602) );
INVx1_ASAP7_75t_L g626 ( .A(n_603), .Y(n_626) );
OAI221xp5_ASAP7_75t_SL g734 ( .A1(n_603), .A2(n_735), .B1(n_737), .B2(n_738), .C(n_741), .Y(n_734) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g753 ( .A(n_606), .Y(n_753) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g702 ( .A(n_608), .B(n_641), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B(n_614), .C(n_618), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OAI32xp33_ASAP7_75t_L g727 ( .A1(n_616), .A2(n_617), .A3(n_680), .B1(n_717), .B2(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g759 ( .A(n_619), .B(n_658), .Y(n_759) );
AND2x2_ASAP7_75t_L g706 ( .A(n_620), .B(n_658), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_620), .B(n_628), .Y(n_724) );
AOI31xp33_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_626), .A3(n_627), .B(n_629), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_625), .B(n_637), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_625), .B(n_635), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_625), .A2(n_655), .B1(n_745), .B2(n_748), .C(n_750), .Y(n_744) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g650 ( .A(n_630), .B(n_651), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_639), .B1(n_642), .B2(n_645), .C1(n_647), .C2(n_648), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g715 ( .A(n_634), .Y(n_715) );
INVx1_ASAP7_75t_L g737 ( .A(n_637), .Y(n_737) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_640), .A2(n_751), .B1(n_753), .B2(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g656 ( .A(n_641), .Y(n_656) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_655), .B2(n_657), .C(n_660), .Y(n_649) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g694 ( .A(n_652), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g746 ( .A(n_652), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g721 ( .A(n_657), .Y(n_721) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g685 ( .A(n_658), .Y(n_685) );
INVx1_ASAP7_75t_L g667 ( .A(n_659), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_662), .B(n_749), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_671), .B2(n_672), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g758 ( .A(n_671), .Y(n_758) );
INVxp33_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_673), .B(n_717), .Y(n_716) );
OAI32xp33_ASAP7_75t_L g707 ( .A1(n_674), .A2(n_708), .A3(n_709), .B1(n_710), .B2(n_711), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_688), .C(n_700), .D(n_712), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_683), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g693 ( .A(n_694), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_697), .A2(n_713), .B1(n_730), .B2(n_733), .C(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g748 ( .A(n_699), .B(n_749), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_704), .B2(n_706), .C(n_707), .Y(n_700) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_709), .B(n_740), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g718 ( .A(n_719), .B(n_729), .C(n_744), .D(n_755), .Y(n_718) );
O2A1O1Ixp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B(n_725), .C(n_727), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g760 ( .A(n_747), .Y(n_760) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .B(n_760), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g776 ( .A(n_761), .Y(n_776) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx14_ASAP7_75t_R g771 ( .A(n_768), .Y(n_771) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
endmodule