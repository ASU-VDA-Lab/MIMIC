module fake_jpeg_15181_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx12_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_30),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

NAND2x1p5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_20),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_46),
.B(n_48),
.Y(n_93)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_51),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_60),
.Y(n_87)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_67),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_23),
.B1(n_34),
.B2(n_33),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_33),
.B1(n_19),
.B2(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_35),
.Y(n_100)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_16),
.B(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_28),
.B1(n_17),
.B2(n_29),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_63),
.A2(n_40),
.B1(n_23),
.B2(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_71),
.B(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_34),
.B1(n_33),
.B2(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_18),
.B1(n_32),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_32),
.B1(n_38),
.B2(n_42),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_89),
.B1(n_95),
.B2(n_64),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_43),
.B(n_27),
.C(n_17),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_20),
.B(n_30),
.C(n_24),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_32),
.B1(n_26),
.B2(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_48),
.B(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_56),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_97),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_49),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_99),
.B1(n_68),
.B2(n_53),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_59),
.B1(n_21),
.B2(n_25),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_21),
.B1(n_25),
.B2(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_68),
.B1(n_58),
.B2(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_102),
.B(n_103),
.Y(n_137)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_22),
.CI(n_55),
.CON(n_103),
.SN(n_103)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_118),
.B1(n_89),
.B2(n_101),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_109),
.A2(n_77),
.B1(n_73),
.B2(n_101),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_111),
.B(n_112),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_81),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_30),
.A3(n_64),
.B1(n_20),
.B2(n_24),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_52),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_0),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_129),
.B(n_130),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_85),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_90),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_65),
.C(n_69),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_82),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_52),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_126),
.B(n_72),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_54),
.Y(n_160)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_20),
.B(n_2),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_1),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_131),
.A2(n_134),
.B(n_141),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_72),
.B(n_75),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_157),
.Y(n_185)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_88),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_88),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_151),
.B(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_153),
.Y(n_170)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AOI22x1_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_75),
.B1(n_80),
.B2(n_87),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_121),
.B1(n_114),
.B2(n_77),
.Y(n_195)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_158),
.Y(n_182)
);

XOR2x2_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_79),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_87),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_156),
.B1(n_134),
.B2(n_131),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_161),
.B1(n_102),
.B2(n_108),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_73),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_98),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_113),
.A2(n_92),
.B1(n_85),
.B2(n_47),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_169),
.B1(n_133),
.B2(n_154),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_103),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_165),
.A2(n_167),
.B(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_123),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_192),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_103),
.C(n_114),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_83),
.C(n_107),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_135),
.B(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_176),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

CKINVDCx12_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_180),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_SL g224 ( 
.A1(n_178),
.A2(n_195),
.B(n_1),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_115),
.B(n_126),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_187),
.B(n_188),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_129),
.B(n_130),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_137),
.A2(n_85),
.B(n_111),
.C(n_130),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_155),
.B1(n_141),
.B2(n_143),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_140),
.B1(n_149),
.B2(n_147),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_138),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_110),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_169),
.A2(n_153),
.B1(n_150),
.B2(n_121),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_197),
.A2(n_200),
.B1(n_206),
.B2(n_214),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_150),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_208),
.C(n_217),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_224),
.B1(n_164),
.B2(n_190),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_169),
.A2(n_146),
.B1(n_127),
.B2(n_112),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_216),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_120),
.B(n_107),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_171),
.B(n_166),
.Y(n_235)
);

NAND2x1_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_179),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_223),
.B(n_185),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_167),
.B(n_170),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_213),
.B(n_188),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_169),
.A2(n_74),
.B1(n_69),
.B2(n_54),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_185),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_69),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_174),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_13),
.C(n_12),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_192),
.C(n_187),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_179),
.A2(n_1),
.B(n_2),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_184),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_242),
.C(n_218),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_198),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_238),
.B1(n_247),
.B2(n_210),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_165),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_232),
.B(n_235),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_178),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_177),
.B(n_183),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_193),
.C(n_181),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_180),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_188),
.B(n_182),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_248),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_261),
.C(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_243),
.B1(n_232),
.B2(n_244),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_172),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_199),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_264),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_213),
.C(n_217),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_262),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_197),
.C(n_205),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_200),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_205),
.B1(n_220),
.B2(n_214),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_231),
.B1(n_259),
.B2(n_268),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_181),
.C(n_176),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_235),
.C(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_270),
.B(n_245),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_275),
.C(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_278),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_241),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_269),
.B(n_262),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_234),
.B1(n_237),
.B2(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_230),
.B1(n_240),
.B2(n_229),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_230),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_285),
.C(n_253),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_238),
.B(n_223),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_266),
.B1(n_193),
.B2(n_188),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_249),
.C(n_190),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_263),
.C(n_267),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_221),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_288),
.B(n_289),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_163),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_295),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_296),
.B1(n_274),
.B2(n_283),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_258),
.B(n_252),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_191),
.C(n_188),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_300),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_3),
.C(n_4),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_282),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_308),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_294),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_279),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_3),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_3),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_272),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_287),
.A3(n_296),
.B1(n_10),
.B2(n_11),
.C1(n_14),
.C2(n_12),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_14),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_3),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

NOR4xp25_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.C(n_302),
.D(n_5),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_4),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_319),
.C(n_307),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_4),
.C(n_5),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_310),
.B1(n_5),
.B2(n_6),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_4),
.B(n_5),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_6),
.B(n_7),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_320),
.C(n_321),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_326),
.B1(n_314),
.B2(n_327),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_315),
.B1(n_6),
.B2(n_8),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_8),
.Y(n_332)
);


endmodule