module real_jpeg_7224_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_0),
.A2(n_161),
.B1(n_165),
.B2(n_168),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_0),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_0),
.B(n_181),
.C(n_185),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_0),
.B(n_77),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_0),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_0),
.B(n_129),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_0),
.B(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_1),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_1),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_1),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_1),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_1),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_2),
.A2(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_2),
.A2(n_66),
.B1(n_213),
.B2(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_2),
.A2(n_66),
.B1(n_85),
.B2(n_221),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_2),
.A2(n_66),
.B1(n_380),
.B2(n_457),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_3),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_102),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_102),
.B1(n_139),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_3),
.A2(n_102),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_4),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_4),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_4),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_4),
.Y(n_370)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_4),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_4),
.Y(n_419)
);

BUFx5_ASAP7_75t_L g443 ( 
.A(n_4),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_5),
.A2(n_55),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_5),
.A2(n_55),
.B1(n_221),
.B2(n_405),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_5),
.A2(n_55),
.B1(n_297),
.B2(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_8),
.A2(n_192),
.B1(n_197),
.B2(n_198),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_8),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_8),
.A2(n_161),
.B1(n_197),
.B2(n_266),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_8),
.A2(n_197),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_8),
.A2(n_197),
.B1(n_418),
.B2(n_420),
.Y(n_417)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_9),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_172),
.B1(n_213),
.B2(n_216),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_11),
.A2(n_172),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_11),
.A2(n_172),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_13),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_13),
.Y(n_215)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_15),
.A2(n_90),
.B1(n_92),
.B2(n_96),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_15),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_15),
.A2(n_96),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_15),
.A2(n_96),
.B1(n_243),
.B2(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_15),
.A2(n_96),
.B1(n_384),
.B2(n_425),
.Y(n_424)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_17),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_17),
.A2(n_223),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_17),
.A2(n_223),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_17),
.A2(n_223),
.B1(n_442),
.B2(n_444),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_18),
.A2(n_285),
.B1(n_289),
.B2(n_290),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_18),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_18),
.A2(n_109),
.B1(n_289),
.B2(n_384),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_18),
.A2(n_289),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_L g469 ( 
.A1(n_18),
.A2(n_289),
.B1(n_364),
.B2(n_470),
.Y(n_469)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_545),
.B(n_548),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_150),
.B(n_544),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_143),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_27),
.B(n_143),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_134),
.C(n_140),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_28),
.A2(n_29),
.B1(n_540),
.B2(n_541),
.Y(n_539)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_67),
.C(n_103),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_30),
.B(n_532),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_31),
.A2(n_56),
.B1(n_58),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_31),
.A2(n_56),
.B1(n_135),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_31),
.A2(n_368),
.B(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_31),
.A2(n_44),
.B1(n_417),
.B2(n_441),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_31),
.A2(n_54),
.B1(n_56),
.B2(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_32),
.A2(n_363),
.B(n_367),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_32),
.B(n_369),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_32),
.A2(n_57),
.B(n_547),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_44),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_43),
.Y(n_345)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_44),
.B(n_168),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_44)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_45),
.Y(n_343)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g280 ( 
.A(n_47),
.Y(n_280)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_48),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_50),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_50),
.Y(n_348)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_50),
.Y(n_378)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_50),
.Y(n_381)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_51),
.Y(n_279)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_56),
.A2(n_441),
.B(n_471),
.Y(n_481)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_57),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_57),
.B(n_469),
.Y(n_468)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_61),
.Y(n_445)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_67),
.A2(n_103),
.B1(n_104),
.B2(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_67),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_89),
.B1(n_97),
.B2(n_98),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_68),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_68),
.A2(n_97),
.B1(n_315),
.B2(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_68),
.A2(n_97),
.B1(n_411),
.B2(n_414),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_68),
.A2(n_89),
.B1(n_97),
.B2(n_521),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_77),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_71),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_73),
.Y(n_412)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_74),
.Y(n_304)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_77),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

AOI22x1_ASAP7_75t_L g446 ( 
.A1(n_77),
.A2(n_141),
.B1(n_319),
.B2(n_447),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_77),
.A2(n_141),
.B1(n_455),
.B2(n_456),
.Y(n_454)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_85),
.B2(n_87),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_83),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_84),
.Y(n_298)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_84),
.Y(n_407)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_90),
.Y(n_272)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_97),
.B(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_97),
.A2(n_315),
.B(n_318),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_99),
.Y(n_413)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_103),
.A2(n_104),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_103),
.B(n_516),
.C(n_519),
.Y(n_527)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_128),
.B(n_130),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_105),
.A2(n_160),
.B(n_169),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_105),
.A2(n_128),
.B1(n_220),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_105),
.A2(n_169),
.B(n_265),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_105),
.A2(n_128),
.B1(n_383),
.B2(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_106),
.B(n_170),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_106),
.A2(n_129),
.B1(n_404),
.B2(n_408),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_106),
.A2(n_129),
.B1(n_408),
.B2(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_106),
.A2(n_129),
.B1(n_424),
.B2(n_460),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_110),
.Y(n_225)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_117),
.A2(n_220),
.B(n_226),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_124),
.B2(n_126),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_122),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_125),
.Y(n_244)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_125),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_125),
.Y(n_400)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_128),
.A2(n_226),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_130),
.Y(n_460)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_134),
.B(n_140),
.Y(n_541)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_141),
.A2(n_271),
.B(n_277),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_141),
.B(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_141),
.A2(n_277),
.B(n_484),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_143),
.B(n_546),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_143),
.B(n_546),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_144),
.Y(n_547)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_147),
.B(n_168),
.Y(n_349)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_538),
.B(n_543),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_510),
.B(n_535),
.Y(n_151)
);

OAI311xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_388),
.A3(n_486),
.B1(n_504),
.C1(n_505),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_333),
.B(n_387),
.Y(n_153)
);

AO21x1_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_306),
.B(n_332),
.Y(n_154)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_259),
.B(n_305),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_229),
.B(n_258),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_189),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_158),
.B(n_189),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_175),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_159),
.A2(n_175),
.B1(n_176),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_159),
.Y(n_256)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx5_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g385 ( 
.A(n_167),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_168),
.A2(n_201),
.B(n_209),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_SL g271 ( 
.A1(n_168),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_SL g363 ( 
.A1(n_168),
.A2(n_349),
.B(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_188),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_217),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_190),
.B(n_218),
.C(n_228),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_201),
.B(n_209),
.Y(n_190)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_196),
.Y(n_397)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_200),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_201),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_201),
.A2(n_394),
.B1(n_398),
.B2(n_399),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_201),
.A2(n_399),
.B(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_212),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_202),
.A2(n_210),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_202),
.A2(n_284),
.B1(n_323),
.B2(n_329),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_202),
.A2(n_355),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_205),
.Y(n_330)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_205),
.Y(n_438)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_215),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_227),
.B2(n_228),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g302 ( 
.A(n_224),
.B(n_303),
.Y(n_302)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_251),
.B(n_257),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_239),
.B(n_250),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_235),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_237),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_249),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_249),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_248),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_248),
.A2(n_283),
.B(n_293),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_261),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_281),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_269),
.B2(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_269),
.C(n_281),
.Y(n_307)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI32xp33_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_297),
.A3(n_298),
.B1(n_299),
.B2(n_302),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_296),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_307),
.B(n_308),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_313),
.B2(n_331),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_312),
.C(n_331),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_313),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_321),
.C(n_322),
.Y(n_357)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_317),
.A2(n_340),
.A3(n_342),
.B1(n_344),
.B2(n_349),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_323),
.Y(n_352)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_334),
.B(n_335),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_360),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_336)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_350),
.B2(n_351),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_339),
.B(n_350),
.Y(n_482)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_347),
.Y(n_346)
);

INVx6_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_357),
.B(n_358),
.C(n_360),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_374),
.B2(n_386),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_361),
.B(n_375),
.C(n_382),
.Y(n_495)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_366),
.Y(n_470)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_373),
.Y(n_420)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_382),
.Y(n_374)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_376),
.Y(n_484)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_377),
.Y(n_457)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_472),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_SL g505 ( 
.A1(n_389),
.A2(n_472),
.B(n_506),
.C(n_509),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_448),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_390),
.B(n_448),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_421),
.C(n_431),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_391),
.B(n_421),
.CI(n_431),
.CON(n_485),
.SN(n_485)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_409),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_392),
.B(n_410),
.C(n_416),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_403),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_393),
.B(n_403),
.Y(n_478)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

INVx4_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_422),
.A2(n_423),
.B1(n_427),
.B2(n_430),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_423),
.B(n_427),
.Y(n_464)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_427),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_427),
.A2(n_430),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_427),
.A2(n_464),
.B(n_467),
.Y(n_513)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.C(n_446),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_432),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_433),
.B(n_435),
.Y(n_494)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_439),
.A2(n_440),
.B1(n_446),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_446),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_449),
.B(n_452),
.C(n_462),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_462),
.B2(n_463),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_458),
.B(n_461),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_459),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_456),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

FAx1_ASAP7_75t_SL g512 ( 
.A(n_461),
.B(n_513),
.CI(n_514),
.CON(n_512),
.SN(n_512)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_461),
.B(n_513),
.C(n_514),
.Y(n_534)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_471),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_485),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_485),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_478),
.C(n_479),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_474),
.A2(n_475),
.B1(n_478),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_478),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_482),
.C(n_483),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_480),
.A2(n_481),
.B1(n_483),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_483),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g551 ( 
.A(n_485),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_499),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_488),
.A2(n_507),
.B(n_508),
.Y(n_506)
);

NOR2x1_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_496),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_496),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.C(n_495),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_502),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_493),
.A2(n_494),
.B1(n_495),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_495),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_501),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_524),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_512),
.B(n_523),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_512),
.B(n_523),
.Y(n_536)
);

BUFx24_ASAP7_75t_SL g552 ( 
.A(n_512),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_516),
.B1(n_518),
.B2(n_522),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_515),
.A2(n_516),
.B1(n_530),
.B2(n_531),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_515),
.B(n_526),
.C(n_530),
.Y(n_542)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_518),
.Y(n_522)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_524),
.A2(n_536),
.B(n_537),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_525),
.B(n_534),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_534),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_527),
.B1(n_528),
.B2(n_529),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_542),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_539),
.B(n_542),
.Y(n_543)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);


endmodule