module fake_jpeg_14753_n_173 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_32),
.Y(n_51)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_14),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_32),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_26),
.B1(n_17),
.B2(n_19),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_50),
.B1(n_30),
.B2(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_29),
.A2(n_17),
.B1(n_14),
.B2(n_19),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_35),
.B1(n_17),
.B2(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_66),
.B1(n_48),
.B2(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_27),
.C(n_34),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_34),
.C(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_45),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_18),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_18),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_79),
.C(n_27),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_31),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_63),
.B(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_48),
.B1(n_43),
.B2(n_37),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_27),
.C(n_34),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_83),
.B(n_89),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_0),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_84),
.B(n_85),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_39),
.B1(n_37),
.B2(n_64),
.Y(n_86)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_48),
.B(n_43),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_53),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_66),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_20),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_53),
.C(n_75),
.Y(n_100)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_13),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_92),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_86),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_103),
.B(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_105),
.C(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_67),
.B1(n_88),
.B2(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_67),
.B1(n_40),
.B2(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_74),
.B1(n_75),
.B2(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_74),
.B1(n_76),
.B2(n_28),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_19),
.B1(n_15),
.B2(n_13),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

OAI321xp33_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_82),
.A3(n_94),
.B1(n_28),
.B2(n_23),
.C(n_24),
.Y(n_115)
);

OAI21x1_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_120),
.B(n_23),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_21),
.B(n_20),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_118),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_123),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_21),
.B(n_15),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_124),
.C(n_65),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_111),
.B(n_16),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_16),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_65),
.C(n_27),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_132),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_102),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_16),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_131),
.B1(n_133),
.B2(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_97),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_103),
.B1(n_1),
.B2(n_2),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_125),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_124),
.C(n_121),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_118),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_147),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_24),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_145),
.B(n_23),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_24),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_131),
.B1(n_130),
.B2(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_128),
.B(n_3),
.Y(n_149)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_155),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_0),
.B(n_4),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_5),
.B(n_7),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_22),
.C(n_5),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_143),
.A3(n_142),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_153),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_153),
.B(n_154),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_164),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_160),
.B(n_7),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_8),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_159),
.C(n_158),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_168),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.C1(n_159),
.C2(n_152),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_164),
.B(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.C(n_167),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_11),
.Y(n_173)
);


endmodule