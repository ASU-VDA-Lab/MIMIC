module fake_jpeg_22263_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_30),
.Y(n_48)
);

NAND3xp33_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_14),
.C(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_19),
.B1(n_14),
.B2(n_20),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_14),
.B1(n_21),
.B2(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_37),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_37),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_27),
.B(n_19),
.C(n_25),
.Y(n_92)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_62),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_35),
.B1(n_32),
.B2(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_18),
.B1(n_16),
.B2(n_21),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_69),
.B1(n_34),
.B2(n_29),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_19),
.B1(n_32),
.B2(n_14),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_48),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_32),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_56),
.Y(n_118)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_83),
.B1(n_88),
.B2(n_100),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_13),
.C(n_12),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_84),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_47),
.B1(n_46),
.B2(n_55),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_46),
.B1(n_48),
.B2(n_53),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_76),
.B(n_75),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_38),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_74),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_28),
.B1(n_21),
.B2(n_18),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_58),
.A2(n_39),
.B1(n_40),
.B2(n_18),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_110),
.B(n_113),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_99),
.B1(n_86),
.B2(n_93),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_59),
.Y(n_139)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_109),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_86),
.B1(n_93),
.B2(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_61),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_66),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_120),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_123),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_27),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_9),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_40),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_80),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_88),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_131),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_78),
.B1(n_59),
.B2(n_90),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_104),
.B1(n_124),
.B2(n_115),
.Y(n_159)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_151),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_150),
.B1(n_122),
.B2(n_104),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_71),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_68),
.B(n_64),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_148),
.B(n_16),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_111),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_16),
.B(n_18),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_71),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_94),
.B1(n_62),
.B2(n_70),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_68),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_123),
.B1(n_122),
.B2(n_106),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_153),
.A2(n_170),
.B1(n_144),
.B2(n_163),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_114),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_126),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_158),
.B(n_166),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_148),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_107),
.B1(n_115),
.B2(n_124),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_116),
.B1(n_111),
.B2(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_119),
.B1(n_63),
.B2(n_89),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_15),
.C(n_23),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_129),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_119),
.B1(n_22),
.B2(n_21),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_70),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_142),
.B(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_180),
.B(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_134),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_136),
.C(n_141),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_165),
.C(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_140),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_202),
.B1(n_162),
.B2(n_170),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_130),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_201),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_127),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_139),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_153),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_163),
.B1(n_155),
.B2(n_154),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_210),
.A2(n_220),
.B1(n_226),
.B2(n_198),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_166),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_182),
.C(n_190),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_179),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_222),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_198),
.B1(n_225),
.B2(n_190),
.Y(n_242)
);

A2O1A1O1Ixp25_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_196),
.B(n_201),
.C(n_152),
.D(n_154),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_192),
.C(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_219),
.C(n_221),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_165),
.C(n_161),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_133),
.B1(n_144),
.B2(n_161),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_156),
.C(n_138),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_203),
.B(n_176),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_156),
.C(n_150),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_205),
.C(n_222),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_137),
.B1(n_27),
.B2(n_28),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_232),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_186),
.Y(n_228)
);

AO22x1_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_241),
.B1(n_24),
.B2(n_13),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_229),
.B(n_243),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_188),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_44),
.Y(n_251)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_195),
.B(n_182),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_20),
.B(n_15),
.Y(n_249)
);

NOR2xp67_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_184),
.Y(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_244),
.B(n_246),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_221),
.B1(n_219),
.B2(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_204),
.C(n_26),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_214),
.A2(n_204),
.B1(n_89),
.B2(n_27),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_254),
.C(n_257),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_249),
.A2(n_23),
.B(n_22),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_228),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_247),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_10),
.B(n_13),
.C(n_11),
.D(n_8),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_44),
.C(n_64),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_236),
.C(n_231),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_44),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_263),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_11),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_253),
.B1(n_248),
.B2(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_230),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_231),
.C(n_68),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_16),
.C(n_28),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_264),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_11),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_276),
.C(n_254),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_15),
.C(n_26),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_8),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_26),
.B1(n_23),
.B2(n_20),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_279),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_292),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_273),
.B1(n_271),
.B2(n_265),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_287),
.B1(n_285),
.B2(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_252),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_250),
.B1(n_17),
.B2(n_22),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_25),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_25),
.C(n_56),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_1),
.C(n_2),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_25),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_277),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_8),
.B(n_53),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_298),
.B(n_302),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_284),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_3),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_284),
.A2(n_1),
.B(n_2),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_2),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_1),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_304),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_3),
.B(n_4),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.C(n_302),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_4),
.B(n_5),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_311),
.B(n_308),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_299),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_313),
.B(n_301),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_4),
.C(n_5),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_7),
.B(n_5),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_6),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_6),
.B(n_7),
.Y(n_318)
);


endmodule