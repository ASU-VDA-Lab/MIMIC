module fake_jpeg_11482_n_580 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_580);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_8),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_55),
.B(n_74),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_56),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_34),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_99),
.Y(n_125)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_8),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_73),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_10),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_7),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_83),
.B(n_44),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_89),
.Y(n_137)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_34),
.B(n_18),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_44),
.B(n_7),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_45),
.B1(n_38),
.B2(n_40),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_117),
.A2(n_120),
.B1(n_121),
.B2(n_136),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_55),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_29),
.B1(n_47),
.B2(n_42),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_58),
.A2(n_52),
.B1(n_29),
.B2(n_47),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_123),
.A2(n_149),
.B(n_174),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_132),
.B(n_148),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_74),
.A2(n_29),
.B1(n_51),
.B2(n_49),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_67),
.A2(n_29),
.B1(n_51),
.B2(n_49),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_142),
.A2(n_35),
.B1(n_27),
.B2(n_28),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_53),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_57),
.A2(n_42),
.B1(n_47),
.B2(n_41),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_57),
.B(n_21),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_158),
.B(n_168),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_21),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_54),
.A2(n_38),
.B1(n_47),
.B2(n_40),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_42),
.B1(n_41),
.B2(n_59),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_66),
.A2(n_41),
.B1(n_42),
.B2(n_40),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_56),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_182),
.Y(n_212)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_88),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_116),
.B(n_0),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_184),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_185),
.B(n_208),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_186),
.A2(n_187),
.B1(n_193),
.B2(n_198),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_82),
.B1(n_78),
.B2(n_71),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_189),
.Y(n_268)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_190),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_121),
.A2(n_94),
.B1(n_107),
.B2(n_103),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g250 ( 
.A1(n_191),
.A2(n_203),
.B1(n_209),
.B2(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_125),
.B(n_37),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_174),
.A2(n_86),
.B1(n_79),
.B2(n_102),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_116),
.B(n_0),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_217),
.Y(n_258)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVx3_ASAP7_75t_SL g270 ( 
.A(n_197),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_129),
.A2(n_113),
.B1(n_81),
.B2(n_96),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_114),
.A2(n_27),
.B1(n_46),
.B2(n_35),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_201),
.Y(n_293)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_202),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_92),
.B1(n_89),
.B2(n_84),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_119),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_128),
.A2(n_62),
.B1(n_64),
.B2(n_37),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_211),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_139),
.A2(n_31),
.B1(n_19),
.B2(n_46),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_213),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_151),
.A2(n_31),
.B1(n_19),
.B2(n_46),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_126),
.B(n_31),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_221),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_133),
.Y(n_216)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_154),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_218),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_130),
.A2(n_28),
.B1(n_19),
.B2(n_35),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_219),
.A2(n_238),
.B1(n_242),
.B2(n_244),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_123),
.A2(n_111),
.B1(n_27),
.B2(n_28),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_220),
.A2(n_232),
.B1(n_237),
.B2(n_240),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_223),
.A2(n_245),
.B1(n_162),
.B2(n_177),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_152),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_224),
.B(n_225),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_161),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_228),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_150),
.B(n_0),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_229),
.B(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_230),
.B(n_231),
.Y(n_283)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_179),
.A2(n_105),
.B1(n_87),
.B2(n_50),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_143),
.B(n_87),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_233),
.B(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_153),
.B(n_105),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_135),
.A2(n_112),
.B1(n_50),
.B2(n_3),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_236),
.A2(n_248),
.B(n_11),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_151),
.A2(n_1),
.B1(n_16),
.B2(n_3),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_137),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_137),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_240)
);

BUFx6f_ASAP7_75t_SL g241 ( 
.A(n_161),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g291 ( 
.A(n_241),
.Y(n_291)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_124),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_134),
.A2(n_1),
.B1(n_15),
.B2(n_5),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_134),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_145),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_246),
.A2(n_247),
.B1(n_156),
.B2(n_176),
.Y(n_295)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_131),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_146),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_266),
.Y(n_302)
);

OA22x2_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_131),
.B1(n_146),
.B2(n_141),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_SL g300 ( 
.A1(n_262),
.A2(n_243),
.B(n_193),
.C(n_187),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_184),
.B(n_147),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_217),
.C(n_248),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_192),
.B(n_164),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_245),
.B1(n_244),
.B2(n_237),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_234),
.B(n_164),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_275),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_234),
.B(n_140),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_184),
.B(n_194),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_194),
.B(n_162),
.Y(n_284)
);

AO22x1_ASAP7_75t_L g285 ( 
.A1(n_225),
.A2(n_167),
.B1(n_127),
.B2(n_178),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_285),
.A2(n_289),
.B(n_297),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_202),
.B(n_178),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_296),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_195),
.B(n_167),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_195),
.B(n_11),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_12),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_295),
.A2(n_299),
.B1(n_221),
.B2(n_241),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_215),
.B(n_176),
.Y(n_296)
);

NOR2x1_ASAP7_75t_R g297 ( 
.A(n_199),
.B(n_11),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_232),
.A2(n_172),
.B1(n_173),
.B2(n_177),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_300),
.A2(n_331),
.B1(n_262),
.B2(n_286),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_259),
.B(n_212),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_303),
.B(n_326),
.Y(n_354)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_287),
.Y(n_304)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_258),
.Y(n_344)
);

AO22x1_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_199),
.B1(n_223),
.B2(n_210),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_307),
.B(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_249),
.Y(n_309)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_310),
.A2(n_317),
.B1(n_278),
.B2(n_298),
.Y(n_345)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_236),
.B1(n_173),
.B2(n_229),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_313),
.A2(n_322),
.B1(n_335),
.B2(n_341),
.Y(n_357)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_269),
.A2(n_217),
.B1(n_228),
.B2(n_190),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_264),
.Y(n_318)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_283),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_323),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_211),
.C(n_185),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_258),
.C(n_281),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_292),
.A2(n_247),
.B1(n_246),
.B2(n_242),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_325),
.Y(n_365)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_256),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_231),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_277),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_330),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_230),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_262),
.A2(n_188),
.B1(n_216),
.B2(n_218),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_259),
.B(n_224),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_334),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_216),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_263),
.A2(n_205),
.B1(n_204),
.B2(n_189),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_275),
.B(n_196),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_337),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_260),
.A2(n_188),
.B(n_201),
.C(n_14),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_338),
.Y(n_374)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_339),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_273),
.B(n_239),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_340),
.A2(n_274),
.B(n_289),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_263),
.A2(n_197),
.B1(n_206),
.B2(n_207),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_342),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_364),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_345),
.A2(n_350),
.B1(n_372),
.B2(n_373),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_348),
.A2(n_319),
.B1(n_279),
.B2(n_257),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_310),
.A2(n_297),
.B1(n_262),
.B2(n_286),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_312),
.B(n_258),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_352),
.B(n_362),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_328),
.A2(n_290),
.B(n_285),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_353),
.A2(n_356),
.B(n_367),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_306),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_289),
.B(n_272),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_260),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_313),
.A2(n_250),
.B1(n_261),
.B2(n_281),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_363),
.A2(n_317),
.B1(n_307),
.B2(n_300),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_282),
.C(n_271),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_308),
.A2(n_284),
.B(n_253),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_328),
.A2(n_285),
.B(n_288),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_368),
.A2(n_375),
.B(n_378),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_304),
.A2(n_270),
.B1(n_253),
.B2(n_267),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_300),
.A2(n_270),
.B1(n_255),
.B2(n_257),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_316),
.A2(n_270),
.B1(n_251),
.B2(n_267),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_311),
.A2(n_279),
.B(n_251),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_379),
.Y(n_417)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_329),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_383),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_320),
.B(n_315),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_406),
.B(n_361),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_393),
.C(n_403),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_396),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_333),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_388),
.B(n_399),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_389),
.A2(n_398),
.B1(n_401),
.B2(n_409),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_302),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_341),
.B1(n_335),
.B2(n_322),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_394),
.A2(n_405),
.B1(n_410),
.B2(n_375),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_302),
.Y(n_395)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_360),
.B(n_333),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_359),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_397),
.B(n_402),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_370),
.A2(n_363),
.B1(n_357),
.B2(n_353),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_354),
.B(n_332),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_352),
.B(n_327),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_390),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_357),
.A2(n_300),
.B1(n_307),
.B2(n_336),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_360),
.B(n_330),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_340),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_359),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_374),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_345),
.A2(n_300),
.B1(n_309),
.B2(n_305),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_361),
.A2(n_334),
.B(n_338),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_346),
.B(n_339),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_407),
.B(n_408),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_347),
.A2(n_337),
.B1(n_325),
.B2(n_324),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_350),
.A2(n_323),
.B1(n_318),
.B2(n_314),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_349),
.Y(n_411)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_411),
.Y(n_424)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_358),
.Y(n_412)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_413),
.A2(n_372),
.B1(n_358),
.B2(n_351),
.Y(n_433)
);

MAJx2_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_364),
.C(n_352),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_388),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_407),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_429),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_418),
.B(n_390),
.Y(n_449)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_367),
.C(n_356),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_391),
.C(n_400),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_428),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_405),
.A2(n_347),
.B1(n_368),
.B2(n_366),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_383),
.A2(n_354),
.B1(n_369),
.B2(n_366),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_431),
.A2(n_433),
.B1(n_380),
.B2(n_404),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_386),
.B(n_326),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_434),
.B(n_437),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_391),
.A2(n_387),
.B(n_382),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_396),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_445),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_393),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_446),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_382),
.B(n_378),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_440),
.A2(n_410),
.B(n_411),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_381),
.A2(n_384),
.B(n_398),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_441),
.A2(n_442),
.B(n_409),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_381),
.A2(n_346),
.B(n_376),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_401),
.A2(n_376),
.B1(n_374),
.B2(n_377),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_443),
.A2(n_394),
.B1(n_389),
.B2(n_413),
.Y(n_463)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_387),
.A2(n_377),
.B1(n_351),
.B2(n_371),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_254),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_448),
.A2(n_419),
.B1(n_416),
.B2(n_429),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_453),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_470),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_395),
.C(n_406),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_456),
.C(n_465),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_444),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_464),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_414),
.B(n_397),
.C(n_402),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_458),
.A2(n_460),
.B(n_473),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_420),
.B(n_412),
.Y(n_459)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_426),
.B(n_371),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_461),
.B(n_474),
.Y(n_493)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_435),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_254),
.C(n_252),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_415),
.B(n_252),
.C(n_293),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_469),
.C(n_425),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_435),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_468),
.A2(n_427),
.B(n_438),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_423),
.B(n_268),
.C(n_293),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_268),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_432),
.A2(n_276),
.B1(n_291),
.B2(n_14),
.Y(n_472)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_441),
.A2(n_291),
.B(n_276),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_436),
.B(n_12),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_476),
.A2(n_464),
.B1(n_455),
.B2(n_462),
.Y(n_518)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_481),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_484),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_437),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_491),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_497),
.Y(n_513)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_488),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_447),
.A2(n_432),
.B1(n_443),
.B2(n_442),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_418),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_494),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_428),
.C(n_440),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_456),
.B(n_440),
.C(n_422),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_495),
.B(n_496),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_469),
.B(n_422),
.C(n_419),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_453),
.B(n_427),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_458),
.A2(n_433),
.B(n_424),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_460),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_455),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_454),
.Y(n_507)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_457),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_500),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_514),
.Y(n_520)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_507),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_480),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_510),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_482),
.B(n_465),
.C(n_467),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_451),
.C(n_466),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_512),
.B(n_515),
.Y(n_533)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_480),
.B(n_466),
.CI(n_468),
.CON(n_514),
.SN(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_483),
.B(n_450),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_470),
.C(n_447),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_517),
.B(n_479),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_518),
.A2(n_488),
.B1(n_462),
.B2(n_463),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_491),
.B(n_449),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_479),
.C(n_494),
.Y(n_523)
);

CKINVDCx14_ASAP7_75t_R g521 ( 
.A(n_504),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_521),
.B(n_526),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_506),
.B(n_477),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_522),
.B(n_529),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_535),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_514),
.Y(n_524)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_524),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_502),
.A2(n_487),
.B1(n_476),
.B2(n_498),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_525),
.A2(n_502),
.B1(n_508),
.B2(n_487),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_483),
.C(n_495),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_496),
.C(n_485),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_527),
.A2(n_531),
.B(n_536),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_484),
.Y(n_528)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_528),
.Y(n_540)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_515),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_513),
.B(n_489),
.C(n_497),
.Y(n_531)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_532),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_512),
.A2(n_490),
.B(n_473),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_524),
.B(n_501),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_538),
.B(n_532),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_533),
.C(n_527),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_547),
.C(n_550),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_490),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_513),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_546),
.B(n_534),
.C(n_520),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_517),
.C(n_501),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_525),
.B(n_505),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_528),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_523),
.B(n_516),
.C(n_519),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_551),
.B(n_553),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_552),
.B(n_555),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_540),
.A2(n_503),
.B1(n_457),
.B2(n_478),
.Y(n_553)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_556),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_545),
.B(n_493),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_557),
.B(n_560),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_541),
.B(n_520),
.C(n_445),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_558),
.A2(n_559),
.B(n_561),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_544),
.C(n_547),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_539),
.A2(n_417),
.B1(n_430),
.B2(n_424),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_417),
.Y(n_561)
);

INVx11_ASAP7_75t_L g564 ( 
.A(n_554),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_564),
.A2(n_565),
.B(n_561),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_554),
.A2(n_550),
.B(n_543),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_567),
.A2(n_538),
.B(n_542),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_569),
.A2(n_570),
.B(n_571),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_566),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_562),
.A2(n_552),
.B(n_555),
.Y(n_571)
);

AO21x2_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_563),
.B(n_568),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_563),
.Y(n_575)
);

AOI322xp5_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_568),
.A3(n_573),
.B1(n_548),
.B2(n_425),
.C1(n_276),
.C2(n_15),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_576),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_15),
.C(n_12),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_578),
.A2(n_13),
.B(n_15),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_13),
.B(n_539),
.Y(n_580)
);


endmodule