module fake_aes_6319_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
INVx1_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
AND2x4_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .Y(n_4) );
NAND3xp33_ASAP7_75t_L g5 ( .A(n_4), .B(n_0), .C(n_1), .Y(n_5) );
AND2x4_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
AOI22xp33_ASAP7_75t_L g7 ( .A1(n_6), .A2(n_4), .B1(n_3), .B2(n_0), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_5), .B(n_4), .Y(n_8) );
AND2x4_ASAP7_75t_L g9 ( .A(n_8), .B(n_3), .Y(n_9) );
OAI211xp5_ASAP7_75t_SL g10 ( .A1(n_9), .A2(n_7), .B(n_2), .C(n_1), .Y(n_10) );
AOI211xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_2), .B(n_8), .C(n_5), .Y(n_11) );
CKINVDCx16_ASAP7_75t_R g12 ( .A(n_11), .Y(n_12) );
OA21x2_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_9), .B(n_10), .Y(n_13) );
endmodule