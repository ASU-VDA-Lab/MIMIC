module fake_netlist_6_2079_n_1729 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1729);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1729;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_81),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_37),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_82),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_37),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_47),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_38),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_28),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_13),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_2),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_26),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_55),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_57),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_74),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_7),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_46),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_64),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_30),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_34),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_60),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_4),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_54),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_89),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_34),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_69),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_51),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_83),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_73),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_18),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_24),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_67),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_20),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_21),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_14),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_19),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_101),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_42),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_75),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_70),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_24),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_92),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_154),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_21),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_97),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_54),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_17),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_113),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_125),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_153),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_138),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_53),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_3),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_3),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_77),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_36),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_27),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_126),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_87),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_146),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_155),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_124),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_47),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_30),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_0),
.Y(n_245)
);

BUFx8_ASAP7_75t_SL g246 ( 
.A(n_43),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_42),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_0),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_102),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_23),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_109),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_18),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_111),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_104),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_147),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_31),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_123),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_72),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_127),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_46),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_20),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_114),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_103),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_62),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_140),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_100),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_41),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_6),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_115),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_68),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_5),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_19),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_39),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_40),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_106),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_41),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_36),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_91),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_16),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_53),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_76),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_51),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_4),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_116),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_118),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_27),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_14),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_107),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_7),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_59),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_12),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_25),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_144),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_35),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_148),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_49),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_135),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_58),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_8),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_28),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_12),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_214),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_246),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_193),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_260),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_195),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_221),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_240),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_286),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_189),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_196),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_198),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_201),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_210),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_213),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_174),
.B(n_1),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_217),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_219),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_223),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_220),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_202),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_227),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_202),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_228),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_239),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_241),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_248),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_200),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_250),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_252),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_170),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_205),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_247),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_274),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_254),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_255),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_256),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_233),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_157),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_161),
.B(n_1),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_194),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_206),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_221),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_208),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_157),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_167),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_159),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_242),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_209),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_215),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_230),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_164),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_231),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_173),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_309),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_181),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_185),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_282),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_190),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_235),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_192),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_177),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_199),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_314),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_317),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_161),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_242),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_361),
.B(n_187),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_328),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_337),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_315),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_329),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_320),
.B(n_187),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_320),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_331),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_312),
.A2(n_266),
.B1(n_285),
.B2(n_169),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_368),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_323),
.A2(n_218),
.B(n_211),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_323),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_332),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_333),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_336),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_340),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_324),
.B(n_360),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_316),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_339),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_374),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_342),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_339),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_376),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_341),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_324),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_364),
.B(n_177),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_344),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_345),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_341),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_343),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_346),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_378),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_343),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_366),
.Y(n_451)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_334),
.B(n_302),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_330),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_379),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_352),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_353),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g458 ( 
.A1(n_453),
.A2(n_302),
.B1(n_156),
.B2(n_204),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_453),
.A2(n_347),
.B1(n_357),
.B2(n_356),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_426),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_396),
.B(n_371),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_426),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_348),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_L g464 ( 
.A(n_396),
.B(n_223),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_372),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_414),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_354),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_414),
.B(n_385),
.Y(n_471)
);

OAI22xp33_ASAP7_75t_L g472 ( 
.A1(n_392),
.A2(n_186),
.B1(n_238),
.B2(n_327),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_439),
.B(n_156),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_424),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_373),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_424),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_439),
.B(n_204),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_431),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_440),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_390),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_393),
.B(n_375),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

BUFx6f_ASAP7_75t_SL g488 ( 
.A(n_431),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_452),
.A2(n_349),
.B1(n_338),
.B2(n_335),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_400),
.Y(n_491)
);

BUFx6f_ASAP7_75t_SL g492 ( 
.A(n_435),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_393),
.B(n_382),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_393),
.B(n_380),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_395),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_395),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_452),
.B(n_360),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_395),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_416),
.B(n_313),
.Y(n_500)
);

INVx4_ASAP7_75t_SL g501 ( 
.A(n_400),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_407),
.B(n_362),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_417),
.A2(n_212),
.B1(n_234),
.B2(n_289),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_407),
.B(n_362),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_452),
.B(n_222),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_436),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_427),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_390),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_438),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_392),
.B(n_212),
.Y(n_512)
);

NOR2x1p5_ASAP7_75t_L g513 ( 
.A(n_388),
.B(n_168),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_387),
.B(n_160),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_387),
.B(n_394),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_433),
.B(n_359),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_433),
.B(n_367),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_438),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_440),
.B(n_234),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_451),
.B(n_384),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_429),
.B(n_298),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_429),
.B(n_379),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_446),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_389),
.B(n_289),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_446),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_448),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_452),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_417),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_394),
.B(n_175),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_455),
.B(n_381),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_397),
.A2(n_325),
.B1(n_326),
.B2(n_191),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_451),
.B(n_381),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_417),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_391),
.B(n_402),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_416),
.B(n_383),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_399),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_405),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_405),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_410),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_399),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_427),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_401),
.B(n_269),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_412),
.B(n_383),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_403),
.B(n_300),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_421),
.B(n_385),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_391),
.Y(n_553)
);

BUFx4f_ASAP7_75t_L g554 ( 
.A(n_452),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_410),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_422),
.B(n_425),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_403),
.B(n_158),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_432),
.B(n_178),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_406),
.B(n_353),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_413),
.B(n_232),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_404),
.B(n_162),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_404),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_410),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_400),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_400),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_417),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_408),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_398),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_441),
.B(n_163),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_415),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_400),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_415),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_409),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_442),
.A2(n_236),
.B1(n_243),
.B2(n_244),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_418),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_411),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_447),
.B(n_178),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_L g579 ( 
.A(n_406),
.B(n_223),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_SL g580 ( 
.A(n_413),
.B(n_168),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_428),
.B(n_165),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_437),
.B(n_166),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_437),
.B(n_176),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_454),
.B(n_182),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_419),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_418),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_418),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_419),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_420),
.B(n_418),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_428),
.B(n_355),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_415),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_420),
.B(n_197),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_437),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_418),
.B(n_207),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_434),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_437),
.B(n_216),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_418),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_L g599 ( 
.A(n_437),
.B(n_223),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_398),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_437),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_461),
.B(n_457),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_461),
.B(n_596),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_486),
.B(n_182),
.Y(n_604)
);

INVx8_ASAP7_75t_L g605 ( 
.A(n_498),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_485),
.A2(n_398),
.B(n_434),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_466),
.B(n_457),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_460),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_466),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_554),
.B(n_223),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_493),
.B(n_457),
.Y(n_611)
);

AND2x6_ASAP7_75t_SL g612 ( 
.A(n_560),
.B(n_251),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_462),
.A2(n_273),
.B1(n_225),
.B2(n_191),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_473),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_468),
.B(n_470),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_473),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_473),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_550),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_554),
.B(n_223),
.Y(n_619)
);

INVx8_ASAP7_75t_L g620 ( 
.A(n_498),
.Y(n_620)
);

NAND3xp33_ASAP7_75t_L g621 ( 
.A(n_538),
.B(n_253),
.C(n_249),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_510),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_475),
.B(n_437),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_538),
.B(n_550),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_510),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_524),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_476),
.B(n_443),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_503),
.B(n_223),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_478),
.B(n_443),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_503),
.B(n_223),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_533),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_560),
.A2(n_270),
.B1(n_277),
.B2(n_281),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_535),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_482),
.B(n_443),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_483),
.B(n_496),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_494),
.B(n_552),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_510),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_523),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

AND2x6_ASAP7_75t_SL g641 ( 
.A(n_560),
.B(n_284),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_533),
.B(n_297),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_508),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_502),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_552),
.A2(n_184),
.B1(n_183),
.B2(n_225),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_511),
.B(n_518),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_532),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_523),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_471),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_520),
.B(n_443),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_558),
.B(n_183),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_539),
.B(n_297),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_525),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_504),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_559),
.A2(n_287),
.B1(n_288),
.B2(n_291),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_459),
.A2(n_273),
.B1(n_267),
.B2(n_259),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_553),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_558),
.B(n_184),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_578),
.B(n_188),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_539),
.A2(n_301),
.B1(n_297),
.B2(n_237),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_527),
.B(n_443),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_541),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_530),
.B(n_443),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_549),
.B(n_297),
.Y(n_664)
);

BUFx6f_ASAP7_75t_SL g665 ( 
.A(n_535),
.Y(n_665)
);

NOR2x2_ASAP7_75t_L g666 ( 
.A(n_505),
.B(n_203),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_484),
.B(n_226),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_531),
.B(n_443),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_578),
.B(n_188),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_549),
.B(n_297),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_523),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_469),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_536),
.B(n_449),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_529),
.B(n_258),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_591),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_566),
.B(n_297),
.Y(n_676)
);

INVx5_ASAP7_75t_L g677 ( 
.A(n_557),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_542),
.B(n_449),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_529),
.B(n_570),
.Y(n_679)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_458),
.B(n_229),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_469),
.Y(n_681)
);

INVx6_ASAP7_75t_L g682 ( 
.A(n_471),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_546),
.B(n_449),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_471),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_535),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_566),
.B(n_532),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_521),
.A2(n_167),
.B1(n_275),
.B2(n_304),
.Y(n_687)
);

AND2x6_ASAP7_75t_SL g688 ( 
.A(n_521),
.B(n_355),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_562),
.B(n_567),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_465),
.A2(n_305),
.B1(n_280),
.B2(n_283),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_568),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_570),
.B(n_258),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_487),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_477),
.B(n_297),
.Y(n_694)
);

AND2x4_ASAP7_75t_SL g695 ( 
.A(n_498),
.B(n_167),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_505),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_557),
.B(n_458),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_487),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_465),
.B(n_259),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_505),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_540),
.B(n_203),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_574),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_512),
.A2(n_279),
.B(n_264),
.C(n_265),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_519),
.B(n_267),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_577),
.B(n_449),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_581),
.B(n_297),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_512),
.B(n_245),
.C(n_280),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_519),
.A2(n_283),
.B1(n_290),
.B2(n_305),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_585),
.B(n_449),
.Y(n_709)
);

OAI221xp5_ASAP7_75t_L g710 ( 
.A1(n_514),
.A2(n_268),
.B1(n_272),
.B2(n_294),
.C(n_171),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_489),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_589),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_464),
.A2(n_444),
.B(n_290),
.C(n_306),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_489),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_575),
.B(n_306),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_463),
.A2(n_276),
.B1(n_172),
.B2(n_179),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_495),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_581),
.B(n_450),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_534),
.B(n_171),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_467),
.B(n_450),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_590),
.B(n_450),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_515),
.B(n_450),
.Y(n_722)
);

OAI22x1_ASAP7_75t_L g723 ( 
.A1(n_584),
.A2(n_509),
.B1(n_547),
.B2(n_537),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_548),
.B(n_450),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_495),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_513),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_497),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_SL g728 ( 
.A1(n_490),
.A2(n_172),
.B1(n_179),
.B2(n_180),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_551),
.B(n_472),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_497),
.Y(n_730)
);

AND2x6_ASAP7_75t_SL g731 ( 
.A(n_556),
.B(n_203),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_464),
.A2(n_292),
.B1(n_224),
.B2(n_261),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_601),
.B(n_444),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_499),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_601),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_565),
.B(n_576),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_474),
.A2(n_398),
.B(n_444),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_565),
.B(n_456),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_565),
.B(n_456),
.Y(n_739)
);

NAND2x1_ASAP7_75t_L g740 ( 
.A(n_576),
.B(n_398),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_488),
.B(n_180),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_499),
.Y(n_742)
);

NOR2x1_ASAP7_75t_R g743 ( 
.A(n_516),
.B(n_278),
.Y(n_743)
);

AO221x1_ASAP7_75t_L g744 ( 
.A1(n_580),
.A2(n_304),
.B1(n_275),
.B2(n_262),
.C(n_263),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_526),
.Y(n_745)
);

INVx8_ASAP7_75t_L g746 ( 
.A(n_488),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_517),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_576),
.B(n_456),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_561),
.B(n_456),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_593),
.B(n_456),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_580),
.A2(n_292),
.B(n_261),
.C(n_307),
.Y(n_751)
);

BUFx12f_ASAP7_75t_L g752 ( 
.A(n_557),
.Y(n_752)
);

AND2x4_ASAP7_75t_SL g753 ( 
.A(n_556),
.B(n_275),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_491),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_594),
.B(n_398),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_598),
.B(n_456),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_543),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_543),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_544),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_474),
.B(n_307),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_481),
.B(n_224),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_481),
.B(n_262),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_492),
.A2(n_557),
.B1(n_579),
.B2(n_500),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_595),
.B(n_491),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_544),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_545),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_720),
.A2(n_600),
.B(n_569),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_634),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_688),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_736),
.A2(n_582),
.B(n_583),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_657),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_624),
.B(n_545),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_611),
.A2(n_600),
.B(n_569),
.Y(n_773)
);

AND2x6_ASAP7_75t_L g774 ( 
.A(n_631),
.B(n_491),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_685),
.B(n_501),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_724),
.A2(n_600),
.B(n_569),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_642),
.A2(n_579),
.B(n_597),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_642),
.A2(n_582),
.B(n_597),
.Y(n_778)
);

AND2x6_ASAP7_75t_L g779 ( 
.A(n_631),
.B(n_763),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_662),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_679),
.A2(n_522),
.B(n_583),
.C(n_599),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_624),
.A2(n_603),
.B(n_729),
.C(n_679),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_729),
.A2(n_522),
.B(n_599),
.C(n_592),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_637),
.B(n_557),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_626),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_699),
.B(n_555),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_699),
.B(n_555),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_602),
.A2(n_480),
.B(n_588),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_618),
.B(n_563),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_764),
.A2(n_480),
.B(n_588),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_626),
.Y(n_791)
);

AO22x1_ASAP7_75t_L g792 ( 
.A1(n_715),
.A2(n_296),
.B1(n_271),
.B2(n_276),
.Y(n_792)
);

AOI22x1_ASAP7_75t_L g793 ( 
.A1(n_614),
.A2(n_592),
.B1(n_563),
.B2(n_571),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_651),
.B(n_571),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_764),
.A2(n_722),
.B(n_697),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_631),
.A2(n_492),
.B1(n_573),
.B2(n_586),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_686),
.A2(n_588),
.B(n_507),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_651),
.B(n_573),
.Y(n_798)
);

AOI21x1_ASAP7_75t_L g799 ( 
.A1(n_652),
.A2(n_501),
.B(n_586),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_686),
.A2(n_491),
.B(n_586),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_658),
.B(n_586),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_608),
.B(n_501),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_631),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_607),
.A2(n_564),
.B(n_528),
.Y(n_804)
);

O2A1O1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_652),
.A2(n_263),
.B(n_271),
.C(n_278),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_664),
.A2(n_293),
.B(n_295),
.C(n_296),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_733),
.A2(n_507),
.B(n_564),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_718),
.A2(n_507),
.B(n_564),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_634),
.A2(n_507),
.B1(n_528),
.B2(n_564),
.Y(n_809)
);

NAND2x1p5_ASAP7_75t_L g810 ( 
.A(n_649),
.B(n_647),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_658),
.B(n_528),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_659),
.B(n_528),
.Y(n_812)
);

AO32x1_ASAP7_75t_L g813 ( 
.A1(n_633),
.A2(n_643),
.A3(n_702),
.B1(n_691),
.B2(n_712),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_692),
.A2(n_303),
.B(n_295),
.C(n_293),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_718),
.A2(n_587),
.B(n_572),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_659),
.B(n_303),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_747),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_649),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_669),
.B(n_587),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_692),
.A2(n_587),
.B(n_572),
.C(n_304),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_669),
.B(n_572),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_604),
.B(n_56),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_660),
.A2(n_152),
.B1(n_136),
.B2(n_133),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_670),
.A2(n_129),
.B(n_128),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_604),
.B(n_2),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_676),
.A2(n_122),
.B(n_119),
.Y(n_826)
);

INVxp33_ASAP7_75t_SL g827 ( 
.A(n_743),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_735),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_684),
.B(n_86),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_721),
.A2(n_110),
.B(n_99),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_721),
.A2(n_677),
.B(n_694),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_677),
.A2(n_98),
.B(n_96),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_677),
.A2(n_94),
.B(n_93),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_674),
.B(n_90),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_677),
.A2(n_85),
.B(n_79),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_674),
.B(n_78),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_615),
.A2(n_5),
.B(n_8),
.C(n_9),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_694),
.A2(n_71),
.B(n_66),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_640),
.Y(n_839)
);

OAI21xp33_ASAP7_75t_L g840 ( 
.A1(n_719),
.A2(n_645),
.B(n_715),
.Y(n_840)
);

BUFx2_ASAP7_75t_SL g841 ( 
.A(n_665),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_609),
.A2(n_61),
.B(n_10),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_660),
.A2(n_52),
.B1(n_10),
.B2(n_11),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_609),
.A2(n_9),
.B(n_11),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_701),
.B(n_15),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_636),
.A2(n_15),
.B(n_22),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_644),
.B(n_52),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_628),
.A2(n_22),
.B(n_23),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_606),
.A2(n_25),
.B(n_26),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_704),
.A2(n_29),
.B(n_31),
.Y(n_850)
);

BUFx8_ASAP7_75t_L g851 ( 
.A(n_665),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_628),
.A2(n_29),
.B(n_32),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_682),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_646),
.A2(n_32),
.B(n_33),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_630),
.A2(n_39),
.B(n_40),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_654),
.B(n_44),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_704),
.A2(n_44),
.B(n_45),
.C(n_48),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_653),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_719),
.B(n_48),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_656),
.B(n_50),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_675),
.B(n_50),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_753),
.B(n_689),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_754),
.A2(n_610),
.B(n_619),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_682),
.A2(n_647),
.B1(n_680),
.B2(n_605),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_754),
.A2(n_610),
.B(n_619),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_754),
.A2(n_755),
.B(n_709),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_754),
.A2(n_755),
.B(n_705),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_703),
.A2(n_761),
.B(n_760),
.C(n_762),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_725),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_753),
.B(n_741),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_623),
.A2(n_683),
.B(n_678),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_621),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_680),
.B(n_616),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_617),
.B(n_622),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_625),
.B(n_638),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_639),
.B(n_648),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_734),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_627),
.A2(n_650),
.B(n_668),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_629),
.A2(n_673),
.B(n_635),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_630),
.A2(n_713),
.B(n_766),
.Y(n_880)
);

CKINVDCx10_ASAP7_75t_R g881 ( 
.A(n_667),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_671),
.B(n_742),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_745),
.B(n_714),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_703),
.A2(n_710),
.B(n_751),
.C(n_655),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_672),
.B(n_717),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_681),
.B(n_698),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_661),
.A2(n_663),
.B(n_749),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_693),
.B(n_727),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_711),
.A2(n_765),
.B(n_759),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_730),
.B(n_757),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_750),
.A2(n_739),
.B(n_738),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_758),
.A2(n_706),
.B(n_707),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_682),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_605),
.B(n_620),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_751),
.A2(n_655),
.B(n_632),
.C(n_716),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_748),
.A2(n_706),
.B(n_756),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_696),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_740),
.A2(n_737),
.B(n_700),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_667),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_735),
.A2(n_605),
.B(n_620),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_726),
.A2(n_752),
.B1(n_667),
.B2(n_620),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_735),
.A2(n_695),
.B(n_613),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_735),
.A2(n_690),
.B1(n_687),
.B2(n_723),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_708),
.A2(n_632),
.B(n_732),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_612),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_732),
.A2(n_744),
.B(n_746),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_728),
.A2(n_746),
.B1(n_666),
.B2(n_641),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_746),
.A2(n_720),
.B(n_611),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_731),
.A2(n_624),
.B(n_603),
.C(n_729),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_624),
.B(n_603),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_624),
.B(n_521),
.C(n_459),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_603),
.B(n_679),
.Y(n_913)
);

AND2x4_ASAP7_75t_SL g914 ( 
.A(n_696),
.B(n_427),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_624),
.B(n_603),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_624),
.A2(n_603),
.B(n_729),
.C(n_396),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_642),
.A2(n_664),
.B(n_652),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_624),
.B(n_603),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_637),
.B(n_624),
.Y(n_921)
);

OAI22xp33_ASAP7_75t_L g922 ( 
.A1(n_603),
.A2(n_624),
.B1(n_618),
.B2(n_679),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_637),
.B(n_624),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_657),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_927)
);

INVx11_ASAP7_75t_L g928 ( 
.A(n_752),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_603),
.B(n_679),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_657),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_624),
.B(n_603),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_679),
.A2(n_624),
.B1(n_729),
.B2(n_637),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_649),
.Y(n_936)
);

AND2x2_ASAP7_75t_SL g937 ( 
.A(n_753),
.B(n_416),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_618),
.B(n_624),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_624),
.A2(n_679),
.B(n_694),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_746),
.B(n_605),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_637),
.B(n_624),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_618),
.B(n_624),
.Y(n_944)
);

INVx11_ASAP7_75t_L g945 ( 
.A(n_752),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_634),
.Y(n_946)
);

OAI22x1_ASAP7_75t_L g947 ( 
.A1(n_624),
.A2(n_618),
.B1(n_679),
.B2(n_584),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_657),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_720),
.A2(n_611),
.B(n_724),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_624),
.B(n_603),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_910),
.B(n_915),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_921),
.B(n_924),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_896),
.A2(n_891),
.B(n_799),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_795),
.A2(n_918),
.B(n_873),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_873),
.A2(n_782),
.B(n_880),
.Y(n_955)
);

NOR2x1_ASAP7_75t_SL g956 ( 
.A(n_803),
.B(n_834),
.Y(n_956)
);

AO31x2_ASAP7_75t_L g957 ( 
.A1(n_940),
.A2(n_783),
.A3(n_781),
.B(n_820),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_821),
.A2(n_811),
.B(n_801),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_840),
.A2(n_904),
.B1(n_912),
.B2(n_843),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_916),
.A2(n_868),
.B(n_777),
.Y(n_960)
);

CKINVDCx16_ASAP7_75t_R g961 ( 
.A(n_941),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_934),
.A2(n_950),
.B1(n_910),
.B2(n_933),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_915),
.B(n_920),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_911),
.A2(n_919),
.B(n_917),
.Y(n_964)
);

AO31x2_ASAP7_75t_L g965 ( 
.A1(n_923),
.A2(n_927),
.A3(n_949),
.B(n_926),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_920),
.B(n_933),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_913),
.A2(n_929),
.B(n_865),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_950),
.A2(n_938),
.B1(n_944),
.B2(n_922),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_943),
.B(n_789),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_772),
.B(n_859),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_772),
.B(n_839),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_851),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_870),
.B(n_845),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_770),
.A2(n_887),
.B(n_878),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_851),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_860),
.A2(n_895),
.B(n_855),
.C(n_852),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_797),
.A2(n_800),
.B(n_793),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_863),
.A2(n_778),
.B(n_786),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_930),
.A2(n_935),
.B(n_939),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_803),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_858),
.Y(n_981)
);

NOR2xp67_ASAP7_75t_L g982 ( 
.A(n_948),
.B(n_771),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_871),
.A2(n_879),
.B(n_831),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_883),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_825),
.B(n_794),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_787),
.A2(n_798),
.B(n_942),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_883),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_848),
.A2(n_909),
.B(n_884),
.C(n_850),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_803),
.B(n_853),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_L g990 ( 
.A1(n_822),
.A2(n_812),
.B(n_932),
.C(n_836),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_931),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_808),
.A2(n_867),
.B(n_866),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_941),
.Y(n_993)
);

OAI21x1_ASAP7_75t_L g994 ( 
.A1(n_790),
.A2(n_804),
.B(n_807),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_908),
.A2(n_819),
.B(n_784),
.Y(n_995)
);

AOI21xp33_ASAP7_75t_L g996 ( 
.A1(n_816),
.A2(n_947),
.B(n_872),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_869),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_818),
.A2(n_936),
.B(n_788),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_928),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_882),
.A2(n_876),
.B(n_875),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_882),
.A2(n_876),
.B(n_875),
.Y(n_1001)
);

AO31x2_ASAP7_75t_L g1002 ( 
.A1(n_857),
.A2(n_814),
.A3(n_846),
.B(n_854),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_767),
.A2(n_776),
.B(n_773),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_785),
.B(n_791),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_824),
.A2(n_837),
.B(n_805),
.C(n_806),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_818),
.A2(n_936),
.B(n_828),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_817),
.B(n_925),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_864),
.B(n_829),
.Y(n_1008)
);

NOR2xp67_ASAP7_75t_SL g1009 ( 
.A(n_841),
.B(n_853),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_829),
.B(n_768),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_889),
.A2(n_815),
.B(n_874),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_823),
.A2(n_856),
.B(n_844),
.C(n_906),
.Y(n_1012)
);

AOI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_862),
.A2(n_780),
.B(n_897),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_903),
.A2(n_902),
.B(n_861),
.C(n_842),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_898),
.A2(n_892),
.B(n_809),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_885),
.A2(n_886),
.B(n_888),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_885),
.Y(n_1017)
);

AOI221x1_ASAP7_75t_L g1018 ( 
.A1(n_796),
.A2(n_838),
.B1(n_826),
.B2(n_830),
.C(n_946),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_901),
.B(n_899),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_849),
.A2(n_810),
.B(n_900),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_886),
.A2(n_888),
.B(n_890),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_847),
.A2(n_890),
.B(n_893),
.C(n_877),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_810),
.A2(n_775),
.B(n_802),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_779),
.B(n_802),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_832),
.A2(n_835),
.B(n_833),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_779),
.A2(n_775),
.B(n_774),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_894),
.A2(n_774),
.B(n_813),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_774),
.A2(n_813),
.B(n_779),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_774),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_779),
.B(n_792),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_941),
.A2(n_937),
.B(n_914),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_945),
.Y(n_1032)
);

AOI211x1_ASAP7_75t_L g1033 ( 
.A1(n_907),
.A2(n_769),
.B(n_881),
.C(n_905),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_905),
.A2(n_827),
.B(n_896),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_821),
.A2(n_811),
.B(n_801),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_921),
.B(n_637),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_771),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_793),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_771),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_911),
.A2(n_919),
.B(n_917),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_910),
.B(n_915),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_910),
.B(n_915),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_793),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_795),
.A2(n_891),
.B(n_896),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_910),
.B(n_915),
.Y(n_1045)
);

O2A1O1Ixp5_ASAP7_75t_L g1046 ( 
.A1(n_825),
.A2(n_940),
.B(n_859),
.C(n_694),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_795),
.A2(n_891),
.B(n_896),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_938),
.B(n_944),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_910),
.B(n_915),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_839),
.Y(n_1050)
);

NAND2x1_ASAP7_75t_L g1051 ( 
.A(n_774),
.B(n_631),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_803),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_771),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_938),
.B(n_944),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_L g1055 ( 
.A(n_779),
.B(n_631),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_896),
.A2(n_891),
.B(n_799),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_934),
.A2(n_915),
.B1(n_920),
.B2(n_910),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_803),
.B(n_631),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_774),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_839),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_912),
.A2(n_840),
.B1(n_624),
.B2(n_938),
.Y(n_1061)
);

INVx8_ASAP7_75t_L g1062 ( 
.A(n_941),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_910),
.B(n_915),
.Y(n_1063)
);

OA21x2_ASAP7_75t_L g1064 ( 
.A1(n_880),
.A2(n_917),
.B(n_911),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_911),
.A2(n_919),
.B(n_917),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_910),
.B(n_915),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_825),
.A2(n_940),
.B(n_859),
.C(n_694),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_921),
.B(n_637),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_910),
.B(n_915),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_795),
.A2(n_918),
.B(n_873),
.Y(n_1070)
);

AND2x2_ASAP7_75t_SL g1071 ( 
.A(n_912),
.B(n_680),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_910),
.B(n_915),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_803),
.B(n_631),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_911),
.A2(n_919),
.B(n_917),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_896),
.A2(n_891),
.B(n_799),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_911),
.A2(n_919),
.B(n_917),
.Y(n_1076)
);

OA22x2_ASAP7_75t_L g1077 ( 
.A1(n_840),
.A2(n_560),
.B1(n_934),
.B2(n_618),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_793),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_940),
.A2(n_783),
.A3(n_781),
.B(n_795),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_910),
.B(n_915),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_931),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_803),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_911),
.A2(n_919),
.B(n_917),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_896),
.A2(n_891),
.B(n_799),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_911),
.A2(n_919),
.B(n_917),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_934),
.B(n_782),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_839),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_900),
.B(n_853),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_795),
.A2(n_918),
.B(n_873),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_896),
.A2(n_891),
.B(n_799),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_803),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_896),
.A2(n_891),
.B(n_799),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_785),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_795),
.A2(n_918),
.B(n_873),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_851),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_896),
.A2(n_891),
.B(n_799),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_803),
.B(n_631),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1020),
.A2(n_1056),
.B(n_953),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_951),
.B(n_963),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_966),
.B(n_1041),
.Y(n_1100)
);

NOR2x1_ASAP7_75t_SL g1101 ( 
.A(n_1059),
.B(n_1008),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1042),
.B(n_1045),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1071),
.A2(n_1077),
.B1(n_959),
.B2(n_1048),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_972),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_960),
.A2(n_955),
.B(n_1015),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1065),
.A2(n_1076),
.B(n_1074),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_975),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1000),
.A2(n_1001),
.B(n_995),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1049),
.B(n_1063),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_993),
.B(n_1032),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_981),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1066),
.B(n_1069),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1072),
.B(n_1080),
.Y(n_1114)
);

BUFx4_ASAP7_75t_SL g1115 ( 
.A(n_972),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_952),
.B(n_1036),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_962),
.B(n_1057),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_1068),
.B(n_991),
.Y(n_1118)
);

INVx5_ASAP7_75t_L g1119 ( 
.A(n_1059),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1083),
.A2(n_1085),
.B(n_986),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1050),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1020),
.A2(n_1084),
.B(n_1096),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_1062),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_999),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_SL g1125 ( 
.A(n_1059),
.B(n_999),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_978),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_968),
.B(n_1048),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_975),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_1007),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1060),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1055),
.A2(n_1064),
.B(n_990),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_1093),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1071),
.A2(n_1077),
.B1(n_959),
.B2(n_1054),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_SL g1134 ( 
.A(n_1059),
.B(n_1008),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_1062),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1004),
.Y(n_1136)
);

OR2x6_ASAP7_75t_L g1137 ( 
.A(n_1062),
.B(n_1031),
.Y(n_1137)
);

CKINVDCx11_ASAP7_75t_R g1138 ( 
.A(n_1081),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1087),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1054),
.B(n_1061),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1058),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_973),
.A2(n_1019),
.B1(n_969),
.B2(n_976),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1037),
.Y(n_1143)
);

AND2x6_ASAP7_75t_L g1144 ( 
.A(n_1029),
.B(n_1088),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_976),
.A2(n_988),
.B1(n_971),
.B2(n_987),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1053),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1039),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_997),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_990),
.A2(n_1064),
.B(n_998),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_954),
.A2(n_1070),
.B(n_1094),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1026),
.B(n_1023),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1093),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_988),
.A2(n_984),
.B1(n_970),
.B2(n_1086),
.Y(n_1153)
);

OAI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1030),
.A2(n_985),
.B1(n_1010),
.B2(n_961),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1017),
.B(n_1086),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1016),
.B(n_1021),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_980),
.Y(n_1157)
);

BUFx2_ASAP7_75t_R g1158 ( 
.A(n_1095),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1089),
.A2(n_983),
.B(n_1044),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_982),
.B(n_996),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_993),
.B(n_1034),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1073),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_967),
.B(n_1014),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1073),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1033),
.A2(n_1095),
.B1(n_1024),
.B2(n_989),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1091),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1013),
.B(n_1002),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1097),
.Y(n_1168)
);

BUFx2_ASAP7_75t_SL g1169 ( 
.A(n_1052),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1082),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1002),
.B(n_1091),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1082),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1014),
.B(n_1012),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1082),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_989),
.B(n_1051),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1088),
.B(n_980),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_L g1177 ( 
.A1(n_1046),
.A2(n_1067),
.B(n_1027),
.C(n_1005),
.Y(n_1177)
);

INVx5_ASAP7_75t_L g1178 ( 
.A(n_1088),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1044),
.A2(n_1047),
.B(n_983),
.Y(n_1179)
);

BUFx4f_ASAP7_75t_L g1180 ( 
.A(n_1009),
.Y(n_1180)
);

AOI21xp33_ASAP7_75t_L g1181 ( 
.A1(n_1046),
.A2(n_1067),
.B(n_1022),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1047),
.A2(n_974),
.B(n_1003),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1038),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1002),
.B(n_956),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1079),
.B(n_1002),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1079),
.B(n_957),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1079),
.B(n_957),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1079),
.B(n_957),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1006),
.B(n_1018),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_957),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_958),
.B(n_1035),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1028),
.A2(n_992),
.B1(n_1011),
.B2(n_1078),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1075),
.B(n_1092),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_965),
.B(n_1038),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1090),
.B(n_1025),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_L g1196 ( 
.A(n_1043),
.B(n_965),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_994),
.Y(n_1197)
);

AO21x2_ASAP7_75t_L g1198 ( 
.A1(n_974),
.A2(n_977),
.B(n_965),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_965),
.B(n_1036),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_951),
.B(n_963),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_981),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_981),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_952),
.B(n_509),
.Y(n_1203)
);

AOI22x1_ASAP7_75t_L g1204 ( 
.A1(n_960),
.A2(n_947),
.B1(n_904),
.B2(n_908),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_981),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_981),
.Y(n_1207)
);

AND3x2_ASAP7_75t_L g1208 ( 
.A(n_1048),
.B(n_860),
.C(n_912),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1053),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_SL g1210 ( 
.A(n_976),
.B(n_840),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_975),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_981),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1036),
.B(n_1068),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1007),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_951),
.B(n_963),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_999),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_993),
.B(n_1032),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1004),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_993),
.B(n_1032),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_1055),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1036),
.B(n_1068),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1061),
.B(n_934),
.Y(n_1225)
);

BUFx5_ASAP7_75t_L g1226 ( 
.A(n_1088),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1058),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1053),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1062),
.B(n_941),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_964),
.A2(n_1040),
.B(n_979),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1036),
.B(n_1068),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1103),
.B(n_1133),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1121),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1130),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1139),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1201),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1123),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1202),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1207),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1099),
.B(n_1100),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1099),
.A2(n_1113),
.B1(n_1100),
.B2(n_1110),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1132),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1136),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1210),
.A2(n_1225),
.B1(n_1140),
.B2(n_1127),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1136),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1177),
.A2(n_1181),
.B(n_1149),
.Y(n_1248)
);

INVxp67_ASAP7_75t_L g1249 ( 
.A(n_1118),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1210),
.A2(n_1140),
.B1(n_1127),
.B2(n_1142),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1112),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1183),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1160),
.A2(n_1110),
.B1(n_1218),
.B2(n_1102),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1102),
.A2(n_1114),
.B1(n_1218),
.B2(n_1113),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1183),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1174),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1183),
.Y(n_1257)
);

OA21x2_ASAP7_75t_L g1258 ( 
.A1(n_1181),
.A2(n_1131),
.B(n_1179),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1146),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1183),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1208),
.A2(n_1117),
.B1(n_1173),
.B2(n_1204),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1165),
.A2(n_1233),
.B1(n_1213),
.B2(n_1224),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1137),
.B(n_1176),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1114),
.A2(n_1200),
.B1(n_1223),
.B2(n_1178),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1117),
.A2(n_1173),
.B(n_1153),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1209),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1098),
.A2(n_1122),
.B(n_1182),
.Y(n_1267)
);

INVx1_ASAP7_75t_SL g1268 ( 
.A(n_1138),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1148),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1105),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1131),
.A2(n_1179),
.B(n_1104),
.Y(n_1271)
);

AOI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1196),
.A2(n_1109),
.B(n_1126),
.Y(n_1272)
);

BUFx12f_ASAP7_75t_L g1273 ( 
.A(n_1219),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1206),
.Y(n_1274)
);

BUFx8_ASAP7_75t_SL g1275 ( 
.A(n_1108),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1200),
.A2(n_1116),
.B1(n_1203),
.B2(n_1221),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1229),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1221),
.B(n_1129),
.Y(n_1278)
);

OR2x6_ASAP7_75t_L g1279 ( 
.A(n_1151),
.B(n_1137),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1212),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1178),
.A2(n_1216),
.B1(n_1155),
.B2(n_1154),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1137),
.A2(n_1153),
.B1(n_1145),
.B2(n_1161),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1180),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1126),
.A2(n_1182),
.B(n_1194),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1174),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1157),
.Y(n_1286)
);

AND2x2_ASAP7_75t_SL g1287 ( 
.A(n_1163),
.B(n_1180),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1115),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1119),
.B(n_1125),
.Y(n_1289)
);

CKINVDCx8_ASAP7_75t_R g1290 ( 
.A(n_1169),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1166),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1155),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1152),
.Y(n_1293)
);

INVxp67_ASAP7_75t_SL g1294 ( 
.A(n_1176),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1171),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1145),
.A2(n_1150),
.B1(n_1163),
.B2(n_1199),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1101),
.A2(n_1134),
.B1(n_1151),
.B2(n_1226),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1159),
.A2(n_1232),
.B(n_1214),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1156),
.A2(n_1120),
.B(n_1191),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1162),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1151),
.A2(n_1143),
.B1(n_1231),
.B2(n_1147),
.Y(n_1301)
);

AO21x1_ASAP7_75t_L g1302 ( 
.A1(n_1156),
.A2(n_1194),
.B(n_1189),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1167),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1231),
.A2(n_1220),
.B1(n_1222),
.B2(n_1111),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1124),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1190),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1106),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1170),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1106),
.A2(n_1187),
.B1(n_1186),
.B2(n_1185),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1111),
.A2(n_1220),
.B1(n_1222),
.B2(n_1135),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1119),
.B(n_1135),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1226),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1231),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1185),
.A2(n_1184),
.B1(n_1189),
.B2(n_1188),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1188),
.B(n_1226),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1158),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1172),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1175),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1141),
.Y(n_1319)
);

INVx6_ASAP7_75t_L g1320 ( 
.A(n_1175),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1164),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1164),
.B(n_1168),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1168),
.B(n_1227),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1128),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1192),
.B(n_1198),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1144),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1175),
.B(n_1198),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1211),
.A2(n_1197),
.B1(n_1228),
.B2(n_1230),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1193),
.B(n_1197),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_1158),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1215),
.A2(n_1107),
.B1(n_1205),
.B2(n_1217),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1193),
.B(n_1195),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1120),
.A2(n_1214),
.B(n_1104),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1121),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1174),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1115),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1199),
.B(n_1140),
.Y(n_1337)
);

INVx5_ASAP7_75t_L g1338 ( 
.A(n_1119),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1116),
.B(n_1136),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1146),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1121),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1303),
.B(n_1337),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1295),
.B(n_1337),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1295),
.B(n_1315),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1267),
.A2(n_1272),
.B(n_1284),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1306),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1245),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1313),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1279),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1265),
.A2(n_1302),
.A3(n_1307),
.B(n_1333),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1315),
.B(n_1309),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1309),
.B(n_1296),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1302),
.Y(n_1353)
);

BUFx2_ASAP7_75t_SL g1354 ( 
.A(n_1338),
.Y(n_1354)
);

AND2x4_ASAP7_75t_SL g1355 ( 
.A(n_1279),
.B(n_1263),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1327),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1314),
.B(n_1296),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1320),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1247),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1314),
.B(n_1299),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1265),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1292),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1320),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1242),
.B(n_1243),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1264),
.A2(n_1267),
.B(n_1281),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1244),
.Y(n_1366)
);

AO21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1282),
.A2(n_1262),
.B(n_1261),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1279),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1254),
.B(n_1253),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1246),
.B(n_1250),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1234),
.B(n_1246),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1331),
.A2(n_1325),
.B(n_1261),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1271),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1234),
.B(n_1332),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1325),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1251),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1287),
.A2(n_1263),
.B1(n_1301),
.B2(n_1276),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1320),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1339),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1332),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1238),
.B(n_1287),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1269),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1294),
.B(n_1286),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1318),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1274),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1277),
.Y(n_1386)
);

OR2x6_ASAP7_75t_L g1387 ( 
.A(n_1263),
.B(n_1312),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1329),
.A2(n_1258),
.B(n_1248),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1280),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1252),
.A2(n_1255),
.B(n_1257),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1249),
.B(n_1298),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1313),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1278),
.B(n_1293),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1235),
.B(n_1236),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1291),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1237),
.B(n_1240),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1321),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1241),
.B(n_1341),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1334),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1252),
.A2(n_1255),
.B(n_1260),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1328),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1326),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1318),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1300),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1318),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1318),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1364),
.B(n_1297),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1351),
.B(n_1319),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1357),
.A2(n_1330),
.B1(n_1310),
.B2(n_1290),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1369),
.B(n_1283),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1390),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1344),
.B(n_1356),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1391),
.B(n_1304),
.Y(n_1414)
);

NOR2x1_ASAP7_75t_SL g1415 ( 
.A(n_1354),
.B(n_1338),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1390),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1353),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1373),
.Y(n_1418)
);

INVxp33_ASAP7_75t_L g1419 ( 
.A(n_1379),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1353),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1369),
.B(n_1283),
.Y(n_1421)
);

AOI211xp5_ASAP7_75t_L g1422 ( 
.A1(n_1370),
.A2(n_1316),
.B(n_1268),
.C(n_1340),
.Y(n_1422)
);

NOR4xp25_ASAP7_75t_SL g1423 ( 
.A(n_1402),
.B(n_1336),
.C(n_1288),
.D(n_1290),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1399),
.Y(n_1424)
);

INVx5_ASAP7_75t_L g1425 ( 
.A(n_1349),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1390),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1362),
.B(n_1308),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1367),
.A2(n_1305),
.B1(n_1259),
.B2(n_1266),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1343),
.B(n_1352),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1375),
.B(n_1259),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1349),
.B(n_1338),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1401),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1343),
.B(n_1317),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1376),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1375),
.B(n_1266),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1342),
.B(n_1338),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1352),
.B(n_1285),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1374),
.B(n_1285),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1400),
.B(n_1285),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1400),
.B(n_1256),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1342),
.B(n_1305),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1387),
.B(n_1355),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1368),
.Y(n_1443)
);

NOR2x1_ASAP7_75t_L g1444 ( 
.A(n_1361),
.B(n_1358),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1429),
.B(n_1347),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1422),
.B(n_1370),
.C(n_1402),
.Y(n_1446)
);

AOI211xp5_ASAP7_75t_L g1447 ( 
.A1(n_1422),
.A2(n_1410),
.B(n_1408),
.C(n_1360),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1429),
.B(n_1347),
.Y(n_1448)
);

NOR3xp33_ASAP7_75t_L g1449 ( 
.A(n_1410),
.B(n_1392),
.C(n_1348),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1413),
.B(n_1368),
.Y(n_1450)
);

NOR3xp33_ASAP7_75t_SL g1451 ( 
.A(n_1411),
.B(n_1336),
.C(n_1288),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1408),
.B(n_1360),
.C(n_1377),
.Y(n_1452)
);

OAI221xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1428),
.A2(n_1357),
.B1(n_1371),
.B2(n_1361),
.C(n_1386),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1419),
.B(n_1386),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1424),
.B(n_1359),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1423),
.B(n_1330),
.Y(n_1456)
);

OAI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1411),
.A2(n_1421),
.B1(n_1441),
.B2(n_1393),
.C(n_1348),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_SL g1458 ( 
.A(n_1425),
.B(n_1358),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1424),
.B(n_1366),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1409),
.B(n_1372),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1441),
.A2(n_1367),
.B1(n_1371),
.B2(n_1355),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1434),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1421),
.A2(n_1363),
.B1(n_1378),
.B2(n_1392),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1433),
.B(n_1395),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1437),
.A2(n_1381),
.B1(n_1363),
.B2(n_1378),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1433),
.B(n_1381),
.Y(n_1466)
);

NAND4xp25_ASAP7_75t_L g1467 ( 
.A(n_1427),
.B(n_1383),
.C(n_1394),
.D(n_1398),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1437),
.B(n_1372),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1430),
.B(n_1405),
.C(n_1383),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1416),
.A2(n_1388),
.B(n_1345),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1430),
.B(n_1382),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1443),
.B(n_1372),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1435),
.B(n_1382),
.Y(n_1473)
);

NAND4xp25_ASAP7_75t_L g1474 ( 
.A(n_1435),
.B(n_1396),
.C(n_1394),
.D(n_1398),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1439),
.B(n_1372),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1440),
.B(n_1380),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1440),
.B(n_1350),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1414),
.A2(n_1363),
.B1(n_1378),
.B2(n_1387),
.Y(n_1478)
);

AOI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1417),
.A2(n_1397),
.B1(n_1385),
.B2(n_1389),
.C(n_1396),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1436),
.B(n_1385),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1431),
.A2(n_1289),
.B(n_1365),
.Y(n_1481)
);

OAI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1436),
.A2(n_1407),
.B1(n_1404),
.B2(n_1406),
.C(n_1384),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_SL g1483 ( 
.A(n_1423),
.B(n_1270),
.C(n_1324),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1414),
.A2(n_1389),
.B1(n_1346),
.B2(n_1403),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1460),
.B(n_1412),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1462),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1480),
.B(n_1417),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1477),
.B(n_1420),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1470),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1462),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1470),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1460),
.B(n_1416),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1457),
.B(n_1438),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1471),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1470),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1475),
.B(n_1432),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1475),
.B(n_1468),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1472),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1468),
.B(n_1432),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1470),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1477),
.Y(n_1501)
);

INVxp67_ASAP7_75t_SL g1502 ( 
.A(n_1469),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1482),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1420),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1450),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1445),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1469),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1448),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1458),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_1484),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1484),
.Y(n_1511)
);

AND2x4_ASAP7_75t_SL g1512 ( 
.A(n_1449),
.B(n_1442),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1455),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1459),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1479),
.B(n_1426),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1509),
.B(n_1425),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1490),
.Y(n_1517)
);

AOI211xp5_ASAP7_75t_L g1518 ( 
.A1(n_1503),
.A2(n_1446),
.B(n_1447),
.C(n_1452),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1503),
.A2(n_1446),
.B(n_1447),
.C(n_1507),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1490),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1514),
.B(n_1454),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1502),
.B(n_1467),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1485),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_L g1524 ( 
.A(n_1507),
.B(n_1444),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1514),
.B(n_1273),
.Y(n_1525)
);

NOR2x1p5_ASAP7_75t_SL g1526 ( 
.A(n_1491),
.B(n_1418),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1502),
.B(n_1467),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1507),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1507),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1497),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1510),
.B(n_1476),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1511),
.B(n_1476),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1490),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1490),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1501),
.B(n_1425),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1486),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1425),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1493),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1491),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1497),
.B(n_1425),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1499),
.B(n_1474),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1511),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1503),
.B(n_1466),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1513),
.B(n_1273),
.Y(n_1546)
);

INVxp67_ASAP7_75t_SL g1547 ( 
.A(n_1503),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1504),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1494),
.B(n_1474),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1487),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1497),
.B(n_1425),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1505),
.B(n_1425),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1529),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1537),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1547),
.B(n_1493),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1537),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1540),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1540),
.Y(n_1559)
);

INVx3_ASAP7_75t_SL g1560 ( 
.A(n_1516),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1517),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1539),
.B(n_1513),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1519),
.B(n_1509),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1517),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1517),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1528),
.B(n_1498),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1535),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1535),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1535),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1520),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1518),
.B(n_1506),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1523),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1524),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1518),
.A2(n_1515),
.B(n_1452),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1521),
.A2(n_1456),
.B1(n_1483),
.B2(n_1461),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1545),
.B(n_1522),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1520),
.Y(n_1577)
);

INVxp67_ASAP7_75t_SL g1578 ( 
.A(n_1524),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1530),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1522),
.B(n_1515),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1530),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1527),
.B(n_1492),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1545),
.B(n_1506),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1534),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1534),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1549),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1529),
.A2(n_1453),
.B1(n_1489),
.B2(n_1509),
.Y(n_1587)
);

AOI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1527),
.A2(n_1551),
.B1(n_1550),
.B2(n_1549),
.C(n_1544),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1544),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1542),
.B(n_1498),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1542),
.B(n_1496),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1552),
.B(n_1496),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_L g1593 ( 
.A(n_1525),
.B(n_1509),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1531),
.B(n_1508),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1531),
.B(n_1508),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1552),
.B(n_1496),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1593),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1574),
.A2(n_1551),
.B1(n_1550),
.B2(n_1548),
.C(n_1489),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1586),
.B(n_1546),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1563),
.B(n_1275),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1571),
.B(n_1593),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1556),
.B(n_1532),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1523),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1560),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1572),
.A2(n_1541),
.B(n_1523),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1555),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1582),
.B(n_1543),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1555),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1561),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1554),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1563),
.A2(n_1516),
.B1(n_1509),
.B2(n_1512),
.Y(n_1612)
);

AND3x1_ASAP7_75t_L g1613 ( 
.A(n_1575),
.B(n_1451),
.C(n_1458),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1562),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1557),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1560),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1573),
.B(n_1516),
.Y(n_1617)
);

AND2x4_ASAP7_75t_SL g1618 ( 
.A(n_1566),
.B(n_1516),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1564),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1566),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1572),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1532),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1583),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1587),
.A2(n_1481),
.B(n_1543),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1557),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1589),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1578),
.B(n_1526),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1591),
.B(n_1523),
.Y(n_1628)
);

NOR3xp33_ASAP7_75t_SL g1629 ( 
.A(n_1588),
.B(n_1595),
.C(n_1594),
.Y(n_1629)
);

NAND2x1_ASAP7_75t_SL g1630 ( 
.A(n_1572),
.B(n_1553),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1558),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1558),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1611),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1613),
.A2(n_1575),
.B1(n_1580),
.B2(n_1582),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1618),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1620),
.B(n_1591),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1626),
.Y(n_1637)
);

OAI22xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1602),
.A2(n_1580),
.B1(n_1587),
.B2(n_1579),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1607),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1629),
.A2(n_1589),
.B(n_1559),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1602),
.A2(n_1624),
.B1(n_1597),
.B2(n_1623),
.Y(n_1641)
);

AOI32xp33_ASAP7_75t_L g1642 ( 
.A1(n_1613),
.A2(n_1590),
.A3(n_1579),
.B1(n_1581),
.B2(n_1512),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1614),
.B(n_1596),
.Y(n_1643)
);

AOI322xp5_ASAP7_75t_L g1644 ( 
.A1(n_1599),
.A2(n_1581),
.A3(n_1592),
.B1(n_1596),
.B2(n_1590),
.C1(n_1489),
.C2(n_1488),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1612),
.A2(n_1600),
.B(n_1601),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

OAI322xp33_ASAP7_75t_L g1647 ( 
.A1(n_1608),
.A2(n_1559),
.A3(n_1585),
.B1(n_1584),
.B2(n_1570),
.C1(n_1577),
.C2(n_1569),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1618),
.Y(n_1648)
);

OAI322xp33_ASAP7_75t_L g1649 ( 
.A1(n_1608),
.A2(n_1585),
.A3(n_1584),
.B1(n_1577),
.B2(n_1570),
.C1(n_1568),
.C2(n_1569),
.Y(n_1649)
);

OAI31xp33_ASAP7_75t_L g1650 ( 
.A1(n_1622),
.A2(n_1512),
.A3(n_1553),
.B(n_1592),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1616),
.B(n_1572),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1607),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1609),
.Y(n_1653)
);

OAI32xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1603),
.A2(n_1533),
.A3(n_1568),
.B1(n_1565),
.B2(n_1564),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1616),
.A2(n_1512),
.B1(n_1533),
.B2(n_1488),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1609),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1494),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1635),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1635),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1651),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1639),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1617),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1646),
.B(n_1633),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1641),
.B(n_1617),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1637),
.B(n_1615),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1651),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1652),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1636),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1648),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1653),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1645),
.B(n_1275),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1656),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1640),
.B(n_1617),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1643),
.B(n_1617),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1638),
.B(n_1627),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1641),
.B(n_1615),
.Y(n_1676)
);

AO21x1_ASAP7_75t_L g1677 ( 
.A1(n_1675),
.A2(n_1634),
.B(n_1627),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1676),
.A2(n_1671),
.B(n_1664),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1659),
.A2(n_1669),
.B(n_1662),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1663),
.A2(n_1654),
.B1(n_1647),
.B2(n_1649),
.C(n_1642),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1673),
.A2(n_1650),
.B1(n_1655),
.B2(n_1657),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1673),
.B(n_1644),
.Y(n_1682)
);

AOI211xp5_ASAP7_75t_L g1683 ( 
.A1(n_1668),
.A2(n_1604),
.B(n_1627),
.C(n_1625),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1658),
.B(n_1625),
.Y(n_1684)
);

NOR3x1_ASAP7_75t_L g1685 ( 
.A(n_1665),
.B(n_1621),
.C(n_1631),
.Y(n_1685)
);

NAND4xp75_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1604),
.C(n_1621),
.D(n_1632),
.Y(n_1686)
);

NOR2xp67_ASAP7_75t_L g1687 ( 
.A(n_1660),
.B(n_1627),
.Y(n_1687)
);

AOI22x1_ASAP7_75t_L g1688 ( 
.A1(n_1678),
.A2(n_1666),
.B1(n_1660),
.B2(n_1674),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1677),
.A2(n_1670),
.B(n_1672),
.C(n_1667),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1679),
.B(n_1674),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1685),
.B(n_1666),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1681),
.B(n_1660),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1682),
.B(n_1665),
.Y(n_1693)
);

AOI211x1_ASAP7_75t_L g1694 ( 
.A1(n_1684),
.A2(n_1672),
.B(n_1670),
.C(n_1667),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1683),
.B(n_1687),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1680),
.B(n_1661),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1686),
.B(n_1661),
.Y(n_1697)
);

NAND5xp2_ASAP7_75t_L g1698 ( 
.A(n_1693),
.B(n_1632),
.C(n_1631),
.D(n_1628),
.E(n_1481),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_SL g1699 ( 
.A(n_1696),
.B(n_1324),
.C(n_1630),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1689),
.A2(n_1619),
.B1(n_1610),
.B2(n_1598),
.C(n_1628),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1691),
.Y(n_1701)
);

NAND5xp2_ASAP7_75t_L g1702 ( 
.A(n_1692),
.B(n_1465),
.C(n_1478),
.D(n_1289),
.E(n_1630),
.Y(n_1702)
);

OAI211xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1689),
.A2(n_1697),
.B(n_1688),
.C(n_1690),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1701),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1703),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1700),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1698),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1699),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1702),
.Y(n_1709)
);

NAND5xp2_ASAP7_75t_L g1710 ( 
.A(n_1708),
.B(n_1695),
.C(n_1694),
.D(n_1311),
.E(n_1270),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1704),
.Y(n_1711)
);

NOR2xp67_ASAP7_75t_L g1712 ( 
.A(n_1705),
.B(n_1619),
.Y(n_1712)
);

OAI311xp33_ASAP7_75t_L g1713 ( 
.A1(n_1706),
.A2(n_1536),
.A3(n_1538),
.B1(n_1606),
.C1(n_1487),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1707),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1714),
.Y(n_1715)
);

AND2x2_ASAP7_75t_SL g1716 ( 
.A(n_1714),
.B(n_1709),
.Y(n_1716)
);

NOR2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1710),
.B(n_1598),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1715),
.A2(n_1711),
.B1(n_1712),
.B2(n_1610),
.Y(n_1718)
);

NAND4xp25_ASAP7_75t_L g1719 ( 
.A(n_1718),
.B(n_1716),
.C(n_1717),
.D(n_1713),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1567),
.B1(n_1565),
.B2(n_1541),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1719),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1721),
.B(n_1239),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1720),
.A2(n_1606),
.B(n_1567),
.Y(n_1723)
);

INVxp33_ASAP7_75t_L g1724 ( 
.A(n_1723),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1722),
.A2(n_1541),
.B1(n_1536),
.B2(n_1538),
.C(n_1500),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1724),
.A2(n_1725),
.B(n_1415),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1726),
.Y(n_1727)
);

AOI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1727),
.A2(n_1495),
.B1(n_1491),
.B2(n_1500),
.C(n_1463),
.Y(n_1728)
);

AOI211xp5_ASAP7_75t_L g1729 ( 
.A1(n_1728),
.A2(n_1256),
.B(n_1335),
.C(n_1491),
.Y(n_1729)
);


endmodule