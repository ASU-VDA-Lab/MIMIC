module fake_jpeg_26504_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AND2x4_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_5),
.Y(n_6)
);

BUFx10_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx11_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_0),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_15),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_L g16 ( 
.A1(n_6),
.A2(n_12),
.B1(n_9),
.B2(n_8),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_6),
.B1(n_9),
.B2(n_8),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_29),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_14),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_19),
.C(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_25),
.B1(n_21),
.B2(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_11),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_7),
.B(n_11),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_34),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_39),
.B1(n_2),
.B2(n_4),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_25),
.B1(n_17),
.B2(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_36),
.B(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_39),
.Y(n_44)
);


endmodule