module fake_ibex_926_n_1186 (n_151, n_147, n_85, n_167, n_128, n_208, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_224, n_183, n_67, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_214, n_79, n_81, n_35, n_159, n_202, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_228, n_1186);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_224;
input n_183;
input n_67;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_214;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;
input n_228;

output n_1186;

wire n_1084;
wire n_599;
wire n_822;
wire n_778;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1104;
wire n_1011;
wire n_992;
wire n_1148;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_1110;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_1182;
wire n_926;
wire n_1097;
wire n_1079;
wire n_1031;
wire n_1143;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_845;
wire n_972;
wire n_1100;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_1162;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_1125;
wire n_634;
wire n_733;
wire n_991;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_930;
wire n_336;
wire n_1018;
wire n_258;
wire n_861;
wire n_959;
wire n_1106;
wire n_1044;
wire n_1129;
wire n_449;
wire n_1138;
wire n_547;
wire n_1134;
wire n_727;
wire n_1131;
wire n_1077;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_1174;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_1147;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_1098;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_317;
wire n_375;
wire n_340;
wire n_280;
wire n_708;
wire n_901;
wire n_1096;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_1166;
wire n_1181;
wire n_1140;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_1144;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_348;
wire n_1109;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1112;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_1172;
wire n_1099;
wire n_598;
wire n_825;
wire n_740;
wire n_1169;
wire n_386;
wire n_549;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_1055;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_1103;
wire n_1161;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1177;
wire n_1068;
wire n_496;
wire n_301;
wire n_325;
wire n_617;
wire n_434;
wire n_1184;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_1141;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_1168;
wire n_289;
wire n_716;
wire n_865;
wire n_1130;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_1179;
wire n_933;
wire n_1081;
wire n_1153;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_1155;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_1117;
wire n_1101;
wire n_518;
wire n_367;
wire n_1052;
wire n_852;
wire n_789;
wire n_1133;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_1178;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_1116;
wire n_623;
wire n_585;
wire n_1030;
wire n_1094;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_1082;
wire n_1137;
wire n_660;
wire n_524;
wire n_349;
wire n_849;
wire n_765;
wire n_857;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_1120;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_1180;
wire n_619;
wire n_1089;
wire n_536;
wire n_1124;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_922;
wire n_1171;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_1183;
wire n_253;
wire n_234;
wire n_300;
wire n_1151;
wire n_1135;
wire n_973;
wire n_1146;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_1038;
wire n_1092;
wire n_999;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1142;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1173;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_433;
wire n_439;
wire n_299;
wire n_704;
wire n_1126;
wire n_1007;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_1063;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_1115;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_553;
wire n_554;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_955;
wire n_1170;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_1057;
wire n_1049;
wire n_763;
wire n_1086;
wire n_745;
wire n_1158;
wire n_329;
wire n_1149;
wire n_447;
wire n_1176;
wire n_940;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_1160;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_1033;
wire n_1118;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_1114;
wire n_409;
wire n_1093;
wire n_582;
wire n_978;
wire n_818;
wire n_1167;
wire n_653;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_744;
wire n_817;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_1107;
wire n_381;
wire n_1073;
wire n_1108;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_1111;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_1128;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_440;
wire n_268;
wire n_858;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_729;
wire n_430;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_1145;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_1113;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_1164;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_866;
wire n_958;
wire n_1175;
wire n_485;
wire n_1139;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_1159;
wire n_1119;
wire n_903;
wire n_1154;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_1095;
wire n_455;
wire n_1136;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_1091;
wire n_885;
wire n_588;
wire n_513;
wire n_877;
wire n_1121;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_528;
wire n_1005;
wire n_1102;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_1150;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_1165;
wire n_1185;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_1122;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_912;
wire n_921;
wire n_890;
wire n_1058;
wire n_1105;
wire n_1163;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_1123;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_231;
wire n_298;
wire n_587;
wire n_1035;
wire n_760;
wire n_1157;
wire n_751;
wire n_806;
wire n_1127;
wire n_932;
wire n_657;
wire n_764;
wire n_1156;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_947;
wire n_559;
wire n_425;
wire n_1050;

INVx1_ASAP7_75t_L g229 ( 
.A(n_34),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_94),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_147),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_109),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_77),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_150),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_99),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_81),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_L g242 ( 
.A(n_103),
.B(n_32),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_151),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_142),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_167),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_111),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_2),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_86),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_47),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_53),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_194),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_149),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_202),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_1),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_32),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_18),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_41),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_47),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_118),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_132),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_186),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_207),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_9),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_12),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_164),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_218),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_58),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_155),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_213),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_180),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_126),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_8),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_189),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_146),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_152),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_82),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_166),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_80),
.B(n_160),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_188),
.B(n_135),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_88),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_179),
.B(n_105),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_136),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_12),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_162),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_181),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_191),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_217),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_204),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_42),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_156),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_192),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_125),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_107),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_39),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_90),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_84),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_115),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_177),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_168),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_3),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_139),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_48),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_123),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_44),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_54),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_221),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_144),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_128),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_35),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_101),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_52),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_226),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_159),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_210),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_120),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_193),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_65),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_17),
.B(n_97),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_28),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_104),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_93),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_1),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_165),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_190),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_170),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_53),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_176),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_31),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_169),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_117),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_0),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_110),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_48),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_178),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_214),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_201),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_209),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_108),
.Y(n_346)
);

BUFx2_ASAP7_75t_SL g347 ( 
.A(n_24),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_76),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_175),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_24),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_141),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_143),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_73),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_112),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_92),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_5),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_183),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_38),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_26),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_49),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_0),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_196),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_161),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_74),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_6),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_33),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_130),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_174),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_51),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_7),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_13),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_95),
.Y(n_372)
);

BUFx8_ASAP7_75t_SL g373 ( 
.A(n_223),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_200),
.B(n_11),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_129),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_28),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_133),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_58),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_66),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_46),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_71),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_91),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_79),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_89),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_41),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_220),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_57),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_114),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_208),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_17),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_87),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_67),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_96),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_57),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_172),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_336),
.B(n_2),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_276),
.Y(n_397)
);

OAI22xp33_ASAP7_75t_L g398 ( 
.A1(n_273),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_308),
.B(n_6),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_310),
.Y(n_400)
);

XNOR2x2_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_7),
.Y(n_401)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_243),
.A2(n_113),
.B(n_227),
.Y(n_402)
);

BUFx12f_ASAP7_75t_L g403 ( 
.A(n_284),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_276),
.Y(n_404)
);

OAI21x1_ASAP7_75t_L g405 ( 
.A1(n_243),
.A2(n_106),
.B(n_224),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_276),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_394),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_8),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_394),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_394),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_9),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

CKINVDCx11_ASAP7_75t_R g418 ( 
.A(n_369),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_233),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g420 ( 
.A1(n_254),
.A2(n_116),
.B(n_222),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_251),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_373),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_251),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_302),
.B(n_10),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_248),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_306),
.Y(n_427)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_276),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g429 ( 
.A(n_316),
.B(n_64),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_229),
.B(n_10),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_256),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_257),
.B(n_11),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_14),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_270),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_376),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_344),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_317),
.Y(n_437)
);

OAI22x1_ASAP7_75t_SL g438 ( 
.A1(n_369),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_254),
.A2(n_122),
.B(n_219),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_327),
.B(n_15),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_316),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_282),
.Y(n_445)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_344),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_371),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_373),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_250),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_232),
.B(n_68),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_259),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_334),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

INVx5_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_260),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_360),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_262),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_321),
.B(n_282),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_365),
.B(n_19),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_395),
.B(n_19),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_370),
.B(n_20),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_283),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_283),
.Y(n_475)
);

OAI22x1_ASAP7_75t_SL g476 ( 
.A1(n_249),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_301),
.B(n_22),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_230),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_333),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_234),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_231),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_285),
.A2(n_375),
.B1(n_269),
.B2(n_279),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_321),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_347),
.B(n_23),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_337),
.B(n_23),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_236),
.Y(n_486)
);

INVx5_ASAP7_75t_L g487 ( 
.A(n_353),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_353),
.B(n_69),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_237),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_363),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_363),
.B(n_25),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_238),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_285),
.B(n_26),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_375),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_239),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_245),
.B(n_27),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_287),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_266),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_291),
.B(n_27),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_449),
.Y(n_500)
);

INVx8_ASAP7_75t_L g501 ( 
.A(n_494),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

OAI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_484),
.A2(n_297),
.B1(n_313),
.B2(n_312),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_485),
.B(n_253),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_415),
.B(n_241),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_425),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_429),
.B(n_488),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_494),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_406),
.B(n_242),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_451),
.Y(n_512)
);

AO21x2_ASAP7_75t_L g513 ( 
.A1(n_405),
.A2(n_261),
.B(n_258),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_492),
.B(n_496),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_492),
.B(n_264),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_451),
.B(n_319),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_460),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_411),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_422),
.Y(n_519)
);

AND3x2_ASAP7_75t_L g520 ( 
.A(n_450),
.B(n_298),
.C(n_374),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_404),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_400),
.Y(n_522)
);

AND3x2_ASAP7_75t_L g523 ( 
.A(n_467),
.B(n_289),
.C(n_278),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_426),
.B(n_249),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_419),
.B(n_330),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_426),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_339),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_417),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_432),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_462),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_492),
.B(n_292),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_462),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_464),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_492),
.B(n_293),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_464),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_468),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_419),
.B(n_294),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_496),
.B(n_300),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_424),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_468),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_416),
.Y(n_548)
);

BUFx6f_ASAP7_75t_SL g549 ( 
.A(n_435),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_445),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_445),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_471),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_478),
.B(n_303),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_471),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_475),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_481),
.B(n_304),
.Y(n_557)
);

NOR2x1p5_ASAP7_75t_L g558 ( 
.A(n_403),
.B(n_350),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_479),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_480),
.B(n_309),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_490),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_429),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_L g563 ( 
.A(n_429),
.B(n_286),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_407),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_436),
.Y(n_565)
);

AND3x2_ASAP7_75t_L g566 ( 
.A(n_422),
.B(n_325),
.C(n_323),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_436),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_436),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_436),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_498),
.Y(n_570)
);

INVx8_ASAP7_75t_L g571 ( 
.A(n_403),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_429),
.B(n_235),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_486),
.B(n_356),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_431),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_448),
.B(n_311),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_448),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_429),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_434),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_437),
.Y(n_579)
);

BUFx4f_ASAP7_75t_L g580 ( 
.A(n_493),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_442),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_489),
.B(n_329),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_495),
.B(n_331),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_418),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_488),
.B(n_240),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_487),
.B(n_332),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_452),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_456),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_396),
.B(n_366),
.C(n_361),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_427),
.B(n_378),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_427),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_487),
.B(n_340),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_453),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_453),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_499),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_453),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_409),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_412),
.B(n_342),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_457),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_461),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_SL g602 ( 
.A(n_433),
.B(n_311),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_457),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_470),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_487),
.B(n_444),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_457),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_472),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_458),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_458),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_482),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g612 ( 
.A1(n_402),
.A2(n_351),
.B(n_346),
.Y(n_612)
);

AO21x2_ASAP7_75t_L g613 ( 
.A1(n_477),
.A2(n_491),
.B(n_440),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_458),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_421),
.B(n_244),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_497),
.B(n_367),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_423),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_458),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_418),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_487),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_488),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_399),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_465),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_465),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_463),
.Y(n_625)
);

BUFx6f_ASAP7_75t_SL g626 ( 
.A(n_488),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_476),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_447),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_441),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_466),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_488),
.B(n_246),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_441),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_517),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_603),
.B(n_247),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_613),
.B(n_420),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_571),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_577),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_599),
.A2(n_622),
.B1(n_512),
.B2(n_536),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_599),
.B(n_252),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_617),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_621),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_548),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_615),
.B(n_255),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_580),
.B(n_263),
.Y(n_644)
);

CKINVDCx6p67_ASAP7_75t_R g645 ( 
.A(n_571),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_580),
.B(n_265),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_584),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_574),
.B(n_267),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_550),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_552),
.Y(n_650)
);

OR2x6_ASAP7_75t_SL g651 ( 
.A(n_627),
.B(n_438),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_578),
.B(n_579),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_553),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_587),
.B(n_588),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_519),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_500),
.B(n_268),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_595),
.B(n_271),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_555),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_538),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_601),
.B(n_272),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_598),
.B(n_315),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_531),
.B(n_532),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_556),
.Y(n_663)
);

NOR2x1p5_ASAP7_75t_L g664 ( 
.A(n_516),
.B(n_401),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_605),
.B(n_439),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_509),
.B(n_318),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_596),
.B(n_318),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_563),
.B(n_439),
.C(n_392),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_591),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_608),
.B(n_274),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_619),
.B(n_528),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_535),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_539),
.B(n_275),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_591),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_589),
.B(n_443),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_573),
.B(n_277),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_541),
.B(n_280),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_576),
.B(n_398),
.Y(n_678)
);

INVxp33_ASAP7_75t_L g679 ( 
.A(n_524),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_542),
.B(n_281),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_543),
.B(n_288),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_543),
.B(n_290),
.Y(n_682)
);

AND3x4_ASAP7_75t_L g683 ( 
.A(n_584),
.B(n_326),
.C(n_398),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_602),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_551),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_560),
.B(n_295),
.Y(n_686)
);

INVxp67_ASAP7_75t_SL g687 ( 
.A(n_563),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_560),
.B(n_296),
.Y(n_688)
);

INVxp33_ASAP7_75t_L g689 ( 
.A(n_575),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_559),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_505),
.B(n_526),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_505),
.B(n_299),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_570),
.B(n_305),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_544),
.B(n_590),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_561),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_522),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_508),
.B(n_320),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_547),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_506),
.B(n_307),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_551),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_544),
.B(n_314),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_519),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_504),
.B(n_324),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_510),
.B(n_328),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_501),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_514),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_504),
.B(n_335),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_611),
.A2(n_322),
.B1(n_343),
.B2(n_345),
.Y(n_708)
);

NOR2x1p5_ASAP7_75t_L g709 ( 
.A(n_558),
.B(n_343),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_510),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_510),
.B(n_338),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_508),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_SL g713 ( 
.A(n_549),
.B(n_345),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_616),
.B(n_455),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_602),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_554),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_557),
.Y(n_717)
);

NAND2x1p5_ASAP7_75t_L g718 ( 
.A(n_557),
.B(n_455),
.Y(n_718)
);

BUFx6f_ASAP7_75t_SL g719 ( 
.A(n_628),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_503),
.B(n_348),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_582),
.B(n_349),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_582),
.B(n_352),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_583),
.B(n_354),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_583),
.B(n_364),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_501),
.A2(n_362),
.B1(n_377),
.B2(n_384),
.Y(n_725)
);

BUFx12f_ASAP7_75t_SL g726 ( 
.A(n_549),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_625),
.B(n_368),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_SL g728 ( 
.A1(n_523),
.A2(n_362),
.B1(n_377),
.B2(n_372),
.Y(n_728)
);

BUFx6f_ASAP7_75t_SL g729 ( 
.A(n_501),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_616),
.B(n_382),
.C(n_383),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_566),
.B(n_586),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_606),
.B(n_29),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_566),
.B(n_388),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_586),
.B(n_391),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_620),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_520),
.B(n_393),
.Y(n_736)
);

AND2x6_ASAP7_75t_SL g737 ( 
.A(n_520),
.B(n_30),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_620),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_585),
.B(n_397),
.Y(n_739)
);

AND2x2_ASAP7_75t_SL g740 ( 
.A(n_572),
.B(n_30),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_592),
.B(n_397),
.Y(n_741)
);

AO221x1_ASAP7_75t_L g742 ( 
.A1(n_572),
.A2(n_474),
.B1(n_466),
.B2(n_34),
.C(n_35),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_631),
.B(n_397),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_507),
.A2(n_446),
.B1(n_473),
.B2(n_454),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_515),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_626),
.B(n_631),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_515),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_635),
.A2(n_507),
.B(n_513),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_691),
.B(n_672),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_635),
.A2(n_540),
.B(n_537),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_698),
.B(n_502),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_687),
.A2(n_525),
.B1(n_529),
.B2(n_533),
.Y(n_752)
);

BUFx4f_ASAP7_75t_L g753 ( 
.A(n_645),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_668),
.A2(n_612),
.B(n_511),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_642),
.A2(n_525),
.B(n_546),
.C(n_545),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_726),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_729),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_696),
.Y(n_758)
);

BUFx8_ASAP7_75t_L g759 ( 
.A(n_729),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_652),
.B(n_518),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_665),
.A2(n_533),
.B(n_530),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_654),
.B(n_534),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_640),
.B(n_534),
.Y(n_763)
);

NOR2x1_ASAP7_75t_L g764 ( 
.A(n_636),
.B(n_629),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_659),
.B(n_632),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_740),
.A2(n_446),
.B1(n_428),
.B2(n_454),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_670),
.B(n_33),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_670),
.B(n_36),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_633),
.B(n_36),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_662),
.B(n_37),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_694),
.B(n_710),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_735),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_638),
.B(n_37),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_716),
.A2(n_597),
.B(n_564),
.Y(n_774)
);

OAI21xp33_ASAP7_75t_L g775 ( 
.A1(n_678),
.A2(n_466),
.B(n_474),
.Y(n_775)
);

NOR2x2_ASAP7_75t_L g776 ( 
.A(n_725),
.B(n_38),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_717),
.A2(n_600),
.B(n_565),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_715),
.B(n_40),
.Y(n_778)
);

NOR2x1p5_ASAP7_75t_SL g779 ( 
.A(n_685),
.B(n_565),
.Y(n_779)
);

AO22x1_ASAP7_75t_L g780 ( 
.A1(n_689),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_649),
.A2(n_474),
.B(n_473),
.C(n_623),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_738),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_738),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_699),
.B(n_43),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_712),
.B(n_44),
.Y(n_785)
);

AO21x1_ASAP7_75t_L g786 ( 
.A1(n_732),
.A2(n_609),
.B(n_567),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_737),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_650),
.A2(n_597),
.B(n_568),
.C(n_623),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_653),
.A2(n_594),
.B(n_569),
.C(n_618),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_637),
.B(n_521),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_667),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_708),
.A2(n_666),
.B1(n_661),
.B2(n_684),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_699),
.B(n_45),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_637),
.B(n_521),
.Y(n_794)
);

AO21x1_ASAP7_75t_L g795 ( 
.A1(n_739),
.A2(n_581),
.B(n_604),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_697),
.B(n_45),
.Y(n_796)
);

AO21x1_ASAP7_75t_L g797 ( 
.A1(n_743),
.A2(n_581),
.B(n_607),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_658),
.A2(n_610),
.B(n_609),
.C(n_618),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_666),
.B(n_46),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_639),
.B(n_50),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_655),
.Y(n_801)
);

OAI21xp33_ASAP7_75t_L g802 ( 
.A1(n_679),
.A2(n_630),
.B(n_624),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_721),
.B(n_722),
.Y(n_803)
);

AOI211xp5_ASAP7_75t_L g804 ( 
.A1(n_728),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_671),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_681),
.B(n_54),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_702),
.B(n_55),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_664),
.B(n_55),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_713),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_682),
.B(n_56),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_686),
.B(n_56),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_720),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_675),
.B(n_59),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_663),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_688),
.B(n_61),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_704),
.B(n_62),
.Y(n_816)
);

AO21x1_ASAP7_75t_L g817 ( 
.A1(n_746),
.A2(n_62),
.B(n_63),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_669),
.Y(n_818)
);

BUFx2_ASAP7_75t_L g819 ( 
.A(n_647),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_745),
.A2(n_614),
.B(n_593),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_709),
.B(n_70),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_634),
.B(n_72),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_674),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_690),
.A2(n_228),
.B(n_78),
.C(n_83),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_648),
.A2(n_75),
.B(n_85),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_706),
.A2(n_742),
.B1(n_730),
.B2(n_736),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_657),
.A2(n_98),
.B(n_100),
.Y(n_827)
);

OAI21xp33_ASAP7_75t_L g828 ( 
.A1(n_692),
.A2(n_102),
.B(n_119),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_747),
.B(n_121),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_711),
.B(n_124),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_660),
.A2(n_127),
.B(n_131),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_733),
.B(n_216),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_695),
.A2(n_138),
.B(n_140),
.Y(n_833)
);

AND2x4_ASAP7_75t_L g834 ( 
.A(n_656),
.B(n_215),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_676),
.B(n_643),
.Y(n_835)
);

INVx11_ASAP7_75t_L g836 ( 
.A(n_719),
.Y(n_836)
);

O2A1O1Ixp5_ASAP7_75t_L g837 ( 
.A1(n_723),
.A2(n_724),
.B(n_734),
.C(n_741),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_641),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_673),
.B(n_148),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_677),
.B(n_154),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_680),
.B(n_157),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_731),
.A2(n_163),
.B(n_171),
.C(n_173),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_719),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_701),
.A2(n_714),
.B(n_703),
.C(n_707),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_693),
.B(n_212),
.Y(n_845)
);

INVx5_ASAP7_75t_L g846 ( 
.A(n_641),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_727),
.A2(n_646),
.B(n_644),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_700),
.A2(n_184),
.B(n_185),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_718),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_744),
.A2(n_195),
.B(n_197),
.C(n_198),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_758),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_748),
.A2(n_754),
.B(n_803),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_759),
.Y(n_853)
);

CKINVDCx6p67_ASAP7_75t_R g854 ( 
.A(n_757),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_805),
.B(n_683),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_761),
.A2(n_750),
.B(n_835),
.Y(n_856)
);

INVx6_ASAP7_75t_SL g857 ( 
.A(n_785),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_763),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_791),
.B(n_651),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_753),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_799),
.B(n_203),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_755),
.A2(n_844),
.B(n_752),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_773),
.B(n_771),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_792),
.B(n_807),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_796),
.B(n_762),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_785),
.B(n_787),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_838),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_785),
.B(n_757),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_819),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_751),
.A2(n_766),
.B1(n_826),
.B2(n_793),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_784),
.A2(n_811),
.B1(n_810),
.B2(n_806),
.Y(n_871)
);

AO31x2_ASAP7_75t_L g872 ( 
.A1(n_795),
.A2(n_797),
.A3(n_786),
.B(n_817),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_787),
.B(n_801),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_820),
.A2(n_777),
.B(n_774),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_812),
.A2(n_815),
.B(n_816),
.C(n_839),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_759),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_756),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_837),
.A2(n_788),
.B(n_789),
.Y(n_878)
);

INVx5_ASAP7_75t_L g879 ( 
.A(n_843),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_769),
.B(n_834),
.Y(n_880)
);

OAI22x1_ASAP7_75t_L g881 ( 
.A1(n_787),
.A2(n_776),
.B1(n_808),
.B2(n_813),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_846),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_SL g883 ( 
.A(n_809),
.B(n_846),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_770),
.Y(n_884)
);

INVx3_ASAP7_75t_SL g885 ( 
.A(n_813),
.Y(n_885)
);

NOR2x1_ASAP7_75t_R g886 ( 
.A(n_822),
.B(n_836),
.Y(n_886)
);

OAI21x1_ASAP7_75t_L g887 ( 
.A1(n_790),
.A2(n_794),
.B(n_831),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_840),
.A2(n_841),
.B(n_830),
.C(n_824),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_834),
.B(n_822),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_849),
.B(n_772),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_845),
.A2(n_847),
.B(n_798),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_821),
.B(n_804),
.Y(n_892)
);

OAI21x1_ASAP7_75t_L g893 ( 
.A1(n_825),
.A2(n_827),
.B(n_802),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_800),
.B(n_832),
.Y(n_894)
);

AO31x2_ASAP7_75t_L g895 ( 
.A1(n_842),
.A2(n_850),
.A3(n_781),
.B(n_848),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_775),
.A2(n_778),
.B(n_779),
.C(n_828),
.Y(n_896)
);

OAI221xp5_ASAP7_75t_L g897 ( 
.A1(n_804),
.A2(n_764),
.B1(n_765),
.B2(n_823),
.C(n_818),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_782),
.B(n_783),
.Y(n_898)
);

AND2x6_ASAP7_75t_L g899 ( 
.A(n_780),
.B(n_829),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_803),
.A2(n_749),
.B(n_768),
.C(n_767),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_749),
.B(n_805),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_748),
.A2(n_635),
.B(n_563),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_749),
.B(n_805),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_SL g904 ( 
.A1(n_833),
.A2(n_562),
.B(n_687),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_748),
.A2(n_635),
.B(n_563),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_753),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_749),
.B(n_805),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_803),
.A2(n_749),
.B(n_768),
.C(n_767),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_749),
.B(n_603),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_749),
.A2(n_760),
.B1(n_762),
.B2(n_814),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_758),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_805),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_753),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_805),
.B(n_527),
.Y(n_914)
);

AND2x6_ASAP7_75t_L g915 ( 
.A(n_822),
.B(n_834),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_749),
.B(n_805),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_749),
.B(n_705),
.Y(n_917)
);

AO31x2_ASAP7_75t_L g918 ( 
.A1(n_748),
.A2(n_795),
.A3(n_797),
.B(n_786),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_805),
.B(n_633),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_805),
.B(n_622),
.Y(n_920)
);

AOI21xp33_ASAP7_75t_L g921 ( 
.A1(n_749),
.A2(n_679),
.B(n_527),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_803),
.A2(n_749),
.B(n_768),
.C(n_767),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

AO31x2_ASAP7_75t_L g924 ( 
.A1(n_748),
.A2(n_795),
.A3(n_797),
.B(n_786),
.Y(n_924)
);

AND2x2_ASAP7_75t_SL g925 ( 
.A(n_753),
.B(n_524),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_749),
.A2(n_760),
.B1(n_762),
.B2(n_814),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_805),
.A2(n_524),
.B1(n_725),
.B2(n_633),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_749),
.A2(n_760),
.B1(n_762),
.B2(n_814),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_803),
.A2(n_749),
.B(n_768),
.C(n_767),
.Y(n_929)
);

AOI21xp33_ASAP7_75t_L g930 ( 
.A1(n_749),
.A2(n_679),
.B(n_527),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_785),
.Y(n_931)
);

BUFx8_ASAP7_75t_L g932 ( 
.A(n_819),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_749),
.B(n_805),
.Y(n_933)
);

INVx8_ASAP7_75t_L g934 ( 
.A(n_785),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_749),
.B(n_805),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_749),
.B(n_805),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_749),
.B(n_705),
.Y(n_937)
);

BUFx5_ASAP7_75t_L g938 ( 
.A(n_758),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_SL g939 ( 
.A1(n_805),
.A2(n_725),
.B(n_708),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_749),
.B(n_705),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_833),
.A2(n_748),
.B(n_824),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_805),
.A2(n_524),
.B1(n_725),
.B2(n_633),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_759),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_749),
.B(n_805),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_785),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_792),
.A2(n_611),
.B1(n_683),
.B2(n_773),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_753),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_749),
.B(n_805),
.Y(n_948)
);

BUFx2_ASAP7_75t_L g949 ( 
.A(n_857),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_900),
.A2(n_922),
.B(n_908),
.Y(n_950)
);

NOR2x1_ASAP7_75t_R g951 ( 
.A(n_853),
.B(n_943),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_901),
.B(n_903),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_934),
.B(n_868),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_907),
.B(n_916),
.Y(n_954)
);

NAND3xp33_ASAP7_75t_L g955 ( 
.A(n_875),
.B(n_929),
.C(n_862),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_906),
.B(n_945),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_874),
.A2(n_893),
.B(n_887),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_934),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_910),
.A2(n_926),
.B1(n_928),
.B2(n_915),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_932),
.Y(n_960)
);

BUFx2_ASAP7_75t_R g961 ( 
.A(n_877),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_912),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_939),
.B(n_855),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_915),
.A2(n_946),
.B1(n_892),
.B2(n_864),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_851),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_851),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_879),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_857),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_867),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_865),
.Y(n_970)
);

INVx5_ASAP7_75t_SL g971 ( 
.A(n_854),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_868),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_904),
.A2(n_896),
.B(n_871),
.Y(n_973)
);

OR2x6_ASAP7_75t_L g974 ( 
.A(n_876),
.B(n_860),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_911),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_SL g976 ( 
.A(n_945),
.B(n_915),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_891),
.A2(n_856),
.B(n_941),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_915),
.A2(n_925),
.B1(n_881),
.B2(n_863),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_879),
.Y(n_979)
);

BUFx2_ASAP7_75t_R g980 ( 
.A(n_923),
.Y(n_980)
);

INVx6_ASAP7_75t_L g981 ( 
.A(n_932),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_878),
.B(n_870),
.C(n_888),
.Y(n_982)
);

OR2x6_ASAP7_75t_L g983 ( 
.A(n_947),
.B(n_913),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_L g984 ( 
.A1(n_880),
.A2(n_886),
.B(n_889),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_879),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_869),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_933),
.B(n_935),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_882),
.Y(n_988)
);

BUFx4f_ASAP7_75t_L g989 ( 
.A(n_885),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_894),
.A2(n_884),
.B(n_897),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_931),
.B(n_861),
.C(n_927),
.Y(n_991)
);

OA21x2_ASAP7_75t_L g992 ( 
.A1(n_918),
.A2(n_924),
.B(n_872),
.Y(n_992)
);

OA21x2_ASAP7_75t_L g993 ( 
.A1(n_918),
.A2(n_924),
.B(n_872),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_917),
.Y(n_994)
);

NOR2xp67_ASAP7_75t_SL g995 ( 
.A(n_914),
.B(n_920),
.Y(n_995)
);

OA21x2_ASAP7_75t_L g996 ( 
.A1(n_895),
.A2(n_898),
.B(n_909),
.Y(n_996)
);

BUFx12f_ASAP7_75t_L g997 ( 
.A(n_873),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_942),
.A2(n_948),
.B1(n_944),
.B2(n_936),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_866),
.Y(n_999)
);

AO21x2_ASAP7_75t_L g1000 ( 
.A1(n_921),
.A2(n_930),
.B(n_938),
.Y(n_1000)
);

NAND3xp33_ASAP7_75t_L g1001 ( 
.A(n_883),
.B(n_919),
.C(n_937),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_940),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_890),
.B(n_859),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_899),
.B(n_906),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_899),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_L g1006 ( 
.A(n_899),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_900),
.A2(n_922),
.B(n_929),
.C(n_908),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_852),
.A2(n_905),
.B(n_902),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_858),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_906),
.B(n_753),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_901),
.B(n_903),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_900),
.A2(n_922),
.B(n_908),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_906),
.B(n_753),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_901),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_853),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_906),
.B(n_945),
.Y(n_1016)
);

BUFx12f_ASAP7_75t_L g1017 ( 
.A(n_853),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_912),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_900),
.A2(n_922),
.B(n_908),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_900),
.A2(n_922),
.B(n_908),
.Y(n_1020)
);

BUFx2_ASAP7_75t_R g1021 ( 
.A(n_853),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_901),
.B(n_903),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_901),
.B(n_903),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_965),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_962),
.Y(n_1025)
);

BUFx4f_ASAP7_75t_SL g1026 ( 
.A(n_1017),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_966),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_987),
.B(n_970),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_966),
.Y(n_1029)
);

AO21x2_ASAP7_75t_L g1030 ( 
.A1(n_977),
.A2(n_1008),
.B(n_973),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_1018),
.Y(n_1031)
);

INVx5_ASAP7_75t_L g1032 ( 
.A(n_969),
.Y(n_1032)
);

OAI22xp33_ASAP7_75t_SL g1033 ( 
.A1(n_959),
.A2(n_976),
.B1(n_1006),
.B2(n_1009),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1023),
.B(n_952),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_1008),
.A2(n_957),
.B(n_1019),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_SL g1036 ( 
.A(n_1021),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_986),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_954),
.B(n_1011),
.Y(n_1038)
);

AO21x2_ASAP7_75t_L g1039 ( 
.A1(n_950),
.A2(n_1020),
.B(n_1012),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_1015),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_1005),
.B(n_1004),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_975),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_1014),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_997),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_959),
.Y(n_1045)
);

AO21x2_ASAP7_75t_L g1046 ( 
.A1(n_982),
.A2(n_955),
.B(n_1007),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1022),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_998),
.B(n_963),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_980),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1006),
.A2(n_978),
.B1(n_964),
.B2(n_1001),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_L g1051 ( 
.A(n_1010),
.Y(n_1051)
);

BUFx4f_ASAP7_75t_SL g1052 ( 
.A(n_960),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_985),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_996),
.Y(n_1054)
);

BUFx5_ASAP7_75t_L g1055 ( 
.A(n_956),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_1032),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1045),
.A2(n_991),
.B1(n_1001),
.B2(n_995),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_1055),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_1032),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1050),
.A2(n_1016),
.B(n_956),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1055),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1039),
.B(n_992),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1024),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1039),
.B(n_992),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1039),
.B(n_993),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1024),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1045),
.A2(n_972),
.B1(n_991),
.B2(n_953),
.Y(n_1067)
);

OAI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_1048),
.A2(n_990),
.B1(n_984),
.B2(n_976),
.C(n_994),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_1054),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1029),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1034),
.B(n_958),
.Y(n_1071)
);

AND3x1_ASAP7_75t_L g1072 ( 
.A(n_1036),
.B(n_967),
.C(n_979),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1029),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1028),
.B(n_1000),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_1028),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1027),
.B(n_994),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1063),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1075),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1063),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_1075),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_1062),
.B(n_1035),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1066),
.B(n_1047),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1066),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_1069),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1062),
.B(n_1035),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_1056),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_1060),
.B(n_1059),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1067),
.A2(n_1068),
.B1(n_1057),
.B2(n_1033),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1062),
.B(n_1030),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_1076),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_1058),
.Y(n_1091)
);

NAND4xp25_ASAP7_75t_L g1092 ( 
.A(n_1068),
.B(n_1038),
.C(n_1003),
.D(n_1049),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1071),
.B(n_1040),
.Y(n_1093)
);

OAI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1060),
.A2(n_972),
.B1(n_953),
.B2(n_1043),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1077),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1077),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_1087),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1089),
.B(n_1064),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1079),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1082),
.B(n_1070),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1089),
.B(n_1064),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1079),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1085),
.B(n_1064),
.Y(n_1103)
);

NAND4xp25_ASAP7_75t_L g1104 ( 
.A(n_1088),
.B(n_1067),
.C(n_1003),
.D(n_1074),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1078),
.B(n_1073),
.Y(n_1105)
);

AND2x2_ASAP7_75t_SL g1106 ( 
.A(n_1091),
.B(n_1072),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1083),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1080),
.B(n_1090),
.Y(n_1108)
);

OR2x6_ASAP7_75t_L g1109 ( 
.A(n_1087),
.B(n_1086),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1084),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1108),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1096),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1098),
.B(n_1091),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1098),
.B(n_1085),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1096),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1099),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1100),
.B(n_1093),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1101),
.B(n_1065),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1099),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1095),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1102),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_1109),
.B(n_1097),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1101),
.B(n_1074),
.Y(n_1123)
);

NOR3xp33_ASAP7_75t_L g1124 ( 
.A(n_1104),
.B(n_1092),
.C(n_1094),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1109),
.B(n_1086),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1103),
.B(n_1065),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1107),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1112),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1122),
.B(n_1097),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1111),
.B(n_1103),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1115),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1116),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_SL g1133 ( 
.A(n_1125),
.B(n_1106),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1119),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1124),
.A2(n_1106),
.B1(n_1109),
.B2(n_1072),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1113),
.Y(n_1136)
);

AOI21xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1122),
.A2(n_1040),
.B(n_1109),
.Y(n_1137)
);

OAI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_1117),
.A2(n_1126),
.B(n_1118),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1114),
.B(n_1081),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1125),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1118),
.B(n_1081),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1120),
.Y(n_1142)
);

INVxp33_ASAP7_75t_L g1143 ( 
.A(n_1137),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_1135),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1140),
.A2(n_1122),
.B1(n_1136),
.B2(n_1138),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1130),
.A2(n_1126),
.B1(n_1127),
.B2(n_1121),
.C(n_1031),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1133),
.A2(n_1081),
.B1(n_1123),
.B2(n_1110),
.Y(n_1147)
);

OAI32xp33_ASAP7_75t_L g1148 ( 
.A1(n_1140),
.A2(n_1086),
.A3(n_1037),
.B1(n_1059),
.B2(n_1061),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_1129),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1129),
.A2(n_1033),
.B(n_1025),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_SL g1151 ( 
.A(n_1148),
.B(n_951),
.Y(n_1151)
);

XNOR2xp5_ASAP7_75t_L g1152 ( 
.A(n_1143),
.B(n_1129),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1149),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1146),
.B(n_1141),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1144),
.A2(n_1141),
.B1(n_1128),
.B2(n_1134),
.C(n_1132),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1145),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1150),
.A2(n_1142),
.B(n_951),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1147),
.B(n_1142),
.Y(n_1158)
);

NAND4xp25_ASAP7_75t_SL g1159 ( 
.A(n_1156),
.B(n_1139),
.C(n_981),
.D(n_961),
.Y(n_1159)
);

OAI211xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1153),
.A2(n_1132),
.B(n_1131),
.C(n_981),
.Y(n_1160)
);

NOR3xp33_ASAP7_75t_L g1161 ( 
.A(n_1157),
.B(n_968),
.C(n_949),
.Y(n_1161)
);

NOR3x1_ASAP7_75t_L g1162 ( 
.A(n_1154),
.B(n_1026),
.C(n_1052),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1152),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_1151),
.B(n_1044),
.Y(n_1164)
);

AOI211xp5_ASAP7_75t_L g1165 ( 
.A1(n_1159),
.A2(n_1155),
.B(n_1158),
.C(n_1044),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1163),
.B(n_1131),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1161),
.A2(n_1139),
.B1(n_1081),
.B2(n_1041),
.Y(n_1167)
);

NOR4xp25_ASAP7_75t_L g1168 ( 
.A(n_1160),
.B(n_1002),
.C(n_988),
.D(n_1042),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1164),
.A2(n_1041),
.B1(n_1046),
.B2(n_1044),
.Y(n_1169)
);

NOR2x1p5_ASAP7_75t_SL g1170 ( 
.A(n_1162),
.B(n_1055),
.Y(n_1170)
);

NOR2x1_ASAP7_75t_L g1171 ( 
.A(n_1166),
.B(n_958),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1167),
.B(n_1105),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_L g1173 ( 
.A(n_1170),
.B(n_974),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1165),
.B(n_971),
.C(n_999),
.Y(n_1174)
);

NOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1168),
.B(n_974),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1172),
.B(n_1169),
.Y(n_1176)
);

XNOR2x1_ASAP7_75t_L g1177 ( 
.A(n_1175),
.B(n_1013),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1176),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1178),
.Y(n_1179)
);

AOI22x1_ASAP7_75t_L g1180 ( 
.A1(n_1179),
.A2(n_1174),
.B1(n_1177),
.B2(n_1171),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1180),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1181),
.A2(n_1173),
.B1(n_971),
.B2(n_989),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1182),
.A2(n_989),
.B1(n_1053),
.B2(n_972),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1183),
.B(n_983),
.Y(n_1184)
);

BUFx24_ASAP7_75t_SL g1185 ( 
.A(n_1184),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1185),
.A2(n_1051),
.B(n_983),
.Y(n_1186)
);


endmodule