module real_aes_11629_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_1369;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_0), .A2(n_20), .B1(n_529), .B2(n_539), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_0), .A2(n_232), .B1(n_365), .B2(n_542), .Y(n_609) );
INVx1_ASAP7_75t_L g928 ( .A(n_1), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_1), .A2(n_136), .B1(n_794), .B2(n_801), .Y(n_938) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_2), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_2), .A2(n_25), .B1(n_390), .B2(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g706 ( .A(n_3), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_4), .A2(n_167), .B1(n_542), .B2(n_552), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_4), .A2(n_167), .B1(n_524), .B2(n_807), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_5), .A2(n_12), .B1(n_514), .B2(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g953 ( .A(n_5), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_6), .A2(n_111), .B1(n_390), .B2(n_798), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_6), .A2(n_111), .B1(n_524), .B2(n_674), .Y(n_991) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_7), .Y(n_262) );
INVx1_ASAP7_75t_L g397 ( .A(n_7), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_7), .B(n_188), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_7), .B(n_344), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_8), .A2(n_57), .B1(n_1017), .B2(n_1021), .Y(n_1016) );
INVx1_ASAP7_75t_L g1234 ( .A(n_9), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_9), .A2(n_177), .B1(n_1281), .B2(n_1285), .Y(n_1280) );
AOI22xp33_ASAP7_75t_SL g1260 ( .A1(n_10), .A2(n_49), .B1(n_1257), .B2(n_1261), .Y(n_1260) );
INVx1_ASAP7_75t_L g1315 ( .A(n_10), .Y(n_1315) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_11), .A2(n_202), .B1(n_376), .B2(n_377), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_11), .A2(n_202), .B1(n_406), .B2(n_417), .Y(n_463) );
INVx1_ASAP7_75t_L g954 ( .A(n_12), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_13), .A2(n_91), .B1(n_604), .B2(n_677), .Y(n_1354) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_13), .A2(n_91), .B1(n_650), .B2(n_1369), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_14), .A2(n_171), .B1(n_376), .B2(n_377), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_14), .A2(n_171), .B1(n_404), .B2(n_406), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_15), .A2(n_198), .B1(n_793), .B2(n_794), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_15), .A2(n_198), .B1(n_413), .B2(n_805), .Y(n_804) );
AO22x2_ASAP7_75t_L g692 ( .A1(n_16), .A2(n_693), .B1(n_761), .B2(n_762), .Y(n_692) );
INVx1_ASAP7_75t_L g761 ( .A(n_16), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_17), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_18), .A2(n_131), .B1(n_440), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_18), .A2(n_131), .B1(n_604), .B2(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g293 ( .A(n_19), .Y(n_293) );
INVx1_ASAP7_75t_L g594 ( .A(n_20), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_21), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_22), .A2(n_65), .B1(n_1021), .B2(n_1035), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_23), .A2(n_241), .B1(n_731), .B2(n_732), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_23), .A2(n_241), .B1(n_744), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g926 ( .A(n_24), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_24), .A2(n_247), .B1(n_390), .B2(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g315 ( .A(n_25), .Y(n_315) );
INVx1_ASAP7_75t_L g427 ( .A(n_26), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_26), .A2(n_127), .B1(n_336), .B2(n_454), .Y(n_458) );
XNOR2xp5_ASAP7_75t_L g557 ( .A(n_27), .B(n_558), .Y(n_557) );
INVxp67_ASAP7_75t_SL g643 ( .A(n_28), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_28), .A2(n_194), .B1(n_686), .B2(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g277 ( .A(n_29), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g1033 ( .A1(n_29), .A2(n_128), .B1(n_1005), .B2(n_1013), .Y(n_1033) );
INVx2_ASAP7_75t_L g285 ( .A(n_30), .Y(n_285) );
OR2x2_ASAP7_75t_L g1278 ( .A(n_30), .B(n_1272), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_31), .A2(n_214), .B1(n_376), .B2(n_820), .Y(n_819) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_31), .Y(n_850) );
INVx1_ASAP7_75t_L g1339 ( .A(n_32), .Y(n_1339) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_32), .A2(n_115), .B1(n_673), .B2(n_1353), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_33), .A2(n_181), .B1(n_705), .B2(n_833), .Y(n_832) );
OAI211xp5_ASAP7_75t_SL g836 ( .A1(n_33), .A2(n_546), .B(n_837), .C(n_840), .Y(n_836) );
BUFx2_ASAP7_75t_L g331 ( .A(n_34), .Y(n_331) );
BUFx2_ASAP7_75t_L g372 ( .A(n_34), .Y(n_372) );
INVx1_ASAP7_75t_L g668 ( .A(n_34), .Y(n_668) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_34), .B(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g878 ( .A(n_35), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_35), .A2(n_207), .B1(n_336), .B2(n_801), .Y(n_893) );
INVx1_ASAP7_75t_L g1058 ( .A(n_36), .Y(n_1058) );
INVx1_ASAP7_75t_L g1332 ( .A(n_37), .Y(n_1332) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_37), .A2(n_96), .B1(n_727), .B2(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1346 ( .A(n_38), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_38), .A2(n_44), .B1(n_677), .B2(n_1351), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_39), .A2(n_170), .B1(n_454), .B2(n_794), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_39), .A2(n_170), .B1(n_301), .B2(n_825), .Y(n_824) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_40), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_40), .A2(n_123), .B1(n_349), .B2(n_641), .Y(n_640) );
INVxp33_ASAP7_75t_L g976 ( .A(n_41), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_41), .A2(n_149), .B1(n_789), .B2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g607 ( .A(n_42), .Y(n_607) );
INVx1_ASAP7_75t_L g1096 ( .A(n_43), .Y(n_1096) );
INVx1_ASAP7_75t_L g1341 ( .A(n_44), .Y(n_1341) );
INVx1_ASAP7_75t_L g431 ( .A(n_45), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_45), .A2(n_229), .B1(n_377), .B2(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g281 ( .A(n_46), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_46), .A2(n_187), .B1(n_336), .B2(n_379), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_47), .A2(n_240), .B1(n_406), .B2(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_47), .A2(n_172), .B1(n_365), .B2(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g699 ( .A(n_48), .Y(n_699) );
INVx1_ASAP7_75t_L g1279 ( .A(n_49), .Y(n_1279) );
XNOR2xp5_ASAP7_75t_L g765 ( .A(n_50), .B(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_50), .A2(n_104), .B1(n_1005), .B2(n_1013), .Y(n_1038) );
INVx1_ASAP7_75t_L g1331 ( .A(n_51), .Y(n_1331) );
AOI22xp33_ASAP7_75t_SL g1360 ( .A1(n_51), .A2(n_69), .B1(n_1361), .B2(n_1363), .Y(n_1360) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_52), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_53), .A2(n_211), .B1(n_793), .B2(n_794), .Y(n_821) );
INVx1_ASAP7_75t_L g847 ( .A(n_53), .Y(n_847) );
INVxp33_ASAP7_75t_L g968 ( .A(n_54), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_54), .A2(n_89), .B1(n_746), .B2(n_825), .Y(n_993) );
INVx1_ASAP7_75t_L g497 ( .A(n_55), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_55), .A2(n_172), .B1(n_527), .B2(n_529), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_56), .A2(n_178), .B1(n_263), .B2(n_365), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_56), .A2(n_174), .B1(n_461), .B2(n_805), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_58), .A2(n_235), .B1(n_301), .B2(n_461), .Y(n_943) );
INVx1_ASAP7_75t_L g949 ( .A(n_58), .Y(n_949) );
INVx1_ASAP7_75t_L g606 ( .A(n_59), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g1062 ( .A1(n_60), .A2(n_114), .B1(n_1005), .B2(n_1013), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_61), .A2(n_205), .B1(n_659), .B2(n_801), .Y(n_1262) );
INVx1_ASAP7_75t_L g1298 ( .A(n_61), .Y(n_1298) );
INVx1_ASAP7_75t_L g775 ( .A(n_62), .Y(n_775) );
INVx1_ASAP7_75t_L g573 ( .A(n_63), .Y(n_573) );
INVx1_ASAP7_75t_L g778 ( .A(n_64), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_64), .A2(n_125), .B1(n_390), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1251 ( .A(n_66), .Y(n_1251) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_66), .A2(n_110), .B1(n_831), .B2(n_1289), .C(n_1290), .Y(n_1288) );
INVx1_ASAP7_75t_L g965 ( .A(n_67), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_68), .A2(n_245), .B1(n_376), .B2(n_377), .Y(n_888) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_68), .A2(n_245), .B1(n_514), .B2(n_827), .Y(n_896) );
OAI222xp33_ASAP7_75t_L g1327 ( .A1(n_69), .A2(n_155), .B1(n_236), .B2(n_306), .C1(n_311), .C2(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g449 ( .A(n_70), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g466 ( .A1(n_70), .A2(n_81), .B1(n_417), .B2(n_418), .Y(n_466) );
INVx1_ASAP7_75t_L g491 ( .A(n_71), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_71), .A2(n_161), .B1(n_538), .B2(n_539), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_72), .A2(n_147), .B1(n_336), .B2(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_72), .A2(n_147), .B1(n_301), .B2(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_73), .A2(n_102), .B1(n_311), .B2(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_73), .A2(n_102), .B1(n_349), .B2(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g362 ( .A(n_74), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_74), .A2(n_94), .B1(n_417), .B2(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g578 ( .A(n_75), .Y(n_578) );
OAI211xp5_ASAP7_75t_SL g610 ( .A1(n_75), .A2(n_544), .B(n_546), .C(n_611), .Y(n_610) );
AO22x2_ASAP7_75t_L g957 ( .A1(n_76), .A2(n_958), .B1(n_995), .B2(n_996), .Y(n_957) );
INVx1_ASAP7_75t_L g995 ( .A(n_76), .Y(n_995) );
CKINVDCx5p33_ASAP7_75t_R g1249 ( .A(n_77), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1321 ( .A1(n_78), .A2(n_1322), .B1(n_1371), .B2(n_1372), .Y(n_1321) );
CKINVDCx5p33_ASAP7_75t_R g1372 ( .A(n_78), .Y(n_1372) );
INVxp67_ASAP7_75t_SL g700 ( .A(n_79), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g736 ( .A1(n_79), .A2(n_193), .B1(n_727), .B2(n_737), .Y(n_736) );
AO22x2_ASAP7_75t_L g861 ( .A1(n_80), .A2(n_862), .B1(n_901), .B2(n_902), .Y(n_861) );
INVxp67_ASAP7_75t_L g901 ( .A(n_80), .Y(n_901) );
INVx1_ASAP7_75t_L g447 ( .A(n_81), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_82), .Y(n_1055) );
INVx1_ASAP7_75t_L g853 ( .A(n_83), .Y(n_853) );
INVx1_ASAP7_75t_L g329 ( .A(n_84), .Y(n_329) );
INVx1_ASAP7_75t_L g1272 ( .A(n_84), .Y(n_1272) );
INVxp33_ASAP7_75t_SL g713 ( .A(n_85), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_85), .A2(n_186), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g702 ( .A(n_86), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_86), .A2(n_176), .B1(n_732), .B2(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g842 ( .A(n_87), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_88), .A2(n_192), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_88), .A2(n_192), .B1(n_748), .B2(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g964 ( .A(n_89), .Y(n_964) );
INVx1_ASAP7_75t_L g522 ( .A(n_90), .Y(n_522) );
OAI211xp5_ASAP7_75t_SL g543 ( .A1(n_90), .A2(n_544), .B(n_546), .C(n_547), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_92), .A2(n_183), .B1(n_306), .B2(n_311), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_92), .A2(n_183), .B1(n_346), .B2(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g567 ( .A(n_93), .Y(n_567) );
INVxp67_ASAP7_75t_L g370 ( .A(n_94), .Y(n_370) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_95), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_95), .A2(n_233), .B1(n_662), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g1335 ( .A(n_96), .Y(n_1335) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_97), .A2(n_117), .B1(n_1005), .B2(n_1013), .Y(n_1004) );
INVx1_ASAP7_75t_L g598 ( .A(n_98), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_99), .A2(n_138), .B1(n_514), .B2(n_831), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_99), .A2(n_138), .B1(n_542), .B2(n_552), .Y(n_835) );
INVx1_ASAP7_75t_L g930 ( .A(n_100), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g950 ( .A1(n_100), .A2(n_175), .B1(n_641), .B2(n_951), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_101), .A2(n_201), .B1(n_1005), .B2(n_1013), .Y(n_1042) );
INVx1_ASAP7_75t_L g865 ( .A(n_103), .Y(n_865) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_103), .A2(n_215), .B1(n_417), .B2(n_418), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_105), .A2(n_130), .B1(n_1021), .B2(n_1035), .Y(n_1039) );
INVx1_ASAP7_75t_L g1026 ( .A(n_106), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_107), .A2(n_134), .B1(n_758), .B2(n_1353), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_107), .A2(n_134), .B1(n_654), .B2(n_1365), .Y(n_1364) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_108), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_108), .A2(n_182), .B1(n_406), .B2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_109), .A2(n_200), .B1(n_383), .B2(n_793), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_109), .A2(n_200), .B1(n_413), .B2(n_414), .Y(n_895) );
INVx1_ASAP7_75t_L g1241 ( .A(n_110), .Y(n_1241) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_112), .A2(n_222), .B1(n_376), .B2(n_377), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_112), .A2(n_222), .B1(n_686), .B2(n_831), .Y(n_941) );
INVx1_ASAP7_75t_L g577 ( .A(n_113), .Y(n_577) );
OAI22xp33_ASAP7_75t_SL g612 ( .A1(n_113), .A2(n_145), .B1(n_263), .B2(n_552), .Y(n_612) );
INVx1_ASAP7_75t_L g1338 ( .A(n_115), .Y(n_1338) );
INVx1_ASAP7_75t_L g254 ( .A(n_116), .Y(n_254) );
INVx1_ASAP7_75t_L g446 ( .A(n_118), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_118), .A2(n_197), .B1(n_414), .B2(n_461), .Y(n_465) );
AO22x1_ASAP7_75t_SL g1023 ( .A1(n_119), .A2(n_208), .B1(n_1005), .B2(n_1013), .Y(n_1023) );
INVx1_ASAP7_75t_L g1094 ( .A(n_120), .Y(n_1094) );
AO221x2_ASAP7_75t_L g1052 ( .A1(n_121), .A2(n_237), .B1(n_1017), .B2(n_1053), .C(n_1054), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_122), .A2(n_181), .B1(n_263), .B2(n_365), .Y(n_843) );
OAI22xp33_ASAP7_75t_L g852 ( .A1(n_122), .A2(n_211), .B1(n_527), .B2(n_529), .Y(n_852) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_123), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_124), .Y(n_874) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_125), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_126), .A2(n_146), .B1(n_1257), .B2(n_1258), .Y(n_1256) );
AOI221xp5_ASAP7_75t_L g1299 ( .A1(n_126), .A2(n_239), .B1(n_404), .B2(n_1300), .C(n_1301), .Y(n_1299) );
INVx1_ASAP7_75t_L g434 ( .A(n_127), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_129), .A2(n_154), .B1(n_654), .B2(n_656), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_129), .A2(n_154), .B1(n_673), .B2(n_674), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_132), .A2(n_239), .B1(n_383), .B2(n_801), .Y(n_1255) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_132), .A2(n_146), .B1(n_1303), .B2(n_1304), .Y(n_1302) );
XOR2xp5_ASAP7_75t_L g468 ( .A(n_133), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g969 ( .A(n_135), .Y(n_969) );
INVx1_ASAP7_75t_L g925 ( .A(n_136), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_137), .A2(n_143), .B1(n_376), .B2(n_816), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_137), .A2(n_143), .B1(n_524), .B2(n_827), .Y(n_826) );
OAI22xp33_ASAP7_75t_L g779 ( .A1(n_139), .A2(n_178), .B1(n_527), .B2(n_529), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_139), .A2(n_210), .B1(n_801), .B2(n_802), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_140), .A2(n_231), .B1(n_1021), .B2(n_1035), .Y(n_1043) );
INVxp33_ASAP7_75t_L g962 ( .A(n_141), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_141), .A2(n_148), .B1(n_524), .B2(n_831), .Y(n_994) );
INVx1_ASAP7_75t_L g570 ( .A(n_142), .Y(n_570) );
INVx1_ASAP7_75t_L g966 ( .A(n_144), .Y(n_966) );
INVx1_ASAP7_75t_L g582 ( .A(n_145), .Y(n_582) );
INVxp33_ASAP7_75t_L g961 ( .A(n_148), .Y(n_961) );
INVxp33_ASAP7_75t_L g978 ( .A(n_149), .Y(n_978) );
INVx1_ASAP7_75t_L g593 ( .A(n_150), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g600 ( .A1(n_150), .A2(n_166), .B1(n_527), .B2(n_538), .Y(n_600) );
INVx1_ASAP7_75t_L g480 ( .A(n_151), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_152), .A2(n_227), .B1(n_660), .B2(n_793), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_152), .A2(n_227), .B1(n_301), .B2(n_461), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_153), .A2(n_213), .B1(n_379), .B2(n_794), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_153), .A2(n_213), .B1(n_301), .B2(n_899), .Y(n_990) );
INVx1_ASAP7_75t_L g1343 ( .A(n_155), .Y(n_1343) );
INVx1_ASAP7_75t_L g1273 ( .A(n_156), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_157), .A2(n_223), .B1(n_1017), .B2(n_1021), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_158), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_158), .B(n_254), .Y(n_1012) );
AND3x2_ASAP7_75t_L g1020 ( .A(n_158), .B(n_254), .C(n_1009), .Y(n_1020) );
INVxp33_ASAP7_75t_SL g632 ( .A(n_159), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_159), .A2(n_224), .B1(n_650), .B2(n_659), .Y(n_658) );
INVxp33_ASAP7_75t_L g979 ( .A(n_160), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_160), .A2(n_164), .B1(n_793), .B2(n_794), .Y(n_988) );
INVx1_ASAP7_75t_L g494 ( .A(n_161), .Y(n_494) );
INVx1_ASAP7_75t_L g773 ( .A(n_162), .Y(n_773) );
INVx2_ASAP7_75t_L g267 ( .A(n_163), .Y(n_267) );
INVx1_ASAP7_75t_L g974 ( .A(n_164), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_165), .Y(n_1246) );
INVx1_ASAP7_75t_L g596 ( .A(n_166), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_168), .A2(n_196), .B1(n_789), .B2(n_790), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_168), .A2(n_196), .B1(n_524), .B2(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g1028 ( .A(n_169), .Y(n_1028) );
INVx1_ASAP7_75t_L g1009 ( .A(n_173), .Y(n_1009) );
OAI211xp5_ASAP7_75t_L g782 ( .A1(n_174), .A2(n_544), .B(n_546), .C(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g929 ( .A(n_175), .Y(n_929) );
INVxp33_ASAP7_75t_SL g696 ( .A(n_176), .Y(n_696) );
INVx1_ASAP7_75t_L g1237 ( .A(n_177), .Y(n_1237) );
INVx1_ASAP7_75t_L g884 ( .A(n_179), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_179), .A2(n_221), .B1(n_390), .B2(n_892), .Y(n_891) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_180), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_180), .A2(n_217), .B1(n_680), .B2(n_683), .Y(n_679) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_182), .Y(n_482) );
INVx1_ASAP7_75t_L g476 ( .A(n_184), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_185), .Y(n_429) );
INVxp33_ASAP7_75t_SL g714 ( .A(n_186), .Y(n_714) );
INVx1_ASAP7_75t_L g304 ( .A(n_187), .Y(n_304) );
INVx1_ASAP7_75t_L g269 ( .A(n_188), .Y(n_269) );
INVx2_ASAP7_75t_L g344 ( .A(n_188), .Y(n_344) );
INVx1_ASAP7_75t_L g334 ( .A(n_189), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_189), .A2(n_238), .B1(n_413), .B2(n_414), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_190), .A2(n_219), .B1(n_379), .B2(n_383), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_190), .A2(n_219), .B1(n_400), .B2(n_401), .Y(n_399) );
XNOR2xp5_ASAP7_75t_L g423 ( .A(n_191), .B(n_424), .Y(n_423) );
INVxp33_ASAP7_75t_SL g697 ( .A(n_193), .Y(n_697) );
INVxp33_ASAP7_75t_SL g644 ( .A(n_194), .Y(n_644) );
AO22x2_ASAP7_75t_L g619 ( .A1(n_195), .A2(n_620), .B1(n_689), .B2(n_690), .Y(n_619) );
CKINVDCx14_ASAP7_75t_R g689 ( .A(n_195), .Y(n_689) );
INVx1_ASAP7_75t_L g439 ( .A(n_197), .Y(n_439) );
INVx1_ASAP7_75t_L g868 ( .A(n_199), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_199), .A2(n_244), .B1(n_401), .B2(n_899), .Y(n_898) );
OAI211xp5_ASAP7_75t_L g905 ( .A1(n_199), .A2(n_546), .B(n_906), .C(n_908), .Y(n_905) );
XNOR2xp5_ASAP7_75t_L g918 ( .A(n_201), .B(n_919), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g1090 ( .A1(n_203), .A2(n_204), .B1(n_1091), .B2(n_1092), .C(n_1093), .Y(n_1090) );
AOI222xp33_ASAP7_75t_L g1222 ( .A1(n_203), .A2(n_1223), .B1(n_1319), .B2(n_1321), .C1(n_1373), .C2(n_1377), .Y(n_1222) );
XOR2x1_ASAP7_75t_L g1224 ( .A(n_203), .B(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1312 ( .A(n_205), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g1334 ( .A(n_206), .Y(n_1334) );
INVx1_ASAP7_75t_L g882 ( .A(n_207), .Y(n_882) );
OAI211xp5_ASAP7_75t_L g912 ( .A1(n_207), .A2(n_536), .B(n_913), .C(n_915), .Y(n_912) );
INVx1_ASAP7_75t_L g519 ( .A(n_209), .Y(n_519) );
OAI22xp33_ASAP7_75t_SL g551 ( .A1(n_209), .A2(n_240), .B1(n_263), .B2(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g770 ( .A(n_210), .Y(n_770) );
INVx1_ASAP7_75t_L g629 ( .A(n_212), .Y(n_629) );
INVx1_ASAP7_75t_L g851 ( .A(n_214), .Y(n_851) );
INVx1_ASAP7_75t_L g866 ( .A(n_215), .Y(n_866) );
INVx1_ASAP7_75t_L g1010 ( .A(n_216), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_216), .B(n_1008), .Y(n_1015) );
INVxp33_ASAP7_75t_SL g637 ( .A(n_217), .Y(n_637) );
INVx1_ASAP7_75t_L g564 ( .A(n_218), .Y(n_564) );
INVx1_ASAP7_75t_L g708 ( .A(n_220), .Y(n_708) );
INVx1_ASAP7_75t_L g879 ( .A(n_221), .Y(n_879) );
INVx1_ASAP7_75t_L g623 ( .A(n_224), .Y(n_623) );
INVx1_ASAP7_75t_L g841 ( .A(n_225), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_226), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_228), .Y(n_534) );
INVx1_ASAP7_75t_L g432 ( .A(n_229), .Y(n_432) );
INVx2_ASAP7_75t_L g266 ( .A(n_230), .Y(n_266) );
INVx1_ASAP7_75t_L g584 ( .A(n_232), .Y(n_584) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_233), .Y(n_633) );
INVxp33_ASAP7_75t_SL g723 ( .A(n_234), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_234), .A2(n_248), .B1(n_754), .B2(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g956 ( .A(n_235), .Y(n_956) );
INVx1_ASAP7_75t_L g1344 ( .A(n_236), .Y(n_1344) );
INVxp33_ASAP7_75t_L g354 ( .A(n_238), .Y(n_354) );
BUFx3_ASAP7_75t_L g290 ( .A(n_242), .Y(n_290) );
INVx1_ASAP7_75t_L g323 ( .A(n_242), .Y(n_323) );
BUFx3_ASAP7_75t_L g292 ( .A(n_243), .Y(n_292) );
INVx1_ASAP7_75t_L g318 ( .A(n_243), .Y(n_318) );
INVx1_ASAP7_75t_L g873 ( .A(n_244), .Y(n_873) );
INVx1_ASAP7_75t_L g500 ( .A(n_246), .Y(n_500) );
INVx1_ASAP7_75t_L g923 ( .A(n_247), .Y(n_923) );
INVx1_ASAP7_75t_L g718 ( .A(n_248), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_998), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_257), .Y(n_251) );
AND2x4_ASAP7_75t_L g1320 ( .A(n_252), .B(n_258), .Y(n_1320) );
NOR2xp33_ASAP7_75t_SL g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_SL g1376 ( .A(n_253), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_253), .B(n_255), .Y(n_1382) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_255), .B(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_263), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g371 ( .A(n_260), .B(n_372), .Y(n_371) );
OR2x6_ASAP7_75t_L g556 ( .A(n_260), .B(n_372), .Y(n_556) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g387 ( .A(n_261), .B(n_269), .Y(n_387) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g473 ( .A(n_262), .B(n_357), .Y(n_473) );
INVx8_ASAP7_75t_L g353 ( .A(n_263), .Y(n_353) );
OR2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
OR2x6_ASAP7_75t_L g365 ( .A(n_264), .B(n_356), .Y(n_365) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_264), .Y(n_475) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_264), .Y(n_496) );
INVx2_ASAP7_75t_SL g589 ( .A(n_264), .Y(n_589) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_264), .B(n_1232), .Y(n_1266) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g338 ( .A(n_266), .Y(n_338) );
INVx1_ASAP7_75t_L g351 ( .A(n_266), .Y(n_351) );
INVx2_ASAP7_75t_L g359 ( .A(n_266), .Y(n_359) );
AND2x4_ASAP7_75t_L g369 ( .A(n_266), .B(n_339), .Y(n_369) );
AND2x2_ASAP7_75t_L g382 ( .A(n_266), .B(n_267), .Y(n_382) );
INVx2_ASAP7_75t_L g339 ( .A(n_267), .Y(n_339) );
INVx1_ASAP7_75t_L g348 ( .A(n_267), .Y(n_348) );
INVx1_ASAP7_75t_L g361 ( .A(n_267), .Y(n_361) );
INVx1_ASAP7_75t_L g479 ( .A(n_267), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_267), .B(n_359), .Y(n_485) );
AND2x4_ASAP7_75t_L g347 ( .A(n_268), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g349 ( .A(n_269), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g951 ( .A(n_269), .B(n_350), .Y(n_951) );
XNOR2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_615), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
XOR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_467), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B1(n_422), .B2(n_423), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
XNOR2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AOI211xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_327), .B(n_332), .C(n_373), .Y(n_278) );
NAND4xp25_ASAP7_75t_L g279 ( .A(n_280), .B(n_297), .C(n_314), .D(n_324), .Y(n_279) );
AOI22xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_282), .B1(n_293), .B2(n_294), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_282), .A2(n_316), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_282), .A2(n_316), .B1(n_696), .B2(n_697), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_282), .A2(n_316), .B1(n_925), .B2(n_926), .Y(n_924) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
AND2x6_ASAP7_75t_L g320 ( .A(n_283), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g428 ( .A(n_283), .B(n_286), .Y(n_428) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g307 ( .A(n_284), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_285), .Y(n_296) );
INVx1_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
AND2x2_ASAP7_75t_L g410 ( .A(n_285), .B(n_329), .Y(n_410) );
INVx2_ASAP7_75t_L g421 ( .A(n_285), .Y(n_421) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g400 ( .A(n_287), .Y(n_400) );
INVx2_ASAP7_75t_L g678 ( .A(n_287), .Y(n_678) );
INVx2_ASAP7_75t_SL g682 ( .A(n_287), .Y(n_682) );
BUFx6f_ASAP7_75t_L g745 ( .A(n_287), .Y(n_745) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_287), .Y(n_755) );
INVx1_ASAP7_75t_L g833 ( .A(n_287), .Y(n_833) );
INVx6_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g294 ( .A(n_288), .B(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g413 ( .A(n_288), .Y(n_413) );
INVx2_ASAP7_75t_L g462 ( .A(n_288), .Y(n_462) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_288), .B(n_1270), .Y(n_1269) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_290), .B(n_292), .Y(n_303) );
AND2x4_ASAP7_75t_L g317 ( .A(n_290), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g310 ( .A(n_291), .Y(n_310) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_L g322 ( .A(n_292), .B(n_323), .Y(n_322) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_293), .A2(n_364), .B1(n_366), .B2(n_370), .Y(n_363) );
AOI22xp5_ASAP7_75t_SL g426 ( .A1(n_294), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_426) );
INVx4_ASAP7_75t_L g529 ( .A(n_294), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_294), .A2(n_320), .B1(n_629), .B2(n_630), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_294), .A2(n_320), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_294), .A2(n_320), .B1(n_874), .B2(n_884), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_294), .A2(n_320), .B1(n_922), .B2(n_923), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g975 ( .A1(n_294), .A2(n_320), .B1(n_325), .B2(n_969), .C(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_294), .A2(n_320), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
AND2x4_ASAP7_75t_L g625 ( .A(n_295), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_SL g774 ( .A(n_295), .B(n_626), .Y(n_774) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B(n_305), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_298), .A2(n_434), .B(n_435), .Y(n_433) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x6_ASAP7_75t_L g316 ( .A(n_299), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g326 ( .A(n_299), .Y(n_326) );
INVx1_ASAP7_75t_L g528 ( .A(n_299), .Y(n_528) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x6_ASAP7_75t_L g312 ( .A(n_300), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_301), .Y(n_881) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g325 ( .A(n_302), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g402 ( .A(n_302), .Y(n_402) );
INVx2_ASAP7_75t_L g605 ( .A(n_302), .Y(n_605) );
BUFx6f_ASAP7_75t_L g973 ( .A(n_302), .Y(n_973) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_303), .Y(n_415) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g436 ( .A(n_307), .Y(n_436) );
AOI222xp33_ASAP7_75t_L g531 ( .A1(n_307), .A2(n_312), .B1(n_500), .B2(n_532), .C1(n_534), .C2(n_535), .Y(n_531) );
AOI222xp33_ASAP7_75t_L g603 ( .A1(n_307), .A2(n_312), .B1(n_598), .B2(n_604), .C1(n_606), .C2(n_607), .Y(n_603) );
AOI222xp33_ASAP7_75t_L g846 ( .A1(n_307), .A2(n_312), .B1(n_841), .B2(n_842), .C1(n_847), .C2(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g626 ( .A(n_309), .Y(n_626) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g1284 ( .A(n_310), .Y(n_1284) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI222xp33_ASAP7_75t_L g622 ( .A1(n_312), .A2(n_401), .B1(n_623), .B2(n_624), .C1(n_625), .C2(n_627), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g701 ( .A1(n_312), .A2(n_702), .B1(n_703), .B2(n_706), .C1(n_707), .C2(n_708), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g769 ( .A1(n_312), .A2(n_770), .B1(n_771), .B2(n_773), .C1(n_774), .C2(n_775), .Y(n_769) );
AOI222xp33_ASAP7_75t_L g880 ( .A1(n_312), .A2(n_707), .B1(n_869), .B2(n_870), .C1(n_881), .C2(n_882), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g915 ( .A1(n_312), .A2(n_625), .B1(n_869), .B2(n_870), .Y(n_915) );
AOI222xp33_ASAP7_75t_L g927 ( .A1(n_312), .A2(n_756), .B1(n_774), .B2(n_928), .C1(n_929), .C2(n_930), .Y(n_927) );
AOI222xp33_ASAP7_75t_L g971 ( .A1(n_312), .A2(n_774), .B1(n_965), .B2(n_966), .C1(n_972), .C2(n_974), .Y(n_971) );
BUFx3_ASAP7_75t_L g1287 ( .A(n_313), .Y(n_1287) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_319), .B2(n_320), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_316), .A2(n_320), .B1(n_431), .B2(n_432), .Y(n_430) );
CKINVDCx6p67_ASAP7_75t_R g538 ( .A(n_316), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_316), .A2(n_320), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_316), .A2(n_320), .B1(n_850), .B2(n_851), .Y(n_849) );
AOI22xp5_ASAP7_75t_SL g877 ( .A1(n_316), .A2(n_428), .B1(n_878), .B2(n_879), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_316), .A2(n_428), .B1(n_978), .B2(n_979), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_316), .A2(n_428), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
INVx2_ASAP7_75t_SL g405 ( .A(n_317), .Y(n_405) );
BUFx3_ASAP7_75t_L g417 ( .A(n_317), .Y(n_417) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_317), .Y(n_514) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_317), .Y(n_524) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_317), .Y(n_566) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_317), .Y(n_581) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_317), .Y(n_758) );
INVx1_ASAP7_75t_L g508 ( .A(n_318), .Y(n_508) );
INVx4_ASAP7_75t_L g539 ( .A(n_320), .Y(n_539) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_321), .Y(n_418) );
INVx2_ASAP7_75t_L g583 ( .A(n_321), .Y(n_583) );
INVx1_ASAP7_75t_L g675 ( .A(n_321), .Y(n_675) );
INVx1_ASAP7_75t_L g688 ( .A(n_321), .Y(n_688) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_321), .Y(n_831) );
INVx1_ASAP7_75t_L g946 ( .A(n_321), .Y(n_946) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_322), .Y(n_406) );
INVx1_ASAP7_75t_L g828 ( .A(n_322), .Y(n_828) );
INVx2_ASAP7_75t_L g1307 ( .A(n_322), .Y(n_1307) );
INVx1_ASAP7_75t_L g507 ( .A(n_323), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_324), .B(n_426), .C(n_430), .D(n_433), .Y(n_425) );
BUFx2_ASAP7_75t_L g709 ( .A(n_324), .Y(n_709) );
NAND4xp25_ASAP7_75t_L g876 ( .A(n_324), .B(n_877), .C(n_880), .D(n_883), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g920 ( .A(n_324), .B(n_921), .C(n_924), .D(n_927), .Y(n_920) );
INVx5_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
CKINVDCx8_ASAP7_75t_R g536 ( .A(n_325), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g1326 ( .A(n_325), .B(n_1327), .Y(n_1326) );
AOI211xp5_ASAP7_75t_L g424 ( .A1(n_327), .A2(n_425), .B(n_437), .C(n_450), .Y(n_424) );
OAI31xp33_ASAP7_75t_SL g525 ( .A1(n_327), .A2(n_526), .A3(n_530), .B(n_537), .Y(n_525) );
OAI31xp33_ASAP7_75t_L g599 ( .A1(n_327), .A2(n_600), .A3(n_601), .B(n_602), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_327), .A2(n_768), .B(n_779), .Y(n_767) );
OAI21xp5_ASAP7_75t_SL g844 ( .A1(n_327), .A2(n_845), .B(n_852), .Y(n_844) );
AOI211xp5_ASAP7_75t_L g919 ( .A1(n_327), .A2(n_920), .B(n_931), .C(n_947), .Y(n_919) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
AND2x4_ASAP7_75t_L g634 ( .A(n_328), .B(n_330), .Y(n_634) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g420 ( .A(n_329), .B(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g386 ( .A(n_331), .Y(n_386) );
OR2x6_ASAP7_75t_L g472 ( .A(n_331), .B(n_473), .Y(n_472) );
AOI31xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_352), .A3(n_363), .B(n_371), .Y(n_332) );
AOI211xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_335), .B(n_340), .C(n_345), .Y(n_333) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x6_ASAP7_75t_L g1247 ( .A(n_336), .B(n_1244), .Y(n_1247) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g340 ( .A(n_337), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_337), .Y(n_442) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_337), .Y(n_660) );
BUFx2_ASAP7_75t_L g721 ( .A(n_337), .Y(n_721) );
BUFx3_ASAP7_75t_L g795 ( .A(n_337), .Y(n_795) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g438 ( .A1(n_340), .A2(n_439), .B(n_440), .C(n_443), .Y(n_438) );
CKINVDCx11_ASAP7_75t_R g546 ( .A(n_340), .Y(n_546) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_340), .A2(n_383), .B(n_639), .C(n_640), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g948 ( .A1(n_340), .A2(n_659), .B(n_949), .C(n_950), .Y(n_948) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g550 ( .A(n_342), .Y(n_550) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_343), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g357 ( .A(n_344), .Y(n_357) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g444 ( .A(n_347), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_347), .A2(n_534), .B1(n_535), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_347), .A2(n_548), .B1(n_606), .B2(n_607), .Y(n_611) );
INVx2_ASAP7_75t_L g641 ( .A(n_347), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_347), .A2(n_548), .B1(n_841), .B2(n_842), .Y(n_840) );
HB1xp67_ASAP7_75t_L g1236 ( .A(n_348), .Y(n_1236) );
INVx1_ASAP7_75t_L g549 ( .A(n_350), .Y(n_549) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_351), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g499 ( .A(n_351), .B(n_479), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_354), .B1(n_355), .B2(n_362), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_353), .A2(n_355), .B1(n_446), .B2(n_447), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_353), .A2(n_364), .B1(n_629), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_353), .A2(n_364), .B1(n_699), .B2(n_723), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_353), .A2(n_873), .B1(n_874), .B2(n_875), .Y(n_872) );
AOI22xp33_ASAP7_75t_SL g955 ( .A1(n_353), .A2(n_875), .B1(n_922), .B2(n_956), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_353), .A2(n_364), .B1(n_968), .B2(n_969), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_353), .A2(n_875), .B1(n_1334), .B2(n_1346), .Y(n_1345) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_355), .A2(n_366), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_355), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_355), .A2(n_366), .B1(n_865), .B2(n_866), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g952 ( .A1(n_355), .A2(n_715), .B1(n_953), .B2(n_954), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_355), .A2(n_715), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_355), .A2(n_366), .B1(n_1338), .B2(n_1339), .Y(n_1337) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
AND2x4_ASAP7_75t_L g366 ( .A(n_356), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g553 ( .A(n_356), .Y(n_553) );
AND2x4_ASAP7_75t_L g715 ( .A(n_356), .B(n_367), .Y(n_715) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_358), .Y(n_376) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_358), .Y(n_457) );
INVx1_ASAP7_75t_L g655 ( .A(n_358), .Y(n_655) );
INVx1_ASAP7_75t_L g663 ( .A(n_358), .Y(n_663) );
BUFx2_ASAP7_75t_L g727 ( .A(n_358), .Y(n_727) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_364), .A2(n_366), .B1(n_429), .B2(n_449), .Y(n_448) );
INVx5_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx4_ASAP7_75t_L g875 ( .A(n_365), .Y(n_875) );
INVx5_ASAP7_75t_SL g542 ( .A(n_366), .Y(n_542) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_368), .Y(n_392) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_369), .Y(n_377) );
INVx3_ASAP7_75t_L g489 ( .A(n_369), .Y(n_489) );
INVx1_ASAP7_75t_L g987 ( .A(n_369), .Y(n_987) );
AOI31xp33_ASAP7_75t_L g437 ( .A1(n_371), .A2(n_438), .A3(n_445), .B(n_448), .Y(n_437) );
AOI31xp33_ASAP7_75t_L g635 ( .A1(n_371), .A2(n_636), .A3(n_638), .B(n_642), .Y(n_635) );
AND2x4_ASAP7_75t_L g419 ( .A(n_372), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g516 ( .A(n_372), .B(n_420), .Y(n_516) );
AND2x4_ASAP7_75t_L g1268 ( .A(n_372), .B(n_1269), .Y(n_1268) );
NAND4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_388), .C(n_398), .D(n_411), .Y(n_373) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .C(n_385), .Y(n_374) );
BUFx3_ASAP7_75t_L g1257 ( .A(n_376), .Y(n_1257) );
INVx2_ASAP7_75t_SL g729 ( .A(n_377), .Y(n_729) );
INVx4_ASAP7_75t_L g738 ( .A(n_377), .Y(n_738) );
INVx2_ASAP7_75t_SL g1259 ( .A(n_377), .Y(n_1259) );
BUFx3_ASAP7_75t_L g1261 ( .A(n_377), .Y(n_1261) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g454 ( .A(n_380), .Y(n_454) );
INVx2_ASAP7_75t_SL g793 ( .A(n_380), .Y(n_793) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g801 ( .A(n_381), .Y(n_801) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g652 ( .A(n_382), .Y(n_652) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_385), .B(n_452), .C(n_453), .Y(n_451) );
INVx2_ASAP7_75t_L g734 ( .A(n_385), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g787 ( .A(n_385), .B(n_788), .C(n_792), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g814 ( .A(n_385), .B(n_815), .C(n_817), .Y(n_814) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_385), .B(n_888), .C(n_889), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_385), .B(n_933), .C(n_934), .Y(n_932) );
NAND3xp33_ASAP7_75t_L g981 ( .A(n_385), .B(n_982), .C(n_983), .Y(n_981) );
BUFx3_ASAP7_75t_L g1254 ( .A(n_385), .Y(n_1254) );
AOI33xp33_ASAP7_75t_L g1356 ( .A1(n_385), .A2(n_665), .A3(n_1357), .B1(n_1360), .B2(n_1364), .B3(n_1368), .Y(n_1356) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g394 ( .A(n_386), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g408 ( .A(n_386), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g561 ( .A(n_386), .B(n_562), .Y(n_561) );
AND2x4_ASAP7_75t_L g648 ( .A(n_386), .B(n_387), .Y(n_648) );
OR2x6_ASAP7_75t_L g671 ( .A(n_386), .B(n_562), .Y(n_671) );
BUFx2_ASAP7_75t_L g1318 ( .A(n_386), .Y(n_1318) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_393), .C(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_394), .B(n_456), .C(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g501 ( .A(n_394), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_394), .B(n_891), .C(n_893), .Y(n_890) );
NAND3xp33_ASAP7_75t_L g935 ( .A(n_394), .B(n_936), .C(n_938), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g984 ( .A(n_394), .B(n_985), .C(n_988), .Y(n_984) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x6_ASAP7_75t_L g666 ( .A(n_396), .B(n_667), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_403), .C(n_407), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g686 ( .A(n_405), .Y(n_686) );
INVx1_ASAP7_75t_L g568 ( .A(n_406), .Y(n_568) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_406), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_407), .B(n_460), .C(n_463), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_407), .B(n_804), .C(n_806), .Y(n_803) );
NAND3xp33_ASAP7_75t_L g823 ( .A(n_407), .B(n_824), .C(n_826), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_407), .B(n_895), .C(n_896), .Y(n_894) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_407), .B(n_940), .C(n_941), .Y(n_939) );
NAND3xp33_ASAP7_75t_L g989 ( .A(n_407), .B(n_990), .C(n_991), .Y(n_989) );
AOI33xp33_ASAP7_75t_L g1348 ( .A1(n_407), .A2(n_1349), .A3(n_1350), .B1(n_1352), .B2(n_1354), .B3(n_1355), .Y(n_1348) );
INVx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_SL g502 ( .A1(n_408), .A2(n_503), .B1(n_515), .B2(n_517), .Y(n_502) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g562 ( .A(n_410), .Y(n_562) );
INVx2_ASAP7_75t_SL g1301 ( .A(n_410), .Y(n_1301) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .C(n_419), .Y(n_411) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g533 ( .A(n_415), .Y(n_533) );
INVx1_ASAP7_75t_L g684 ( .A(n_415), .Y(n_684) );
BUFx4f_ASAP7_75t_L g746 ( .A(n_415), .Y(n_746) );
BUFx3_ASAP7_75t_L g756 ( .A(n_415), .Y(n_756) );
INVx1_ASAP7_75t_L g772 ( .A(n_415), .Y(n_772) );
AND2x4_ASAP7_75t_L g1297 ( .A(n_415), .B(n_1277), .Y(n_1297) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_419), .B(n_465), .C(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g585 ( .A(n_419), .Y(n_585) );
AOI33xp33_ASAP7_75t_L g669 ( .A1(n_419), .A2(n_670), .A3(n_672), .B1(n_676), .B2(n_679), .B3(n_685), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_419), .B(n_809), .C(n_810), .Y(n_808) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_419), .B(n_830), .C(n_832), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_419), .B(n_898), .C(n_900), .Y(n_897) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_419), .B(n_943), .C(n_944), .Y(n_942) );
NAND3xp33_ASAP7_75t_L g992 ( .A(n_419), .B(n_993), .C(n_994), .Y(n_992) );
INVx2_ASAP7_75t_L g1293 ( .A(n_420), .Y(n_1293) );
AND2x4_ASAP7_75t_L g1270 ( .A(n_421), .B(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g802 ( .A(n_441), .Y(n_802) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g1363 ( .A(n_442), .Y(n_1363) );
INVx1_ASAP7_75t_L g784 ( .A(n_444), .Y(n_784) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_451), .B(n_455), .C(n_459), .D(n_464), .Y(n_450) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_457), .B(n_1244), .Y(n_1252) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g825 ( .A(n_462), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_557), .B1(n_613), .B2(n_614), .Y(n_467) );
INVx1_ASAP7_75t_L g613 ( .A(n_468), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_525), .C(n_540), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_502), .Y(n_470) );
OAI33xp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .A3(n_481), .B1(n_490), .B2(n_495), .B3(n_501), .Y(n_471) );
OAI33xp33_ASAP7_75t_L g586 ( .A1(n_472), .A2(n_501), .A3(n_587), .B1(n_590), .B2(n_591), .B3(n_595), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_477), .B2(n_480), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g503 ( .A1(n_476), .A2(n_480), .B1(n_504), .B2(n_509), .C(n_513), .Y(n_503) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_477), .A2(n_570), .B1(n_573), .B2(n_588), .Y(n_587) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI22xp33_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_483), .B1(n_486), .B2(n_487), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_483), .A2(n_491), .B1(n_492), .B2(n_494), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_483), .A2(n_492), .B1(n_564), .B2(n_567), .Y(n_590) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g592 ( .A(n_484), .Y(n_592) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g554 ( .A(n_485), .Y(n_554) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g657 ( .A(n_488), .Y(n_657) );
INVx2_ASAP7_75t_L g791 ( .A(n_488), .Y(n_791) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g493 ( .A(n_489), .Y(n_493) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_489), .Y(n_799) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_492), .A2(n_592), .B1(n_593), .B2(n_594), .Y(n_591) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g1243 ( .A(n_493), .B(n_1244), .Y(n_1243) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_498), .B2(n_500), .Y(n_495) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g545 ( .A(n_499), .Y(n_545) );
INVx3_ASAP7_75t_L g597 ( .A(n_499), .Y(n_597) );
INVx2_ASAP7_75t_L g839 ( .A(n_499), .Y(n_839) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g518 ( .A(n_505), .Y(n_518) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g527 ( .A(n_506), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g572 ( .A(n_506), .Y(n_572) );
OR2x2_ASAP7_75t_L g1314 ( .A(n_506), .B(n_1278), .Y(n_1314) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_L g512 ( .A(n_507), .B(n_508), .Y(n_512) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g521 ( .A(n_512), .Y(n_521) );
BUFx4f_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
INVx1_ASAP7_75t_L g914 ( .A(n_512), .Y(n_914) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx4f_ASAP7_75t_L g760 ( .A(n_516), .Y(n_760) );
BUFx4f_ASAP7_75t_L g1349 ( .A(n_516), .Y(n_1349) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_520), .B2(n_522), .C(n_523), .Y(n_517) );
INVx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g749 ( .A(n_524), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_531), .B(n_536), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g805 ( .A(n_533), .Y(n_805) );
INVx1_ASAP7_75t_L g1351 ( .A(n_533), .Y(n_1351) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_536), .B(n_603), .Y(n_602) );
NAND4xp25_ASAP7_75t_SL g621 ( .A(n_536), .B(n_622), .C(n_628), .D(n_631), .Y(n_621) );
NAND3xp33_ASAP7_75t_SL g768 ( .A(n_536), .B(n_769), .C(n_776), .Y(n_768) );
NAND3xp33_ASAP7_75t_SL g845 ( .A(n_536), .B(n_846), .C(n_849), .Y(n_845) );
OAI31xp33_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_543), .A3(n_551), .B(n_555), .Y(n_540) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND4xp25_ASAP7_75t_SL g711 ( .A(n_546), .B(n_712), .C(n_716), .D(n_722), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g863 ( .A(n_546), .B(n_864), .C(n_867), .D(n_872), .Y(n_863) );
NAND4xp25_ASAP7_75t_L g959 ( .A(n_546), .B(n_960), .C(n_963), .D(n_967), .Y(n_959) );
NAND4xp25_ASAP7_75t_SL g1336 ( .A(n_546), .B(n_1337), .C(n_1340), .D(n_1345), .Y(n_1336) );
AOI222xp33_ASAP7_75t_L g716 ( .A1(n_548), .A2(n_706), .B1(n_708), .B2(n_717), .C1(n_718), .C2(n_719), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_548), .A2(n_773), .B1(n_775), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_548), .A2(n_784), .B1(n_869), .B2(n_870), .Y(n_908) );
AND2x4_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
AND2x4_ASAP7_75t_L g871 ( .A(n_549), .B(n_550), .Y(n_871) );
AND2x4_ASAP7_75t_L g1230 ( .A(n_549), .B(n_1231), .Y(n_1230) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
OAI31xp33_ASAP7_75t_SL g608 ( .A1(n_555), .A2(n_609), .A3(n_610), .B(n_612), .Y(n_608) );
AOI221x1_ASAP7_75t_L g693 ( .A1(n_555), .A2(n_694), .B1(n_710), .B2(n_711), .C(n_724), .Y(n_693) );
OAI31xp33_ASAP7_75t_L g780 ( .A1(n_555), .A2(n_781), .A3(n_782), .B(n_785), .Y(n_780) );
OAI31xp33_ASAP7_75t_SL g834 ( .A1(n_555), .A2(n_835), .A3(n_836), .B(n_843), .Y(n_834) );
AOI221x1_ASAP7_75t_L g862 ( .A1(n_555), .A2(n_710), .B1(n_863), .B2(n_876), .C(n_885), .Y(n_862) );
OAI31xp33_ASAP7_75t_L g903 ( .A1(n_555), .A2(n_904), .A3(n_905), .B(n_909), .Y(n_903) );
AOI221x1_ASAP7_75t_L g958 ( .A1(n_555), .A2(n_634), .B1(n_959), .B2(n_970), .C(n_980), .Y(n_958) );
AOI221x1_ASAP7_75t_L g1324 ( .A1(n_555), .A2(n_710), .B1(n_1325), .B2(n_1336), .C(n_1347), .Y(n_1324) );
CKINVDCx16_ASAP7_75t_R g555 ( .A(n_556), .Y(n_555) );
AOI31xp33_ASAP7_75t_L g947 ( .A1(n_556), .A2(n_948), .A3(n_952), .B(n_955), .Y(n_947) );
INVx1_ASAP7_75t_L g614 ( .A(n_557), .Y(n_614) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_599), .C(n_608), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_586), .Y(n_559) );
OAI33xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .A3(n_569), .B1(n_576), .B2(n_579), .B3(n_585), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_567), .B2(n_568), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx4f_ASAP7_75t_L g673 ( .A(n_566), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_571), .A2(n_574), .B1(n_577), .B2(n_578), .Y(n_576) );
OAI221xp5_ASAP7_75t_L g1290 ( .A1(n_571), .A2(n_1246), .B1(n_1249), .B2(n_1291), .C(n_1292), .Y(n_1290) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g1291 ( .A(n_575), .Y(n_1291) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_582), .B1(n_583), .B2(n_584), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_L g1276 ( .A(n_581), .B(n_1277), .Y(n_1276) );
BUFx3_ASAP7_75t_L g1289 ( .A(n_581), .Y(n_1289) );
INVx1_ASAP7_75t_L g750 ( .A(n_583), .Y(n_750) );
INVx1_ASAP7_75t_L g759 ( .A(n_583), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_588), .A2(n_596), .B1(n_597), .B2(n_598), .Y(n_595) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g907 ( .A(n_597), .Y(n_907) );
INVx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g705 ( .A(n_605), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_856), .B2(n_857), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AO22x1_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_764), .B1(n_854), .B2(n_855), .Y(n_617) );
INVx1_ASAP7_75t_L g854 ( .A(n_618), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_691), .B1(n_692), .B2(n_763), .Y(n_618) );
INVx1_ASAP7_75t_L g763 ( .A(n_619), .Y(n_763) );
INVx1_ASAP7_75t_L g690 ( .A(n_620), .Y(n_690) );
AOI211x1_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_634), .B(n_635), .C(n_645), .Y(n_620) );
BUFx4f_ASAP7_75t_L g707 ( .A(n_625), .Y(n_707) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_634), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_641), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_669), .Y(n_645) );
AOI33xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .A3(n_653), .B1(n_658), .B2(n_661), .B3(n_665), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g741 ( .A(n_651), .Y(n_741) );
AND2x4_ASAP7_75t_L g1250 ( .A(n_651), .B(n_1244), .Y(n_1250) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g731 ( .A(n_652), .Y(n_731) );
INVx2_ASAP7_75t_SL g1362 ( .A(n_652), .Y(n_1362) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g664 ( .A(n_657), .Y(n_664) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g789 ( .A(n_663), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_665), .B(n_736), .C(n_739), .Y(n_735) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_665), .B(n_797), .C(n_800), .Y(n_796) );
INVx5_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx6_ASAP7_75t_L g822 ( .A(n_666), .Y(n_822) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x4_ASAP7_75t_L g1244 ( .A(n_668), .B(n_1245), .Y(n_1244) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_671), .Y(n_751) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g762 ( .A(n_693), .Y(n_762) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_695), .B(n_698), .C(n_701), .D(n_709), .Y(n_694) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g1300 ( .A(n_704), .Y(n_1300) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI31xp33_ASAP7_75t_L g910 ( .A1(n_710), .A2(n_911), .A3(n_912), .B(n_916), .Y(n_910) );
AOI222xp33_ASAP7_75t_L g867 ( .A1(n_717), .A2(n_794), .B1(n_868), .B2(n_869), .C1(n_870), .C2(n_871), .Y(n_867) );
AOI222xp33_ASAP7_75t_L g1340 ( .A1(n_717), .A2(n_871), .B1(n_1341), .B2(n_1342), .C1(n_1343), .C2(n_1344), .Y(n_1340) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g732 ( .A(n_720), .Y(n_732) );
INVx1_ASAP7_75t_L g1342 ( .A(n_720), .Y(n_1342) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g963 ( .A1(n_721), .A2(n_784), .B1(n_871), .B2(n_964), .C1(n_965), .C2(n_966), .Y(n_963) );
AND2x4_ASAP7_75t_L g1239 ( .A(n_721), .B(n_1231), .Y(n_1239) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_725), .B(n_735), .C(n_742), .D(n_752), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_730), .C(n_733), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .C(n_751), .Y(n_742) );
INVx4_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g899 ( .A(n_745), .Y(n_899) );
INVx2_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_757), .C(n_760), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g855 ( .A(n_764), .Y(n_855) );
XOR2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_811), .Y(n_764) );
NAND3x1_ASAP7_75t_L g766 ( .A(n_767), .B(n_780), .C(n_786), .Y(n_766) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g848 ( .A(n_772), .Y(n_848) );
AND4x1_ASAP7_75t_L g786 ( .A(n_787), .B(n_796), .C(n_803), .D(n_808), .Y(n_786) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
BUFx6f_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g1370 ( .A(n_795), .Y(n_1370) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g816 ( .A(n_799), .Y(n_816) );
INVx2_ASAP7_75t_L g820 ( .A(n_799), .Y(n_820) );
INVx3_ASAP7_75t_L g892 ( .A(n_799), .Y(n_892) );
INVx2_ASAP7_75t_SL g937 ( .A(n_799), .Y(n_937) );
XOR2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_853), .Y(n_811) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_834), .C(n_844), .Y(n_812) );
AND4x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_818), .C(n_823), .D(n_829), .Y(n_813) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_821), .C(n_822), .Y(n_818) );
AOI33xp33_ASAP7_75t_L g1253 ( .A1(n_822), .A2(n_1254), .A3(n_1255), .B1(n_1256), .B2(n_1260), .B3(n_1262), .Y(n_1253) );
BUFx2_ASAP7_75t_L g1303 ( .A(n_825), .Y(n_1303) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVxp67_ASAP7_75t_SL g856 ( .A(n_857), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .B1(n_957), .B2(n_997), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
AO22x2_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B1(n_917), .B2(n_918), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g909 ( .A(n_864), .Y(n_909) );
INVx1_ASAP7_75t_L g904 ( .A(n_872), .Y(n_904) );
INVxp67_ASAP7_75t_L g911 ( .A(n_877), .Y(n_911) );
INVxp67_ASAP7_75t_L g916 ( .A(n_883), .Y(n_916) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_886), .B(n_903), .C(n_910), .Y(n_902) );
AND4x1_ASAP7_75t_L g886 ( .A(n_887), .B(n_890), .C(n_894), .D(n_897), .Y(n_886) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g1329 ( .A(n_914), .Y(n_1329) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
NAND4xp25_ASAP7_75t_L g931 ( .A(n_932), .B(n_935), .C(n_939), .D(n_942), .Y(n_931) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g997 ( .A(n_957), .Y(n_997) );
INVx1_ASAP7_75t_L g996 ( .A(n_958), .Y(n_996) );
NAND3xp33_ASAP7_75t_L g970 ( .A(n_971), .B(n_975), .C(n_977), .Y(n_970) );
BUFx6f_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
AND2x4_ASAP7_75t_L g1308 ( .A(n_973), .B(n_1309), .Y(n_1308) );
NAND4xp25_ASAP7_75t_L g980 ( .A(n_981), .B(n_984), .C(n_989), .D(n_992), .Y(n_980) );
INVx1_ASAP7_75t_L g1359 ( .A(n_986), .Y(n_1359) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
INVx1_ASAP7_75t_L g1367 ( .A(n_987), .Y(n_1367) );
OAI21xp33_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1221), .B(n_1222), .Y(n_998) );
NOR2x1_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1171), .Y(n_999) );
NAND3xp33_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1104), .C(n_1148), .Y(n_1000) );
AOI211xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1029), .B(n_1068), .C(n_1099), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1002), .B(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1002), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1022), .Y(n_1002) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1003), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1003), .B(n_1066), .Y(n_1088) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1003), .Y(n_1103) );
BUFx6f_ASAP7_75t_L g1118 ( .A(n_1003), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1003), .B(n_1061), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1016), .Y(n_1003) );
AND2x4_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1011), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_1007), .B(n_1012), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1010), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_1008), .Y(n_1381) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1010), .Y(n_1019) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_1011), .B(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1060 ( .A(n_1012), .B(n_1015), .Y(n_1060) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1017), .Y(n_1025) );
BUFx3_ASAP7_75t_L g1091 ( .A(n_1017), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1020), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_1018), .B(n_1020), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1379 ( .A(n_1018), .Y(n_1379) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_1019), .B(n_1020), .Y(n_1021) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1021), .Y(n_1027) );
CKINVDCx6p67_ASAP7_75t_R g1084 ( .A(n_1022), .Y(n_1084) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1022), .B(n_1103), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1022), .B(n_1103), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1022), .B(n_1139), .Y(n_1138) );
CKINVDCx5p33_ASAP7_75t_R g1183 ( .A(n_1022), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1022), .B(n_1216), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1022), .B(n_1080), .Y(n_1220) );
OR2x6_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_1023), .B(n_1024), .Y(n_1123) );
OAI22xp5_ASAP7_75t_SL g1024 ( .A1(n_1025), .A2(n_1026), .B1(n_1027), .B2(n_1028), .Y(n_1024) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1027), .Y(n_1053) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1027), .Y(n_1092) );
A2O1A1Ixp33_ASAP7_75t_L g1029 ( .A1(n_1030), .A2(n_1044), .B(n_1050), .C(n_1064), .Y(n_1029) );
NOR2xp33_ASAP7_75t_L g1219 ( .A(n_1030), .B(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1036), .Y(n_1031) );
CKINVDCx5p33_ASAP7_75t_R g1046 ( .A(n_1032), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1032), .B(n_1047), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_1032), .B(n_1087), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1032), .B(n_1072), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1032), .B(n_1126), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1032), .B(n_1087), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1032), .B(n_1051), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1032), .B(n_1206), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1032), .B(n_1121), .Y(n_1210) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1032), .B(n_1206), .Y(n_1213) );
AND2x4_ASAP7_75t_SL g1032 ( .A(n_1033), .B(n_1034), .Y(n_1032) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1036), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1036), .B(n_1046), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1040), .Y(n_1036) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1037), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1037), .B(n_1041), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
INVxp67_ASAP7_75t_SL g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1041), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1041), .B(n_1048), .Y(n_1121) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1041), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .Y(n_1041) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1045), .B(n_1101), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1045), .B(n_1070), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1179 ( .A1(n_1045), .A2(n_1139), .B1(n_1156), .B2(n_1180), .C(n_1182), .Y(n_1179) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_1045), .B(n_1113), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1047), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1046), .B(n_1072), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1046), .B(n_1077), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1119 ( .A(n_1046), .B(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1046), .B(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1046), .B(n_1121), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1046), .B(n_1052), .Y(n_1162) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1047), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1047), .B(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1047), .B(n_1170), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1049), .Y(n_1047) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1048), .Y(n_1087) );
OAI322xp33_ASAP7_75t_L g1124 ( .A1(n_1050), .A2(n_1125), .A3(n_1127), .B1(n_1129), .B2(n_1130), .C1(n_1131), .C2(n_1133), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1061), .Y(n_1050) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_1051), .B(n_1066), .Y(n_1065) );
BUFx3_ASAP7_75t_L g1070 ( .A(n_1051), .Y(n_1070) );
INVx2_ASAP7_75t_SL g1078 ( .A(n_1051), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_1051), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1051), .B(n_1156), .Y(n_1155) );
INVx2_ASAP7_75t_SL g1051 ( .A(n_1052), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1052), .B(n_1066), .Y(n_1139) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .B1(n_1058), .B2(n_1059), .Y(n_1054) );
BUFx3_ASAP7_75t_L g1095 ( .A(n_1056), .Y(n_1095) );
BUFx6f_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1060), .Y(n_1098) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1061), .Y(n_1066) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1061), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1061), .B(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1061), .Y(n_1156) );
NAND3xp33_ASAP7_75t_L g1163 ( .A(n_1061), .B(n_1164), .C(n_1166), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1063), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1067), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1065), .B(n_1072), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1066), .B(n_1084), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1066), .B(n_1081), .Y(n_1159) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1067), .Y(n_1108) );
A2O1A1Ixp33_ASAP7_75t_L g1186 ( .A1(n_1067), .A2(n_1123), .B(n_1152), .C(n_1187), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1067), .B(n_1192), .Y(n_1191) );
OAI211xp5_ASAP7_75t_L g1211 ( .A1(n_1067), .A2(n_1212), .B(n_1214), .C(n_1217), .Y(n_1211) );
OAI221xp5_ASAP7_75t_L g1068 ( .A1(n_1069), .A2(n_1073), .B1(n_1075), .B2(n_1080), .C(n_1082), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1071), .Y(n_1069) );
NOR3xp33_ASAP7_75t_L g1089 ( .A(n_1070), .B(n_1087), .C(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1070), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1070), .B(n_1159), .Y(n_1198) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1072), .Y(n_1134) );
A2O1A1Ixp33_ASAP7_75t_L g1184 ( .A1(n_1073), .A2(n_1125), .B(n_1185), .C(n_1186), .Y(n_1184) );
OAI211xp5_ASAP7_75t_SL g1173 ( .A1(n_1074), .A2(n_1174), .B(n_1176), .C(n_1179), .Y(n_1173) );
INVx3_ASAP7_75t_L g1194 ( .A(n_1074), .Y(n_1194) );
AOI21xp33_ASAP7_75t_L g1099 ( .A1(n_1075), .A2(n_1100), .B(n_1102), .Y(n_1099) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
NOR2xp33_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1079), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1078), .B(n_1086), .Y(n_1085) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1078), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1078), .B(n_1121), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1078), .B(n_1205), .Y(n_1204) );
INVxp67_ASAP7_75t_L g1216 ( .A(n_1078), .Y(n_1216) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1080), .Y(n_1132) );
INVx2_ASAP7_75t_L g1217 ( .A(n_1080), .Y(n_1217) );
AOI22xp5_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1085), .B1(n_1088), .B2(n_1089), .Y(n_1082) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1083), .Y(n_1109) );
NOR2xp33_ASAP7_75t_L g1114 ( .A(n_1084), .B(n_1115), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1084), .B(n_1088), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1084), .B(n_1103), .Y(n_1203) );
NAND2xp5_ASAP7_75t_SL g1208 ( .A(n_1084), .B(n_1159), .Y(n_1208) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1086), .Y(n_1130) );
AOI222xp33_ASAP7_75t_L g1176 ( .A1(n_1087), .A2(n_1121), .B1(n_1151), .B2(n_1159), .C1(n_1177), .C2(n_1178), .Y(n_1176) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1087), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1088), .B(n_1128), .Y(n_1140) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1088), .Y(n_1201) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1090), .Y(n_1147) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1092), .Y(n_1221) );
OAI22xp33_ASAP7_75t_L g1093 ( .A1(n_1094), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1093) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1101), .Y(n_1190) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1102), .Y(n_1166) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1103), .Y(n_1129) );
OAI31xp33_ASAP7_75t_SL g1104 ( .A1(n_1105), .A2(n_1114), .A3(n_1117), .B(n_1144), .Y(n_1104) );
OAI222xp33_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1107), .B1(n_1108), .B2(n_1109), .C1(n_1110), .C2(n_1112), .Y(n_1105) );
OAI321xp33_ASAP7_75t_L g1188 ( .A1(n_1107), .A2(n_1135), .A3(n_1185), .B1(n_1189), .B2(n_1190), .C(n_1191), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_1110), .A2(n_1150), .B1(n_1153), .B2(n_1154), .Y(n_1149) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1111), .B(n_1175), .Y(n_1218) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1113), .B(n_1127), .Y(n_1175) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
OAI211xp5_ASAP7_75t_SL g1117 ( .A1(n_1118), .A2(n_1119), .B(n_1122), .C(n_1141), .Y(n_1117) );
CKINVDCx14_ASAP7_75t_R g1178 ( .A(n_1118), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1121), .B(n_1162), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1124), .B1(n_1136), .B2(n_1137), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g1177 ( .A(n_1125), .B(n_1128), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1126), .B(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1126), .Y(n_1181) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1128), .B(n_1152), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1132), .B(n_1170), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1134), .B(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1136), .Y(n_1153) );
NAND2xp33_ASAP7_75t_SL g1137 ( .A(n_1138), .B(n_1140), .Y(n_1137) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1139), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1143), .Y(n_1189) );
OAI21xp33_ASAP7_75t_L g1171 ( .A1(n_1144), .A2(n_1172), .B(n_1195), .Y(n_1171) );
INVx3_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
AOI21xp5_ASAP7_75t_L g1148 ( .A1(n_1145), .A2(n_1149), .B(n_1157), .Y(n_1148) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
NOR2xp33_ASAP7_75t_L g1168 ( .A(n_1153), .B(n_1169), .Y(n_1168) );
OAI211xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1160), .B(n_1163), .C(n_1167), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
AOI211xp5_ASAP7_75t_L g1172 ( .A1(n_1173), .A2(n_1183), .B(n_1184), .C(n_1188), .Y(n_1172) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
NOR3xp33_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1207), .C(n_1219), .Y(n_1195) );
OAI221xp5_ASAP7_75t_SL g1196 ( .A1(n_1197), .A2(n_1198), .B1(n_1199), .B2(n_1201), .C(n_1202), .Y(n_1196) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1203), .B(n_1204), .Y(n_1202) );
OAI211xp5_ASAP7_75t_SL g1207 ( .A1(n_1208), .A2(n_1209), .B(n_1211), .C(n_1218), .Y(n_1207) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
HB1xp67_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1263), .Y(n_1225) );
AND4x1_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1240), .C(n_1248), .D(n_1253), .Y(n_1226) );
AOI221xp5_ASAP7_75t_L g1227 ( .A1(n_1228), .A2(n_1234), .B1(n_1235), .B2(n_1237), .C(n_1238), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
AND2x4_ASAP7_75t_L g1235 ( .A(n_1231), .B(n_1236), .Y(n_1235) );
INVx3_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
HB1xp67_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_1241), .A2(n_1242), .B1(n_1246), .B2(n_1247), .Y(n_1240) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_1249), .A2(n_1250), .B1(n_1251), .B2(n_1252), .Y(n_1248) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
AOI21xp33_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1273), .B(n_1274), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1267), .Y(n_1265) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
AND2x4_ASAP7_75t_L g1282 ( .A(n_1270), .B(n_1283), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1270), .B(n_1287), .Y(n_1286) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1270), .Y(n_1310) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
AOI31xp33_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1294), .A3(n_1311), .B(n_1318), .Y(n_1274) );
AOI211xp5_ASAP7_75t_L g1275 ( .A1(n_1276), .A2(n_1279), .B(n_1280), .C(n_1288), .Y(n_1275) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1278), .B(n_1307), .Y(n_1317) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx2_ASAP7_75t_SL g1285 ( .A(n_1286), .Y(n_1285) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
AOI221xp5_ASAP7_75t_L g1294 ( .A1(n_1295), .A2(n_1298), .B1(n_1299), .B2(n_1302), .C(n_1308), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1305), .Y(n_1353) );
INVx2_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_SL g1309 ( .A(n_1310), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1313), .B1(n_1315), .B2(n_1316), .Y(n_1311) );
INVx6_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
INVx4_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
BUFx2_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1322), .Y(n_1371) );
HB1xp67_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
NAND3xp33_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1330), .C(n_1333), .Y(n_1325) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1348), .B(n_1356), .Y(n_1347) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
BUFx2_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
CKINVDCx5p33_ASAP7_75t_R g1374 ( .A(n_1375), .Y(n_1374) );
A2O1A1Ixp33_ASAP7_75t_L g1377 ( .A1(n_1376), .A2(n_1378), .B(n_1380), .C(n_1382), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
endmodule