module fake_jpeg_29519_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_53),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_43),
.B1(n_52),
.B2(n_49),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_48),
.B1(n_53),
.B2(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_73),
.B1(n_44),
.B2(n_3),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_61),
.B1(n_58),
.B2(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_1),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_51),
.B1(n_46),
.B2(n_41),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_45),
.C(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_19),
.B(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_45),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_90),
.B(n_3),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_2),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_89),
.B1(n_7),
.B2(n_9),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_70),
.A2(n_32),
.B1(n_14),
.B2(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_2),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_87),
.B(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_86),
.A2(n_74),
.B1(n_66),
.B2(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_97),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_94),
.B(n_9),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_81),
.B1(n_83),
.B2(n_91),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_101),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_22),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_106),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_7),
.B(n_8),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_12),
.B(n_13),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_110),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_10),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_113),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_20),
.B(n_25),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_101),
.C(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_107),
.C(n_103),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_121),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_115),
.B(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_123),
.C(n_112),
.Y(n_128)
);

AOI211xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_112),
.B(n_114),
.C(n_118),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_102),
.B(n_27),
.Y(n_130)
);


endmodule