module fake_jpeg_15580_n_383 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_383);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_383;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_8),
.B1(n_12),
.B2(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_49),
.B1(n_37),
.B2(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_42),
.B(n_47),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_15),
.B(n_8),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_13),
.B1(n_8),
.B2(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_22),
.B(n_9),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_37),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_61),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_15),
.B(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_30),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_17),
.B1(n_25),
.B2(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_66),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_67),
.B(n_71),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_68),
.A2(n_83),
.B1(n_77),
.B2(n_80),
.Y(n_165)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_17),
.B1(n_30),
.B2(n_14),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_17),
.B1(n_25),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_17),
.B1(n_14),
.B2(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_76),
.B(n_82),
.Y(n_166)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_80),
.B(n_91),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_14),
.B1(n_30),
.B2(n_31),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_84),
.A2(n_95),
.B1(n_115),
.B2(n_5),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_20),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_23),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_25),
.B1(n_22),
.B2(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_29),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_101),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_44),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_106),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_46),
.B(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_26),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_26),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_24),
.B1(n_29),
.B2(n_35),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_9),
.B1(n_12),
.B2(n_5),
.Y(n_133)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_55),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_114),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_24),
.B1(n_35),
.B2(n_28),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_113),
.B(n_129),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_28),
.B1(n_23),
.B2(n_16),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_20),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_118),
.B(n_129),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_24),
.B1(n_28),
.B2(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_121),
.A2(n_128),
.B1(n_137),
.B2(n_146),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_36),
.B1(n_16),
.B2(n_18),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_122),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_148),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_105),
.B1(n_88),
.B2(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_167),
.B1(n_102),
.B2(n_113),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_16),
.B1(n_36),
.B2(n_18),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_20),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_36),
.B1(n_18),
.B2(n_5),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_36),
.B(n_10),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_131),
.A2(n_145),
.B(n_151),
.Y(n_188)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_81),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_6),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_138),
.B(n_149),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_77),
.A2(n_13),
.B1(n_0),
.B2(n_1),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_13),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_147),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_87),
.A2(n_0),
.B1(n_1),
.B2(n_92),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_79),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_159),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_157),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_99),
.A2(n_1),
.B1(n_105),
.B2(n_87),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_165),
.B1(n_117),
.B2(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_72),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_112),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_91),
.A2(n_1),
.B(n_70),
.C(n_114),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_162),
.A2(n_101),
.B(n_90),
.C(n_98),
.Y(n_168)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_89),
.B(n_97),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_102),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_83),
.A2(n_89),
.B1(n_97),
.B2(n_98),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_170),
.A2(n_176),
.B1(n_181),
.B2(n_195),
.Y(n_227)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_203),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_179),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_126),
.B1(n_165),
.B2(n_166),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_116),
.B1(n_118),
.B2(n_167),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_179),
.A2(n_191),
.B1(n_193),
.B2(n_197),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_147),
.C(n_140),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_190),
.C(n_183),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_178),
.C(n_177),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_116),
.B(n_142),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_190),
.B(n_196),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_142),
.B1(n_159),
.B2(n_140),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_160),
.B1(n_162),
.B2(n_153),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_154),
.A2(n_160),
.B1(n_138),
.B2(n_146),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_133),
.B(n_137),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_119),
.A2(n_124),
.B1(n_143),
.B2(n_132),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_124),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_201),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_207),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_156),
.A2(n_158),
.B1(n_120),
.B2(n_135),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

BUFx4f_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_139),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_210),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_144),
.B(n_149),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_123),
.B(n_142),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_217),
.A2(n_233),
.B(n_226),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_171),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_223),
.B(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_194),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_175),
.B(n_183),
.C(n_207),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_226),
.B(n_229),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_177),
.Y(n_229)
);

NAND2x1_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_209),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_237),
.Y(n_263)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_185),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_174),
.B(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_244),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_171),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_186),
.B(n_172),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_247),
.B(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_172),
.B(n_206),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_192),
.A2(n_180),
.B(n_181),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_253),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_192),
.A2(n_200),
.B(n_202),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_238),
.A2(n_212),
.B1(n_169),
.B2(n_208),
.Y(n_259)
);

OAI22x1_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_286),
.B1(n_269),
.B2(n_282),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_260),
.B(n_265),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_261),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_170),
.B1(n_169),
.B2(n_189),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_232),
.B1(n_228),
.B2(n_223),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_246),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_275),
.Y(n_290)
);

OA22x2_ASAP7_75t_L g269 ( 
.A1(n_233),
.A2(n_204),
.B1(n_173),
.B2(n_189),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_269),
.A2(n_239),
.B(n_252),
.C(n_230),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_214),
.B(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_270),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_240),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_282),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_249),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_215),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_285),
.C(n_248),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_227),
.A2(n_250),
.B1(n_247),
.B2(n_218),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_240),
.B1(n_255),
.B2(n_277),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_231),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_284),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_220),
.A2(n_233),
.B1(n_218),
.B2(n_243),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_251),
.B1(n_253),
.B2(n_241),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_234),
.B(n_219),
.Y(n_282)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_225),
.B(n_229),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_287),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_257),
.Y(n_326)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_292),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_294),
.A2(n_298),
.B1(n_306),
.B2(n_307),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_308),
.Y(n_325)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_310),
.B1(n_301),
.B2(n_295),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_277),
.A2(n_232),
.B1(n_228),
.B2(n_245),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_299),
.A2(n_301),
.B(n_265),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_216),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_313),
.C(n_264),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_274),
.B(n_230),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_311),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_255),
.A2(n_236),
.B1(n_238),
.B2(n_267),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_238),
.B1(n_262),
.B2(n_278),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_310),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_256),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_280),
.A2(n_262),
.B1(n_269),
.B2(n_271),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_271),
.B1(n_273),
.B2(n_283),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_264),
.B(n_285),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_256),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_260),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_315),
.A2(n_335),
.B1(n_334),
.B2(n_329),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_290),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_316),
.B1(n_328),
.B2(n_291),
.Y(n_340)
);

NAND2xp33_ASAP7_75t_SL g349 ( 
.A(n_319),
.B(n_303),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_321),
.C(n_322),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_273),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_257),
.Y(n_322)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_281),
.C(n_268),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_326),
.C(n_334),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_327),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_288),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_275),
.C(n_279),
.Y(n_334)
);

XOR2x1_ASAP7_75t_SL g339 ( 
.A(n_319),
.B(n_312),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_339),
.B(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_287),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_344),
.C(n_347),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_299),
.B1(n_309),
.B2(n_308),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_348),
.B1(n_339),
.B2(n_344),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_306),
.C(n_292),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_335),
.A2(n_294),
.B1(n_299),
.B2(n_298),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_345),
.A2(n_349),
.B1(n_331),
.B2(n_332),
.Y(n_362)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_300),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_299),
.B1(n_296),
.B2(n_288),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_345),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_324),
.C(n_315),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_352),
.C(n_331),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_330),
.C(n_328),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_341),
.B(n_325),
.CI(n_330),
.CON(n_353),
.SN(n_353)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_353),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_354),
.A2(n_364),
.B(n_347),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_359),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_333),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_362),
.Y(n_368)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_348),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_361),
.A2(n_363),
.B(n_343),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_352),
.B(n_336),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_366),
.A2(n_364),
.B(n_356),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_367),
.B1(n_354),
.B2(n_361),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_338),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_359),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_371),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_373),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_368),
.A2(n_356),
.B1(n_363),
.B2(n_357),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_375),
.A2(n_365),
.B1(n_351),
.B2(n_338),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_378),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_374),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_358),
.C(n_374),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_358),
.C(n_369),
.Y(n_381)
);

AOI21x1_ASAP7_75t_L g382 ( 
.A1(n_381),
.A2(n_366),
.B(n_337),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_382),
.B(n_337),
.Y(n_383)
);


endmodule