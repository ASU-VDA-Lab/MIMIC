module fake_jpeg_1119_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_55),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_52),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_0),
.Y(n_60)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_55),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_82),
.B1(n_38),
.B2(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_40),
.B1(n_68),
.B2(n_51),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_39),
.B1(n_43),
.B2(n_48),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_48),
.B1(n_43),
.B2(n_42),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_66),
.B(n_68),
.C(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_38),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_63),
.B1(n_64),
.B2(n_49),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_96),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_8),
.B(n_9),
.Y(n_110)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g112 ( 
.A(n_93),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_18),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_41),
.B1(n_50),
.B2(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_98),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_10),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_5),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_20),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_11),
.B1(n_12),
.B2(n_36),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_111),
.B(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_11),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_27),
.B1(n_35),
.B2(n_17),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_12),
.B1(n_24),
.B2(n_28),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_123),
.B1(n_127),
.B2(n_112),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_32),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_108),
.C(n_112),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_19),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_30),
.B1(n_109),
.B2(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_129),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_132),
.C(n_118),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_124),
.B(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_137),
.B(n_135),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_117),
.C(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_128),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_117),
.B(n_120),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_127),
.Y(n_143)
);


endmodule