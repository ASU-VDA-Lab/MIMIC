module fake_netlist_5_2000_n_1093 (n_137, n_210, n_168, n_260, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_268, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_271, n_46, n_233, n_21, n_94, n_203, n_245, n_274, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_267, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_272, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_273, n_270, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_1093);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_268;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_271;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_274;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_272;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_273;
input n_270;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1093;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_318;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_315;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_913;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_1055;
wire n_916;
wire n_452;
wire n_1081;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_718;
wire n_671;
wire n_819;
wire n_302;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_932;
wire n_417;
wire n_946;
wire n_1048;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_757;
wire n_936;
wire n_1090;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_1063;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_943;
wire n_524;
wire n_878;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_992;
wire n_1049;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_919;
wire n_782;
wire n_325;
wire n_449;
wire n_1073;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_1062;
wire n_400;
wire n_962;
wire n_436;
wire n_930;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_482;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_477;
wire n_338;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1028;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_585;
wire n_349;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_1091;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_425;
wire n_513;
wire n_647;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_952;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_931;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_803;
wire n_868;
wire n_1092;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_1004;
wire n_935;
wire n_817;
wire n_1032;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_36),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_129),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_150),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_48),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_126),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_141),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_39),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_39),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_118),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_58),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_143),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_74),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_149),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_101),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_208),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_25),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_234),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_12),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_114),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_72),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_163),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_216),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_273),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_49),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_115),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_6),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_188),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_103),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_170),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_96),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_90),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_241),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_217),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_30),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_24),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_225),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_159),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_125),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_66),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_124),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_75),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_8),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_256),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_182),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_60),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_104),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_218),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_3),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_250),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_32),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_229),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_97),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_148),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_19),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_2),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_174),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_248),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_28),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_276),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_281),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_275),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_282),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_334),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_281),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_277),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_0),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_310),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_312),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_280),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_310),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_327),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_333),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_295),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_295),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_296),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_278),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_307),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_307),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_283),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_0),
.Y(n_373)
);

INVxp33_ASAP7_75t_SL g374 ( 
.A(n_313),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_285),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_279),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_287),
.B(n_1),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_291),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_288),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_371),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_365),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_341),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_370),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_376),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_378),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_363),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_339),
.B(n_335),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_362),
.B(n_322),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_375),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_343),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_364),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_337),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_337),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_381),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_342),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_342),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_344),
.B(n_314),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_347),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_347),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_352),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_354),
.B(n_289),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_346),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_352),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_356),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_356),
.B(n_290),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_357),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_367),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

BUFx10_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_353),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_294),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_318),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_393),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_395),
.B(n_351),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_411),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_411),
.A2(n_299),
.B1(n_300),
.B2(n_298),
.Y(n_444)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_428),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_382),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_412),
.B(n_302),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_304),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_425),
.A2(n_306),
.B1(n_309),
.B2(n_308),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_305),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_425),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

INVx6_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_403),
.A2(n_305),
.B1(n_328),
.B2(n_326),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_387),
.B(n_311),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_398),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_428),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_398),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

NOR2x1p5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_315),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_410),
.B(n_360),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_384),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_407),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_404),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_404),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_423),
.B(n_332),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_SL g474 ( 
.A(n_426),
.B(n_355),
.C(n_317),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_418),
.A2(n_305),
.B1(n_319),
.B2(n_316),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_417),
.B(n_320),
.Y(n_478)
);

NAND3xp33_ASAP7_75t_L g479 ( 
.A(n_405),
.B(n_324),
.C(n_323),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_390),
.Y(n_480)
);

AND3x2_ASAP7_75t_L g481 ( 
.A(n_422),
.B(n_1),
.C(n_2),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_422),
.B(n_361),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_412),
.B(n_305),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_417),
.B(n_325),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_412),
.B(n_336),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_412),
.B(n_305),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_427),
.B(n_331),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_427),
.B(n_330),
.Y(n_492)
);

BUFx10_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_414),
.B(n_47),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_414),
.B(n_3),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

O2A1O1Ixp5_ASAP7_75t_L g498 ( 
.A1(n_453),
.A2(n_420),
.B(n_414),
.C(n_415),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_466),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_414),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_462),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_420),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_431),
.B(n_434),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_470),
.A2(n_415),
.B1(n_416),
.B2(n_409),
.Y(n_505)
);

BUFx5_ASAP7_75t_L g506 ( 
.A(n_487),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_480),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_434),
.B(n_430),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_476),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_454),
.B(n_430),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_442),
.A2(n_430),
.B(n_421),
.C(n_424),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_468),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_496),
.B(n_430),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_475),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_454),
.B(n_430),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_441),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_490),
.B(n_416),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_435),
.B(n_421),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_470),
.A2(n_424),
.B1(n_385),
.B2(n_396),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_472),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_490),
.B(n_383),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_496),
.A2(n_385),
.B1(n_396),
.B2(n_383),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_401),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_435),
.B(n_50),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_438),
.B(n_51),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_478),
.A2(n_401),
.B1(n_419),
.B2(n_53),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_494),
.B(n_4),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_491),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_469),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_466),
.B(n_5),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_448),
.B(n_7),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_438),
.B(n_52),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_432),
.B(n_7),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_491),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_433),
.B(n_10),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_482),
.B(n_11),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_485),
.B(n_54),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_463),
.A2(n_56),
.B1(n_57),
.B2(n_55),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g542 ( 
.A(n_474),
.B(n_59),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_466),
.B(n_11),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_455),
.A2(n_62),
.B1(n_63),
.B2(n_61),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_445),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

INVxp33_ASAP7_75t_L g547 ( 
.A(n_464),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_477),
.A2(n_65),
.B1(n_67),
.B2(n_64),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_459),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_459),
.B(n_68),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_473),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_445),
.B(n_12),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_449),
.B(n_13),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_495),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_461),
.B(n_69),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_451),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_461),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_444),
.B(n_14),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_443),
.B(n_70),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_458),
.B(n_15),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_447),
.B(n_16),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_436),
.B(n_71),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_457),
.B(n_73),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_486),
.B(n_16),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_452),
.B(n_76),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_452),
.B(n_77),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_502),
.B(n_483),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_557),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_560),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_500),
.A2(n_484),
.B(n_479),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_503),
.A2(n_509),
.B(n_526),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_547),
.B(n_560),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_521),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_497),
.B(n_501),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_527),
.A2(n_440),
.B(n_451),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_513),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_508),
.B(n_484),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_558),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_510),
.B(n_533),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_519),
.A2(n_460),
.B1(n_465),
.B2(n_451),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_533),
.B(n_487),
.Y(n_585)
);

AOI21x1_ASAP7_75t_L g586 ( 
.A1(n_540),
.A2(n_440),
.B(n_446),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_499),
.B(n_481),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_498),
.A2(n_487),
.B(n_450),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_531),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_534),
.A2(n_450),
.B(n_446),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_535),
.B(n_450),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_505),
.B(n_439),
.Y(n_592)
);

O2A1O1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_554),
.A2(n_450),
.B(n_19),
.C(n_17),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_L g594 ( 
.A1(n_559),
.A2(n_460),
.B(n_437),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_529),
.Y(n_595)
);

AO32x1_ASAP7_75t_L g596 ( 
.A1(n_548),
.A2(n_17),
.A3(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_535),
.A2(n_446),
.B(n_437),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_564),
.A2(n_79),
.B(n_78),
.Y(n_598)
);

O2A1O1Ixp33_ASAP7_75t_L g599 ( 
.A1(n_559),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_564),
.A2(n_81),
.B(n_80),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_568),
.Y(n_601)
);

INVx6_ASAP7_75t_L g602 ( 
.A(n_514),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_511),
.A2(n_83),
.B(n_82),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_536),
.B(n_467),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_546),
.B(n_467),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_516),
.A2(n_565),
.B(n_569),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_549),
.B(n_493),
.Y(n_607)
);

AND2x4_ASAP7_75t_SL g608 ( 
.A(n_545),
.B(n_493),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_567),
.A2(n_85),
.B(n_84),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_556),
.A2(n_87),
.B(n_86),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_562),
.B(n_22),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_562),
.A2(n_89),
.B(n_88),
.Y(n_612)
);

O2A1O1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_553),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_613)
);

AO22x1_ASAP7_75t_L g614 ( 
.A1(n_563),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_515),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_556),
.A2(n_92),
.B(n_91),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_550),
.A2(n_94),
.B(n_93),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_512),
.A2(n_176),
.B1(n_272),
.B2(n_271),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_517),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_520),
.A2(n_98),
.B(n_95),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_522),
.B(n_26),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_555),
.A2(n_100),
.B(n_99),
.Y(n_622)
);

A2O1A1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_563),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_524),
.B(n_566),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_539),
.B(n_566),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_L g626 ( 
.A(n_541),
.B(n_102),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_514),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_551),
.B(n_27),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_561),
.A2(n_106),
.B(n_105),
.Y(n_629)
);

O2A1O1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_532),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_504),
.A2(n_108),
.B(n_107),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_570),
.B(n_538),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_595),
.B(n_518),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_584),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_574),
.A2(n_561),
.B(n_525),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_606),
.A2(n_523),
.B(n_507),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_591),
.A2(n_529),
.B(n_528),
.Y(n_638)
);

AOI21x1_ASAP7_75t_L g639 ( 
.A1(n_586),
.A2(n_542),
.B(n_543),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_595),
.B(n_552),
.Y(n_640)
);

NOR2x1_ASAP7_75t_SL g641 ( 
.A(n_573),
.B(n_506),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_602),
.Y(n_642)
);

AOI221x1_ASAP7_75t_L g643 ( 
.A1(n_611),
.A2(n_537),
.B1(n_530),
.B2(n_524),
.C(n_544),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_530),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_582),
.B(n_537),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_578),
.A2(n_506),
.B(n_110),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_590),
.A2(n_506),
.B(n_111),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_585),
.A2(n_506),
.B(n_112),
.Y(n_649)
);

AOI221x1_ASAP7_75t_L g650 ( 
.A1(n_597),
.A2(n_506),
.B1(n_32),
.B2(n_33),
.C(n_34),
.Y(n_650)
);

AO31x2_ASAP7_75t_L g651 ( 
.A1(n_618),
.A2(n_506),
.A3(n_33),
.B(n_34),
.Y(n_651)
);

INVx3_ASAP7_75t_SL g652 ( 
.A(n_581),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_625),
.A2(n_187),
.B1(n_270),
.B2(n_269),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_579),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_588),
.A2(n_113),
.B(n_109),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_615),
.B(n_116),
.Y(n_656)
);

NAND3xp33_ASAP7_75t_L g657 ( 
.A(n_592),
.B(n_31),
.C(n_35),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_598),
.A2(n_119),
.B(n_117),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_601),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g660 ( 
.A1(n_612),
.A2(n_121),
.B(n_120),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_619),
.B(n_36),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_620),
.A2(n_192),
.B(n_268),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_600),
.A2(n_191),
.B(n_267),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_629),
.A2(n_190),
.B(n_266),
.Y(n_664)
);

O2A1O1Ixp5_ASAP7_75t_L g665 ( 
.A1(n_580),
.A2(n_189),
.B(n_265),
.C(n_264),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_602),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_609),
.A2(n_186),
.B(n_262),
.Y(n_667)
);

O2A1O1Ixp33_ASAP7_75t_SL g668 ( 
.A1(n_623),
.A2(n_185),
.B(n_261),
.C(n_260),
.Y(n_668)
);

A2O1A1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_626),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_583),
.B(n_274),
.Y(n_670)
);

AOI21x1_ASAP7_75t_L g671 ( 
.A1(n_628),
.A2(n_183),
.B(n_258),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_621),
.A2(n_181),
.B(n_257),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_589),
.A2(n_180),
.B(n_255),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_572),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_608),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_575),
.Y(n_676)
);

AO31x2_ASAP7_75t_L g677 ( 
.A1(n_617),
.A2(n_37),
.A3(n_38),
.B(n_40),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_594),
.A2(n_184),
.B1(n_254),
.B2(n_253),
.Y(n_678)
);

A2O1A1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_613),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_613),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_602),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_593),
.A2(n_193),
.B(n_252),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_587),
.B(n_44),
.Y(n_683)
);

AOI21x1_ASAP7_75t_L g684 ( 
.A1(n_622),
.A2(n_179),
.B(n_251),
.Y(n_684)
);

O2A1O1Ixp5_ASAP7_75t_L g685 ( 
.A1(n_603),
.A2(n_178),
.B(n_249),
.C(n_247),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_610),
.A2(n_177),
.B(n_246),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_587),
.Y(n_687)
);

AOI221x1_ASAP7_75t_L g688 ( 
.A1(n_616),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.C(n_122),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_584),
.B(n_45),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_604),
.A2(n_194),
.B1(n_123),
.B2(n_127),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_645),
.A2(n_599),
.B(n_630),
.C(n_607),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_636),
.B(n_605),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_681),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_676),
.B(n_627),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_636),
.B(n_614),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_644),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_681),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_632),
.B(n_576),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_669),
.A2(n_679),
.B(n_680),
.C(n_599),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_654),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_659),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_681),
.B(n_631),
.Y(n_702)
);

NAND2x1p5_ASAP7_75t_L g703 ( 
.A(n_642),
.B(n_593),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_640),
.B(n_46),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_633),
.B(n_630),
.Y(n_705)
);

BUFx2_ASAP7_75t_SL g706 ( 
.A(n_675),
.Y(n_706)
);

CKINVDCx11_ASAP7_75t_R g707 ( 
.A(n_652),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_674),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_643),
.A2(n_596),
.B1(n_130),
.B2(n_131),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_687),
.B(n_128),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_674),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_646),
.B(n_132),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_635),
.A2(n_596),
.B(n_134),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_682),
.A2(n_596),
.B1(n_135),
.B2(n_136),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_660),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_687),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_683),
.B(n_139),
.Y(n_717)
);

AO21x2_ASAP7_75t_L g718 ( 
.A1(n_638),
.A2(n_140),
.B(n_142),
.Y(n_718)
);

BUFx2_ASAP7_75t_SL g719 ( 
.A(n_642),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_670),
.B(n_144),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_642),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_639),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_666),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_670),
.B(n_145),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_666),
.B(n_146),
.Y(n_725)
);

AOI21xp5_ASAP7_75t_L g726 ( 
.A1(n_648),
.A2(n_147),
.B(n_151),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_666),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_664),
.B(n_152),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_637),
.A2(n_153),
.B(n_154),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_678),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_662),
.A2(n_158),
.B(n_160),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_650),
.B(n_161),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_687),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_647),
.A2(n_649),
.B(n_655),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_657),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_656),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_634),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_641),
.A2(n_169),
.B(n_171),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_661),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_656),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_689),
.B(n_172),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_703),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_740),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_740),
.Y(n_744)
);

BUFx2_ASAP7_75t_R g745 ( 
.A(n_701),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_722),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_696),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_695),
.B(n_651),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_732),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_700),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_693),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_708),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_711),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_692),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_732),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_692),
.A2(n_672),
.B1(n_690),
.B2(n_663),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_740),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_718),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_734),
.A2(n_667),
.B(n_686),
.Y(n_759)
);

OA21x2_ASAP7_75t_L g760 ( 
.A1(n_713),
.A2(n_688),
.B(n_665),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_705),
.A2(n_653),
.B1(n_656),
.B2(n_673),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_718),
.Y(n_762)
);

CKINVDCx6p67_ASAP7_75t_R g763 ( 
.A(n_707),
.Y(n_763)
);

BUFx2_ASAP7_75t_SL g764 ( 
.A(n_693),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_695),
.B(n_677),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_712),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_SL g767 ( 
.A1(n_715),
.A2(n_656),
.B1(n_658),
.B2(n_668),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_703),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_694),
.Y(n_769)
);

CKINVDCx11_ASAP7_75t_R g770 ( 
.A(n_737),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_727),
.Y(n_771)
);

OA21x2_ASAP7_75t_L g772 ( 
.A1(n_714),
.A2(n_685),
.B(n_671),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_693),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_739),
.Y(n_774)
);

AOI21x1_ASAP7_75t_L g775 ( 
.A1(n_728),
.A2(n_684),
.B(n_651),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_704),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_723),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_716),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_712),
.B(n_677),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_698),
.B(n_651),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_691),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_716),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_720),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_720),
.Y(n_784)
);

BUFx2_ASAP7_75t_R g785 ( 
.A(n_719),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_710),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_724),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_724),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_741),
.B(n_677),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_714),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_717),
.B(n_259),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_SL g792 ( 
.A1(n_715),
.A2(n_173),
.B1(n_175),
.B2(n_195),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_710),
.B(n_245),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_721),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_SL g795 ( 
.A1(n_728),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_706),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_721),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_702),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_730),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_697),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_730),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_699),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_768),
.Y(n_803)
);

OA21x2_ASAP7_75t_L g804 ( 
.A1(n_790),
.A2(n_726),
.B(n_729),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_771),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_769),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_790),
.A2(n_738),
.B(n_731),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_748),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_746),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_748),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_768),
.B(n_742),
.Y(n_811)
);

BUFx8_ASAP7_75t_L g812 ( 
.A(n_743),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_759),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_765),
.B(n_736),
.Y(n_814)
);

OAI21x1_ASAP7_75t_L g815 ( 
.A1(n_759),
.A2(n_725),
.B(n_735),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_742),
.B(n_702),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_770),
.B(n_733),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_771),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_797),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_749),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_754),
.B(n_709),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_797),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_755),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_779),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_798),
.B(n_205),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_775),
.A2(n_206),
.B(n_207),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_743),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_765),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_779),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_766),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_794),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_758),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_776),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_758),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_789),
.B(n_209),
.Y(n_836)
);

CKINVDCx8_ASAP7_75t_R g837 ( 
.A(n_764),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_798),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_762),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_789),
.B(n_244),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_766),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_762),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_780),
.B(n_210),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_775),
.A2(n_211),
.B(n_212),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_781),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_756),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_783),
.Y(n_847)
);

OAI21x1_ASAP7_75t_L g848 ( 
.A1(n_772),
.A2(n_219),
.B(n_220),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_802),
.Y(n_849)
);

AO21x2_ASAP7_75t_L g850 ( 
.A1(n_787),
.A2(n_221),
.B(n_222),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_825),
.B(n_810),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_825),
.B(n_802),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_846),
.A2(n_761),
.B(n_792),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_834),
.B(n_787),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_818),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_833),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_833),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_835),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_825),
.B(n_788),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_805),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_835),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_846),
.A2(n_786),
.B1(n_793),
.B2(n_799),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_837),
.A2(n_801),
.B1(n_796),
.B2(n_785),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_838),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_810),
.B(n_788),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_805),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_829),
.B(n_783),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_829),
.B(n_784),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_838),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_830),
.B(n_784),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_816),
.A2(n_786),
.B1(n_793),
.B2(n_817),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_810),
.B(n_774),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_836),
.A2(n_786),
.B1(n_767),
.B2(n_798),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_811),
.B(n_808),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_830),
.B(n_750),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_805),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_806),
.B(n_752),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_839),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_811),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_837),
.A2(n_796),
.B1(n_745),
.B2(n_786),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_820),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_812),
.Y(n_882)
);

AOI221xp5_ASAP7_75t_L g883 ( 
.A1(n_822),
.A2(n_795),
.B1(n_753),
.B2(n_777),
.C(n_791),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_811),
.B(n_757),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_820),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_816),
.A2(n_786),
.B1(n_791),
.B2(n_763),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_808),
.B(n_750),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_839),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_811),
.B(n_757),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_842),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_832),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_803),
.B(n_747),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_803),
.B(n_824),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_845),
.B(n_747),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_838),
.B(n_831),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_819),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_812),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_842),
.B(n_760),
.Y(n_898)
);

OAI221xp5_ASAP7_75t_SL g899 ( 
.A1(n_883),
.A2(n_843),
.B1(n_814),
.B2(n_836),
.C(n_840),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_891),
.B(n_845),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_853),
.B(n_843),
.C(n_849),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_855),
.B(n_854),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_873),
.B(n_849),
.C(n_840),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_SL g904 ( 
.A1(n_862),
.A2(n_814),
.B(n_826),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_877),
.B(n_821),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_874),
.B(n_821),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_SL g907 ( 
.A1(n_886),
.A2(n_826),
.B(n_816),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_874),
.B(n_803),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_856),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_874),
.B(n_892),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_892),
.B(n_887),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_879),
.B(n_803),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_879),
.B(n_824),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_887),
.B(n_841),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_863),
.A2(n_757),
.B1(n_816),
.B2(n_763),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_SL g916 ( 
.A1(n_871),
.A2(n_826),
.B(n_743),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_852),
.B(n_841),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_893),
.B(n_831),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_893),
.B(n_841),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_852),
.B(n_847),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_867),
.B(n_847),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_894),
.B(n_807),
.C(n_804),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_880),
.A2(n_743),
.B1(n_744),
.B2(n_826),
.Y(n_923)
);

OAI221xp5_ASAP7_75t_L g924 ( 
.A1(n_864),
.A2(n_778),
.B1(n_751),
.B2(n_800),
.C(n_773),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_867),
.B(n_847),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_868),
.B(n_823),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_860),
.B(n_838),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_L g928 ( 
.A1(n_875),
.A2(n_800),
.B1(n_819),
.B2(n_823),
.C(n_778),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_866),
.B(n_838),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_896),
.B(n_807),
.C(n_804),
.Y(n_930)
);

OAI21xp33_ASAP7_75t_L g931 ( 
.A1(n_868),
.A2(n_844),
.B(n_848),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_870),
.B(n_809),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_909),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_918),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_918),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_908),
.B(n_876),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_908),
.B(n_895),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_913),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_902),
.B(n_851),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_919),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_906),
.B(n_859),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_919),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_929),
.B(n_895),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_927),
.B(n_895),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_927),
.B(n_895),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_912),
.B(n_851),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_913),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_912),
.B(n_864),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_920),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_910),
.B(n_864),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_911),
.B(n_869),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_917),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_926),
.B(n_869),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_921),
.B(n_869),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_901),
.A2(n_889),
.B1(n_884),
.B2(n_882),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_900),
.B(n_905),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_925),
.B(n_932),
.Y(n_957)
);

BUFx2_ASAP7_75t_SL g958 ( 
.A(n_923),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_947),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_933),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_939),
.B(n_914),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_933),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_939),
.B(n_941),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_949),
.B(n_856),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_934),
.Y(n_965)
);

NAND2xp67_ASAP7_75t_SL g966 ( 
.A(n_944),
.B(n_928),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_937),
.B(n_884),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_934),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_938),
.B(n_872),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_940),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_940),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_949),
.B(n_857),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_952),
.B(n_857),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_942),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_967),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_960),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_962),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_959),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_964),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_964),
.A2(n_955),
.B(n_899),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_969),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_972),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_972),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_959),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_963),
.B(n_952),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_965),
.B(n_937),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_968),
.B(n_943),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_978),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_981),
.B(n_961),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_976),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_980),
.B(n_966),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_981),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_977),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_975),
.B(n_958),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_987),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_994),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_SL g997 ( 
.A1(n_992),
.A2(n_978),
.B(n_984),
.C(n_983),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_993),
.Y(n_998)
);

OR2x6_ASAP7_75t_L g999 ( 
.A(n_991),
.B(n_958),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_990),
.B(n_987),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_996),
.B(n_994),
.C(n_988),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_1000),
.B(n_989),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_999),
.B(n_995),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_998),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_999),
.B(n_986),
.Y(n_1005)
);

OAI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_1003),
.A2(n_988),
.B(n_979),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_1005),
.A2(n_984),
.B1(n_904),
.B2(n_997),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_1001),
.A2(n_982),
.B(n_915),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1004),
.Y(n_1009)
);

AOI211xp5_ASAP7_75t_L g1010 ( 
.A1(n_1002),
.A2(n_924),
.B(n_903),
.C(n_916),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1001),
.A2(n_986),
.B1(n_945),
.B2(n_944),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_1002),
.A2(n_985),
.B(n_973),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_SL g1013 ( 
.A(n_1010),
.B(n_1008),
.C(n_1011),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_1009),
.B(n_764),
.Y(n_1014)
);

NOR3x1_ASAP7_75t_L g1015 ( 
.A(n_1007),
.B(n_907),
.C(n_985),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_1006),
.A2(n_930),
.B1(n_850),
.B2(n_897),
.Y(n_1016)
);

OAI211xp5_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_945),
.B(n_773),
.C(n_931),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_1006),
.B(n_956),
.Y(n_1018)
);

NAND4xp75_ASAP7_75t_L g1019 ( 
.A(n_1015),
.B(n_751),
.C(n_974),
.D(n_971),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_SL g1020 ( 
.A1(n_1013),
.A2(n_970),
.B(n_743),
.Y(n_1020)
);

NAND4xp75_ASAP7_75t_L g1021 ( 
.A(n_1014),
.B(n_973),
.C(n_943),
.D(n_953),
.Y(n_1021)
);

AOI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_1018),
.A2(n_922),
.B1(n_850),
.B2(n_953),
.C(n_954),
.Y(n_1022)
);

NOR4xp25_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_950),
.C(n_951),
.D(n_935),
.Y(n_1023)
);

AOI221xp5_ASAP7_75t_L g1024 ( 
.A1(n_1016),
.A2(n_850),
.B1(n_954),
.B2(n_950),
.C(n_951),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1018),
.B(n_957),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_SL g1026 ( 
.A(n_1017),
.B(n_782),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_1019),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1026),
.A2(n_882),
.B1(n_897),
.B2(n_850),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1025),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_1021),
.A2(n_1020),
.B1(n_1024),
.B2(n_1023),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1022),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1019),
.A2(n_936),
.B1(n_947),
.B2(n_744),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1025),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_935),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_1019),
.A2(n_936),
.B1(n_744),
.B2(n_812),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1025),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_1019),
.A2(n_744),
.B1(n_812),
.B2(n_948),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1019),
.A2(n_744),
.B1(n_948),
.B2(n_957),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1025),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_1019),
.A2(n_782),
.B1(n_942),
.B2(n_828),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1025),
.Y(n_1041)
);

NOR2x1_ASAP7_75t_L g1042 ( 
.A(n_1019),
.B(n_782),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1027),
.B(n_946),
.Y(n_1043)
);

OAI221xp5_ASAP7_75t_SL g1044 ( 
.A1(n_1030),
.A2(n_828),
.B1(n_872),
.B2(n_946),
.C(n_898),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_1042),
.B(n_858),
.Y(n_1045)
);

OAI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1035),
.A2(n_838),
.B1(n_898),
.B2(n_890),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1029),
.B(n_875),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_L g1048 ( 
.A(n_1033),
.B(n_1041),
.C(n_1036),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_827),
.Y(n_1049)
);

NAND4xp75_ASAP7_75t_L g1050 ( 
.A(n_1031),
.B(n_807),
.C(n_804),
.D(n_861),
.Y(n_1050)
);

OAI211xp5_ASAP7_75t_L g1051 ( 
.A1(n_1028),
.A2(n_844),
.B(n_827),
.C(n_848),
.Y(n_1051)
);

NOR2x1_ASAP7_75t_L g1052 ( 
.A(n_1034),
.B(n_858),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_1040),
.B(n_865),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_1037),
.B(n_1032),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_1038),
.B(n_223),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_L g1056 ( 
.A(n_1042),
.B(n_861),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1027),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1027),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_1029),
.B(n_815),
.C(n_813),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1027),
.B(n_890),
.C(n_888),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1043),
.B(n_889),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_1057),
.Y(n_1062)
);

OA22x2_ASAP7_75t_L g1063 ( 
.A1(n_1058),
.A2(n_889),
.B1(n_884),
.B2(n_888),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_SL g1064 ( 
.A1(n_1045),
.A2(n_878),
.B(n_760),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1047),
.Y(n_1065)
);

AND3x1_ASAP7_75t_L g1066 ( 
.A(n_1048),
.B(n_870),
.C(n_859),
.Y(n_1066)
);

NOR2x1_ASAP7_75t_L g1067 ( 
.A(n_1056),
.B(n_224),
.Y(n_1067)
);

XOR2xp5_ASAP7_75t_L g1068 ( 
.A(n_1060),
.B(n_227),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1052),
.Y(n_1069)
);

XNOR2x1_ASAP7_75t_L g1070 ( 
.A(n_1046),
.B(n_228),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1054),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1062),
.Y(n_1072)
);

XOR2xp5_ASAP7_75t_L g1073 ( 
.A(n_1071),
.B(n_1055),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1069),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1067),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1068),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1065),
.Y(n_1077)
);

XOR2xp5_ASAP7_75t_L g1078 ( 
.A(n_1073),
.B(n_1070),
.Y(n_1078)
);

XNOR2xp5_ASAP7_75t_L g1079 ( 
.A(n_1072),
.B(n_1061),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_SL g1080 ( 
.A(n_1074),
.B(n_1044),
.C(n_1053),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1077),
.A2(n_1066),
.B1(n_1063),
.B2(n_1059),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_1078),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1079),
.A2(n_1075),
.B1(n_1076),
.B2(n_1050),
.Y(n_1083)
);

OAI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1083),
.A2(n_1081),
.B1(n_1080),
.B2(n_1049),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1082),
.A2(n_1064),
.B1(n_1049),
.B2(n_1051),
.Y(n_1085)
);

AOI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1082),
.A2(n_878),
.B1(n_813),
.B2(n_881),
.C(n_885),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_1084),
.B(n_1086),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1084),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1088),
.Y(n_1089)
);

AOI222xp33_ASAP7_75t_L g1090 ( 
.A1(n_1087),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.C1(n_235),
.C2(n_236),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1089),
.A2(n_807),
.B1(n_804),
.B2(n_813),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_R g1092 ( 
.A1(n_1091),
.A2(n_1090),
.B1(n_238),
.B2(n_239),
.C(n_242),
.Y(n_1092)
);

AOI211xp5_ASAP7_75t_L g1093 ( 
.A1(n_1092),
.A2(n_237),
.B(n_243),
.C(n_815),
.Y(n_1093)
);


endmodule