module fake_jpeg_3317_n_151 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_151);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_151;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_46),
.B(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_43),
.B1(n_48),
.B2(n_41),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_67),
.B1(n_51),
.B2(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_53),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_43),
.B1(n_48),
.B2(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_79),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_73),
.B1(n_78),
.B2(n_1),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_51),
.B1(n_55),
.B2(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_38),
.B1(n_41),
.B2(n_49),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_42),
.C(n_44),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_0),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_49),
.B(n_47),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_22),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_20),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_111),
.B1(n_89),
.B2(n_8),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_23),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_109),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_16),
.B(n_17),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_24),
.C(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_5),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_85),
.B(n_88),
.Y(n_113)
);

BUFx12f_ASAP7_75t_SL g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_19),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_27),
.B(n_28),
.Y(n_122)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_29),
.B(n_30),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_124),
.CI(n_109),
.CON(n_129),
.SN(n_129)
);

NOR2xp67_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_31),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_123),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_135),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_137),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_143),
.B1(n_126),
.B2(n_127),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_140),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

AOI31xp33_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_114),
.A3(n_120),
.B(n_129),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_128),
.A3(n_129),
.B1(n_121),
.B2(n_132),
.C1(n_116),
.C2(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_32),
.Y(n_151)
);


endmodule