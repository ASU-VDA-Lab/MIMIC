module fake_jpeg_27817_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_17),
.B(n_34),
.C(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_9),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_30),
.B1(n_16),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_56),
.B1(n_18),
.B2(n_21),
.Y(n_79)
);

OR2x4_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_20),
.Y(n_93)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_54),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_30),
.B1(n_21),
.B2(n_28),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_75),
.B1(n_18),
.B2(n_17),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_30),
.B1(n_16),
.B2(n_28),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_57),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_30),
.B1(n_16),
.B2(n_28),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_24),
.B1(n_20),
.B2(n_27),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_66),
.B(n_77),
.Y(n_111)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_31),
.Y(n_82)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_34),
.B1(n_33),
.B2(n_19),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_31),
.B(n_17),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_21),
.B1(n_29),
.B2(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_78),
.B(n_84),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_87),
.B1(n_94),
.B2(n_63),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_22),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_22),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_85),
.A2(n_108),
.B1(n_109),
.B2(n_20),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_20),
.B1(n_23),
.B2(n_3),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_18),
.B1(n_31),
.B2(n_19),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_92),
.B(n_93),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_35),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_117),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_32),
.B1(n_22),
.B2(n_35),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_32),
.B1(n_22),
.B2(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_58),
.B1(n_72),
.B2(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_102),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_64),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_69),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_22),
.B1(n_24),
.B2(n_39),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_114),
.B1(n_49),
.B2(n_47),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_11),
.B(n_12),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_27),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_67),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_47),
.B(n_20),
.C(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_24),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_118),
.A2(n_91),
.B1(n_115),
.B2(n_100),
.Y(n_173)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_121),
.Y(n_161)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_81),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_47),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_144),
.B(n_107),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_139),
.B1(n_141),
.B2(n_122),
.Y(n_177)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_136),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_78),
.A2(n_68),
.B1(n_27),
.B2(n_47),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_23),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_147),
.Y(n_158)
);

AOI22x1_ASAP7_75t_SL g145 ( 
.A1(n_80),
.A2(n_9),
.B1(n_14),
.B2(n_12),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_145),
.A2(n_85),
.B1(n_99),
.B2(n_110),
.Y(n_155)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_113),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_88),
.B(n_84),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_150),
.A2(n_152),
.B(n_153),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_156),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_111),
.B(n_86),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_114),
.B(n_99),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_155),
.A2(n_168),
.B(n_1),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_95),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_104),
.B1(n_81),
.B2(n_96),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_173),
.B1(n_179),
.B2(n_133),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_128),
.C(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_162),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_85),
.C(n_114),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_114),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_115),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_83),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_119),
.B(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_175),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_83),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_180),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_124),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_175),
.B1(n_148),
.B2(n_162),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_91),
.C(n_15),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_4),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_118),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_120),
.B(n_11),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_10),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_199),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_184),
.A2(n_202),
.B1(n_203),
.B2(n_161),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_196),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_138),
.B(n_125),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_205),
.B(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_138),
.B1(n_120),
.B2(n_127),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_194),
.A2(n_170),
.B1(n_155),
.B2(n_148),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_127),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_146),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_136),
.B1(n_134),
.B2(n_3),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_1),
.B(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_207),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_2),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_3),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_209),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_218),
.Y(n_246)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_220),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_196),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_228),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_160),
.B(n_168),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_232),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_231),
.B1(n_235),
.B2(n_203),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_178),
.B1(n_167),
.B2(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_234),
.B1(n_185),
.B2(n_200),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_184),
.A2(n_181),
.B1(n_158),
.B2(n_159),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_183),
.B1(n_198),
.B2(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_204),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_240),
.A2(n_206),
.B1(n_201),
.B2(n_209),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_189),
.C(n_195),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_243),
.C(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_189),
.C(n_195),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_187),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_260),
.Y(n_266)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_250),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_254),
.B1(n_259),
.B2(n_239),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_187),
.C(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_186),
.B1(n_185),
.B2(n_203),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_191),
.C(n_151),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_261),
.C(n_230),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_217),
.A2(n_203),
.B1(n_186),
.B2(n_205),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_258),
.A2(n_217),
.B1(n_225),
.B2(n_223),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_203),
.B1(n_194),
.B2(n_210),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_211),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_150),
.C(n_158),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_213),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_216),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_240),
.B(n_238),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_237),
.B(n_161),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_272),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_271),
.B(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_214),
.B1(n_228),
.B2(n_220),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_274),
.B(n_218),
.Y(n_292)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_163),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_219),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_260),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_235),
.B1(n_222),
.B2(n_214),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_278),
.A2(n_258),
.B1(n_243),
.B2(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_280),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_241),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_287),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_267),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_266),
.B1(n_163),
.B2(n_7),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_247),
.B1(n_252),
.B2(n_261),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_293),
.B1(n_4),
.B2(n_5),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_236),
.C(n_210),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_280),
.C(n_279),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_271),
.B(n_273),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_267),
.B1(n_268),
.B2(n_266),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_265),
.A2(n_163),
.B1(n_5),
.B2(n_7),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_275),
.B(n_264),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_291),
.B(n_283),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_281),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_298),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_283),
.B(n_281),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_4),
.C(n_5),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_304),
.C(n_293),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_7),
.C(n_286),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_7),
.B1(n_288),
.B2(n_289),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_312),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_304),
.B(n_295),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_313),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_305),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_316),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_297),
.C(n_301),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_321),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_322),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_315),
.B(n_317),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_314),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_326),
.B(n_313),
.CI(n_324),
.CON(n_327),
.SN(n_327)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_327),
.Y(n_328)
);


endmodule