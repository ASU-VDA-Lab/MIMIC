module fake_ibex_196_n_784 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_784);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_784;

wire n_599;
wire n_778;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_191;
wire n_593;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_738;
wire n_475;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_698;
wire n_187;
wire n_667;
wire n_682;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_673;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_689;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_262;
wire n_299;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_772;
wire n_768;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_605;
wire n_539;
wire n_179;
wire n_392;
wire n_354;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_164;
wire n_616;
wire n_782;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g155 ( 
.A(n_32),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_58),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_48),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_47),
.Y(n_162)
);

NOR2xp67_ASAP7_75t_L g163 ( 
.A(n_33),
.B(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_93),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_45),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_108),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_26),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_90),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVxp33_ASAP7_75t_SL g179 ( 
.A(n_50),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_36),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_64),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_78),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_46),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_4),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_114),
.Y(n_190)
);

BUFx2_ASAP7_75t_SL g191 ( 
.A(n_106),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_23),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_66),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_135),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_41),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_55),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_77),
.Y(n_199)
);

BUFx2_ASAP7_75t_SL g200 ( 
.A(n_23),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_20),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_43),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_129),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_L g206 ( 
.A(n_91),
.B(n_39),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_16),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_56),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_94),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_35),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_131),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_102),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_7),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_59),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_12),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_3),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_44),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_85),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_52),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_137),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_12),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_25),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_120),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_148),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_51),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_60),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_81),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_67),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_53),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_34),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_18),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_116),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_22),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_92),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_89),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_79),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_6),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_95),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_54),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_142),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_68),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_111),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_29),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_110),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_16),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_72),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_9),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_118),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_99),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_180),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_0),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_174),
.A2(n_73),
.B(n_153),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_37),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g267 ( 
.A1(n_174),
.A2(n_71),
.B(n_152),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_178),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_180),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_155),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_180),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_0),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_155),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_157),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_177),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_195),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_159),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_177),
.A2(n_187),
.B1(n_229),
.B2(n_182),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_172),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_160),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_182),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_195),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_195),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_158),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_195),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_161),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_201),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_165),
.Y(n_295)
);

AND2x4_ASAP7_75t_L g296 ( 
.A(n_183),
.B(n_2),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_197),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_197),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_169),
.B(n_4),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_197),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_5),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_187),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_167),
.B(n_175),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_9),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_197),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_170),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_189),
.B(n_10),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_244),
.B(n_11),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_192),
.B(n_13),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_208),
.B(n_13),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_173),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_220),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_176),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_220),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_181),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_185),
.A2(n_87),
.B(n_151),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_229),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_186),
.Y(n_320)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_188),
.B(n_38),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_220),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_193),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_194),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_235),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_198),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_220),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_207),
.B(n_14),
.Y(n_328)
);

CKINVDCx6p67_ASAP7_75t_R g329 ( 
.A(n_191),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_202),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_203),
.A2(n_88),
.B(n_149),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_204),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_228),
.B(n_237),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_269),
.B(n_258),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_296),
.Y(n_336)
);

AO21x2_ASAP7_75t_L g337 ( 
.A1(n_318),
.A2(n_211),
.B(n_210),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_269),
.B(n_216),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_275),
.B(n_215),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_217),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

OR2x6_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_200),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_266),
.B(n_261),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_263),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_263),
.Y(n_347)
);

NAND3xp33_ASAP7_75t_L g348 ( 
.A(n_264),
.B(n_243),
.C(n_226),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_263),
.Y(n_349)
);

AO22x1_ASAP7_75t_L g350 ( 
.A1(n_285),
.A2(n_254),
.B1(n_251),
.B2(n_179),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_321),
.B(n_219),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_321),
.A2(n_246),
.B1(n_240),
.B2(n_250),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_294),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_305),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_312),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_313),
.B(n_162),
.Y(n_356)
);

AND3x2_ASAP7_75t_L g357 ( 
.A(n_301),
.B(n_156),
.C(n_209),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_315),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_L g359 ( 
.A(n_266),
.B(n_166),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_306),
.Y(n_360)
);

CKINVDCx6p67_ASAP7_75t_R g361 ( 
.A(n_290),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_272),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_276),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_266),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_264),
.B(n_253),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_266),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_276),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_168),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_321),
.B(n_222),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_276),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_290),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_276),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_323),
.B(n_223),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g374 ( 
.A(n_301),
.B(n_310),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_332),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_273),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_280),
.Y(n_378)
);

CKINVDCx11_ASAP7_75t_R g379 ( 
.A(n_325),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_310),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_273),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_281),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_268),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_285),
.B(n_256),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_257),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_270),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_270),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_233),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_271),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_284),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_332),
.B(n_234),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_283),
.B(n_329),
.Y(n_392)
);

NAND3xp33_ASAP7_75t_L g393 ( 
.A(n_277),
.B(n_259),
.C(n_241),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_281),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_283),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_274),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_309),
.B(n_235),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_288),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_279),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_288),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_295),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_279),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_319),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_273),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_282),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_266),
.B(n_171),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_288),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_329),
.B(n_247),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_299),
.B(n_252),
.C(n_221),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_273),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_292),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_308),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_317),
.B(n_184),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_286),
.Y(n_415)
);

INVx5_ASAP7_75t_L g416 ( 
.A(n_298),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_319),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_288),
.Y(n_418)
);

OAI22xp33_ASAP7_75t_L g419 ( 
.A1(n_355),
.A2(n_287),
.B1(n_303),
.B2(n_240),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_317),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_320),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_353),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_339),
.B(n_333),
.Y(n_423)
);

NOR3xp33_ASAP7_75t_L g424 ( 
.A(n_352),
.B(n_397),
.C(n_392),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_351),
.A2(n_303),
.B1(n_287),
.B2(n_369),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_395),
.A2(n_246),
.B1(n_250),
.B2(n_311),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_344),
.A2(n_267),
.B(n_265),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_354),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_341),
.B(n_324),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_385),
.B(n_326),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_334),
.B(n_278),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_348),
.B(n_369),
.C(n_351),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_381),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_365),
.B(n_286),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_361),
.B(n_278),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_364),
.B(n_190),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_402),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_374),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_368),
.B(n_293),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_366),
.B(n_196),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_374),
.A2(n_302),
.B1(n_225),
.B2(n_199),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_380),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_340),
.B(n_164),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_371),
.B(n_393),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_343),
.B(n_17),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_374),
.B(n_265),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_205),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_408),
.B(n_377),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_338),
.B(n_212),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_384),
.A2(n_249),
.B1(n_214),
.B2(n_218),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_358),
.B(n_227),
.Y(n_455)
);

O2A1O1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_335),
.A2(n_267),
.B(n_265),
.C(n_163),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_408),
.B(n_230),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_365),
.B(n_231),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_336),
.B(n_232),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_345),
.A2(n_267),
.B1(n_265),
.B2(n_242),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_388),
.A2(n_331),
.B(n_206),
.C(n_238),
.Y(n_462)
);

NAND2x1_ASAP7_75t_L g463 ( 
.A(n_345),
.B(n_267),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_359),
.B(n_298),
.C(n_255),
.Y(n_464)
);

BUFx8_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_360),
.B(n_255),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_343),
.B(n_331),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_373),
.A2(n_327),
.B1(n_316),
.B2(n_314),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_410),
.Y(n_469)
);

AND2x4_ASAP7_75t_SL g470 ( 
.A(n_378),
.B(n_395),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_405),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_409),
.B(n_298),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_350),
.B(n_17),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_401),
.B(n_289),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_411),
.A2(n_327),
.B1(n_316),
.B2(n_314),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_415),
.B(n_327),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_413),
.Y(n_478)
);

O2A1O1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_391),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_357),
.B(n_289),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_383),
.Y(n_481)
);

OAI221xp5_ASAP7_75t_L g482 ( 
.A1(n_386),
.A2(n_307),
.B1(n_300),
.B2(n_297),
.C(n_291),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_357),
.B(n_289),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_403),
.B(n_40),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_396),
.B(n_389),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_42),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_406),
.B(n_337),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_337),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_423),
.B(n_21),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_437),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_456),
.A2(n_427),
.B(n_461),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_22),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_433),
.B(n_24),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_463),
.A2(n_342),
.B(n_346),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_425),
.A2(n_342),
.B1(n_349),
.B2(n_347),
.Y(n_497)
);

O2A1O1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_419),
.A2(n_418),
.B(n_400),
.C(n_398),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_438),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_24),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_434),
.B(n_25),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_458),
.B(n_445),
.Y(n_502)
);

AO32x1_ASAP7_75t_L g503 ( 
.A1(n_475),
.A2(n_382),
.A3(n_362),
.B1(n_363),
.B2(n_367),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_477),
.B(n_27),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_424),
.A2(n_291),
.B1(n_297),
.B2(n_300),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_447),
.B(n_27),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_441),
.B(n_297),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_421),
.B(n_28),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_481),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_29),
.Y(n_510)
);

BUFx12f_ASAP7_75t_L g511 ( 
.A(n_465),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_454),
.B(n_30),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_444),
.B(n_416),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_435),
.A2(n_300),
.B(n_307),
.C(n_372),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_476),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_R g516 ( 
.A(n_465),
.B(n_31),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_420),
.B(n_32),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_426),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_448),
.B(n_307),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_470),
.Y(n_520)
);

INVx6_ASAP7_75t_L g521 ( 
.A(n_473),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_476),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_455),
.B(n_300),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_476),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_480),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_457),
.B(n_57),
.Y(n_527)
);

A2O1A1Ixp33_ASAP7_75t_L g528 ( 
.A1(n_442),
.A2(n_407),
.B(n_394),
.C(n_370),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_439),
.A2(n_370),
.B(n_62),
.Y(n_529)
);

AO32x1_ASAP7_75t_L g530 ( 
.A1(n_475),
.A2(n_61),
.A3(n_63),
.B1(n_65),
.B2(n_69),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_443),
.A2(n_70),
.B(n_76),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_451),
.B(n_80),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_486),
.A2(n_82),
.B(n_83),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_467),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_483),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_485),
.B(n_96),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_428),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_464),
.A2(n_97),
.B(n_98),
.Y(n_538)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_100),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_L g540 ( 
.A1(n_479),
.A2(n_101),
.B(n_104),
.C(n_105),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_431),
.B(n_154),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_440),
.B(n_107),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_471),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_478),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_429),
.Y(n_545)
);

NOR3xp33_ASAP7_75t_L g546 ( 
.A(n_460),
.B(n_125),
.C(n_127),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_450),
.B(n_139),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_453),
.A2(n_140),
.B(n_144),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_469),
.B(n_472),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_466),
.B(n_474),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_499),
.A2(n_468),
.B1(n_482),
.B2(n_518),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_511),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_491),
.B(n_544),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_521),
.B(n_512),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_505),
.B(n_540),
.C(n_546),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_494),
.B(n_490),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_525),
.Y(n_559)
);

AOI31xp67_ASAP7_75t_L g560 ( 
.A1(n_532),
.A2(n_542),
.A3(n_541),
.B(n_523),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_508),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_519),
.A2(n_501),
.B1(n_534),
.B2(n_504),
.Y(n_562)
);

O2A1O1Ixp5_ASAP7_75t_L g563 ( 
.A1(n_527),
.A2(n_513),
.B(n_500),
.C(n_529),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_521),
.B(n_509),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_493),
.B(n_510),
.Y(n_565)
);

BUFx8_ASAP7_75t_L g566 ( 
.A(n_506),
.Y(n_566)
);

CKINVDCx8_ASAP7_75t_R g567 ( 
.A(n_506),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_498),
.B(n_517),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_522),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_526),
.B(n_535),
.Y(n_570)
);

OAI21x1_ASAP7_75t_SL g571 ( 
.A1(n_538),
.A2(n_539),
.B(n_536),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_519),
.B(n_516),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_537),
.B(n_547),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_524),
.Y(n_574)
);

AO31x2_ASAP7_75t_L g575 ( 
.A1(n_548),
.A2(n_531),
.A3(n_549),
.B(n_533),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_497),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_503),
.A2(n_550),
.B(n_545),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_551),
.A2(n_507),
.B(n_503),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_507),
.B(n_530),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_495),
.Y(n_581)
);

AO31x2_ASAP7_75t_L g582 ( 
.A1(n_514),
.A2(n_488),
.A3(n_462),
.B(n_489),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_534),
.B(n_495),
.Y(n_583)
);

AOI221x1_ASAP7_75t_L g584 ( 
.A1(n_492),
.A2(n_462),
.B1(n_546),
.B2(n_427),
.C(n_514),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_499),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_490),
.A2(n_352),
.B1(n_369),
.B2(n_351),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_534),
.B(n_495),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_490),
.A2(n_352),
.B1(n_369),
.B2(n_351),
.Y(n_588)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_498),
.A2(n_490),
.B(n_452),
.C(n_432),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_499),
.B(n_392),
.Y(n_591)
);

AO31x2_ASAP7_75t_L g592 ( 
.A1(n_514),
.A2(n_488),
.A3(n_462),
.B(n_489),
.Y(n_592)
);

BUFx2_ASAP7_75t_SL g593 ( 
.A(n_515),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_543),
.Y(n_594)
);

A2O1A1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_498),
.A2(n_490),
.B(n_452),
.C(n_432),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_490),
.A2(n_352),
.B1(n_369),
.B2(n_351),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_495),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_511),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_543),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_499),
.B(n_392),
.Y(n_600)
);

A2O1A1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_498),
.A2(n_490),
.B(n_452),
.C(n_432),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_495),
.B(n_422),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_543),
.Y(n_603)
);

AO21x2_ASAP7_75t_L g604 ( 
.A1(n_492),
.A2(n_427),
.B(n_528),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_511),
.Y(n_605)
);

BUFx6f_ASAP7_75t_SL g606 ( 
.A(n_511),
.Y(n_606)
);

AOI21xp33_ASAP7_75t_L g607 ( 
.A1(n_502),
.A2(n_417),
.B(n_403),
.Y(n_607)
);

AO31x2_ASAP7_75t_L g608 ( 
.A1(n_514),
.A2(n_488),
.A3(n_462),
.B(n_489),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_491),
.B(n_423),
.Y(n_609)
);

AO31x2_ASAP7_75t_L g610 ( 
.A1(n_514),
.A2(n_488),
.A3(n_462),
.B(n_489),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_518),
.A2(n_424),
.B1(n_352),
.B2(n_419),
.Y(n_611)
);

CKINVDCx8_ASAP7_75t_R g612 ( 
.A(n_520),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_511),
.B(n_371),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_499),
.A2(n_352),
.B1(n_319),
.B2(n_325),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_496),
.A2(n_449),
.B(n_427),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_534),
.A2(n_369),
.B1(n_351),
.B2(n_424),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_499),
.B(n_355),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_491),
.B(n_423),
.Y(n_618)
);

AND2x2_ASAP7_75t_SL g619 ( 
.A(n_534),
.B(n_283),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_612),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_569),
.Y(n_621)
);

BUFx8_ASAP7_75t_L g622 ( 
.A(n_606),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_576),
.B(n_561),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_569),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_589),
.A2(n_595),
.B(n_601),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_553),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_585),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_591),
.B(n_600),
.Y(n_628)
);

OA21x2_ASAP7_75t_L g629 ( 
.A1(n_579),
.A2(n_584),
.B(n_578),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_594),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_617),
.B(n_611),
.Y(n_631)
);

NOR2x1_ASAP7_75t_R g632 ( 
.A(n_598),
.B(n_605),
.Y(n_632)
);

AO21x1_ASAP7_75t_L g633 ( 
.A1(n_562),
.A2(n_568),
.B(n_557),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_619),
.A2(n_616),
.B1(n_555),
.B2(n_565),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_614),
.B(n_618),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_563),
.A2(n_556),
.B(n_571),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_599),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_554),
.A2(n_603),
.B(n_609),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_559),
.Y(n_639)
);

OA21x2_ASAP7_75t_L g640 ( 
.A1(n_580),
.A2(n_604),
.B(n_560),
.Y(n_640)
);

OAI21x1_ASAP7_75t_SL g641 ( 
.A1(n_570),
.A2(n_574),
.B(n_573),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_590),
.B(n_597),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_569),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_SL g644 ( 
.A1(n_552),
.A2(n_564),
.B(n_572),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_583),
.Y(n_645)
);

OAI21x1_ASAP7_75t_SL g646 ( 
.A1(n_581),
.A2(n_567),
.B(n_566),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_593),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_583),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_587),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_587),
.B(n_607),
.Y(n_650)
);

OA21x2_ASAP7_75t_L g651 ( 
.A1(n_582),
.A2(n_592),
.B(n_610),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_558),
.B(n_613),
.Y(n_652)
);

OA21x2_ASAP7_75t_L g653 ( 
.A1(n_582),
.A2(n_608),
.B(n_575),
.Y(n_653)
);

AO21x2_ASAP7_75t_L g654 ( 
.A1(n_608),
.A2(n_579),
.B(n_578),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_602),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_608),
.B(n_617),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_612),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_585),
.Y(n_658)
);

AO31x2_ASAP7_75t_L g659 ( 
.A1(n_584),
.A2(n_577),
.A3(n_579),
.B(n_615),
.Y(n_659)
);

AO31x2_ASAP7_75t_L g660 ( 
.A1(n_584),
.A2(n_577),
.A3(n_579),
.B(n_615),
.Y(n_660)
);

NAND4xp25_ASAP7_75t_L g661 ( 
.A(n_611),
.B(n_424),
.C(n_614),
.D(n_303),
.Y(n_661)
);

OAI21xp33_ASAP7_75t_SL g662 ( 
.A1(n_579),
.A2(n_321),
.B(n_351),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_576),
.B(n_561),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_586),
.A2(n_588),
.B1(n_596),
.B2(n_424),
.Y(n_664)
);

AO22x1_ASAP7_75t_L g665 ( 
.A1(n_566),
.A2(n_465),
.B1(n_319),
.B2(n_417),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_585),
.B(n_590),
.Y(n_666)
);

INVx8_ASAP7_75t_L g667 ( 
.A(n_606),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_656),
.B(n_631),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_662),
.A2(n_628),
.B(n_635),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_630),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_661),
.A2(n_628),
.B1(n_664),
.B2(n_634),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_634),
.B(n_623),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_627),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_637),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_623),
.B(n_663),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_666),
.B(n_638),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_641),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_639),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_643),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_625),
.B(n_651),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_635),
.B(n_661),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_633),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_659),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_658),
.B(n_642),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_621),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_640),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_652),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_651),
.B(n_653),
.Y(n_688)
);

BUFx8_ASAP7_75t_L g689 ( 
.A(n_622),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_660),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_653),
.B(n_650),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_654),
.B(n_645),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_654),
.B(n_648),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_646),
.B(n_624),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_647),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_691),
.B(n_680),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_691),
.B(n_629),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_681),
.B(n_626),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_668),
.B(n_629),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_677),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_692),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_677),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_693),
.Y(n_703)
);

OAI21xp33_ASAP7_75t_L g704 ( 
.A1(n_671),
.A2(n_644),
.B(n_655),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_685),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_669),
.A2(n_649),
.B1(n_636),
.B2(n_652),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_695),
.Y(n_707)
);

NOR2x1_ASAP7_75t_R g708 ( 
.A(n_689),
.B(n_626),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_688),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_675),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_676),
.B(n_665),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_686),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_709),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_696),
.B(n_683),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_705),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_712),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_696),
.B(n_683),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_696),
.B(n_690),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_710),
.B(n_672),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_700),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_700),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_700),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_700),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_699),
.B(n_697),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_710),
.B(n_672),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_713),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_724),
.B(n_701),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_724),
.B(n_707),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_716),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_714),
.B(n_697),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_720),
.A2(n_711),
.B1(n_706),
.B2(n_702),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_719),
.B(n_707),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_717),
.B(n_718),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_719),
.B(n_725),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_725),
.B(n_703),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_720),
.B(n_711),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_733),
.B(n_718),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_733),
.B(n_730),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_729),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_727),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_728),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_734),
.B(n_715),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_726),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_727),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_732),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_729),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_737),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_739),
.B(n_720),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_742),
.A2(n_736),
.B(n_731),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_739),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_746),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

AOI21xp33_ASAP7_75t_SL g753 ( 
.A1(n_745),
.A2(n_667),
.B(n_736),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_743),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_738),
.A2(n_720),
.B1(n_723),
.B2(n_722),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_749),
.A2(n_753),
.B(n_748),
.C(n_755),
.Y(n_756)
);

AOI221xp5_ASAP7_75t_L g757 ( 
.A1(n_747),
.A2(n_741),
.B1(n_740),
.B2(n_744),
.C(n_738),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_SL g758 ( 
.A1(n_748),
.A2(n_667),
.B(n_721),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_752),
.B(n_708),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_756),
.A2(n_708),
.B(n_667),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_L g761 ( 
.A1(n_757),
.A2(n_754),
.B1(n_673),
.B2(n_704),
.C(n_735),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_SL g762 ( 
.A(n_758),
.B(n_620),
.C(n_657),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_760),
.B(n_759),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_762),
.B(n_632),
.C(n_698),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_763),
.B(n_761),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_764),
.B(n_737),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_765),
.B(n_751),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_766),
.B(n_657),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_768),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_767),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_769),
.B(n_622),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_770),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_771),
.B(n_689),
.C(n_687),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_772),
.Y(n_774)
);

AOI22x1_ASAP7_75t_L g775 ( 
.A1(n_774),
.A2(n_684),
.B1(n_722),
.B2(n_723),
.Y(n_775)
);

NOR3xp33_ASAP7_75t_L g776 ( 
.A(n_773),
.B(n_704),
.C(n_670),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_774),
.B(n_750),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_774),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_694),
.B1(n_682),
.B2(n_721),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_777),
.B(n_694),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_779),
.A2(n_775),
.B(n_776),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_780),
.B(n_694),
.C(n_674),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_781),
.B(n_679),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_783),
.A2(n_782),
.B(n_678),
.Y(n_784)
);


endmodule