module fake_jpeg_974_n_17 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_17);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_17;

wire n_13;
wire n_14;
wire n_16;
wire n_15;

INVx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_7),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_12),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_16)
);

AOI322xp5_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_14),
.A3(n_15),
.B1(n_9),
.B2(n_10),
.C1(n_5),
.C2(n_8),
.Y(n_17)
);


endmodule