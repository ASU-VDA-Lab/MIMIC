module fake_jpeg_8054_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_64),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_21),
.B1(n_25),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_62),
.B1(n_19),
.B2(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_19),
.C(n_33),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_32),
.B1(n_20),
.B2(n_17),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_24),
.B1(n_27),
.B2(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_40),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_32),
.B1(n_25),
.B2(n_33),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_36),
.B1(n_41),
.B2(n_44),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_79),
.B1(n_94),
.B2(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_80),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_41),
.B1(n_43),
.B2(n_42),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_88),
.Y(n_112)
);

BUFx4f_ASAP7_75t_SL g85 ( 
.A(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_24),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_38),
.B1(n_40),
.B2(n_44),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_97),
.B1(n_50),
.B2(n_49),
.Y(n_106)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_100),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_66),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_103),
.C(n_119),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_64),
.C(n_62),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_44),
.B1(n_59),
.B2(n_51),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_106),
.B1(n_116),
.B2(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_44),
.B1(n_53),
.B2(n_43),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_37),
.B1(n_39),
.B2(n_49),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_48),
.C(n_39),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_48),
.Y(n_122)
);

AO21x2_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_90),
.B(n_89),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_39),
.C(n_47),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_127),
.B(n_129),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_42),
.B1(n_43),
.B2(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_149),
.B1(n_150),
.B2(n_154),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_134),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_132),
.A2(n_137),
.B1(n_143),
.B2(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_138),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_144),
.B(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_110),
.B1(n_124),
.B2(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_83),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_53),
.B1(n_86),
.B2(n_42),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_86),
.B1(n_91),
.B2(n_84),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_119),
.A2(n_97),
.B1(n_82),
.B2(n_38),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_82),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_153),
.A2(n_31),
.B1(n_18),
.B2(n_34),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_123),
.A2(n_47),
.B1(n_46),
.B2(n_38),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_123),
.B1(n_103),
.B2(n_101),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_164),
.B1(n_173),
.B2(n_152),
.Y(n_201)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_163),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_101),
.B(n_26),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_168),
.B(n_169),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_40),
.C(n_38),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_126),
.B1(n_104),
.B2(n_120),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_80),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_38),
.C(n_40),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_35),
.B(n_26),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_16),
.B(n_12),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_113),
.B1(n_40),
.B2(n_46),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_181),
.B1(n_182),
.B2(n_135),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_120),
.B1(n_113),
.B2(n_109),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_35),
.B1(n_23),
.B2(n_28),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_179),
.B(n_23),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_148),
.B(n_133),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_100),
.C(n_98),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_47),
.C(n_109),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_18),
.B(n_34),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_180),
.B(n_0),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_47),
.B1(n_46),
.B2(n_28),
.Y(n_181)
);

OAI22x1_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_28),
.B1(n_23),
.B2(n_46),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_150),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_129),
.Y(n_187)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_191),
.Y(n_235)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_200),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_193),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_149),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_206),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_170),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_205),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_179),
.A2(n_134),
.B(n_137),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_161),
.B(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_181),
.B1(n_158),
.B2(n_159),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_180),
.B1(n_182),
.B2(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_34),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_34),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_46),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_109),
.B1(n_47),
.B2(n_10),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_160),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_210),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_164),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_0),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_212),
.A2(n_10),
.B(n_16),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_226),
.B1(n_236),
.B2(n_189),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_218),
.A2(n_234),
.B(n_198),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_159),
.B1(n_183),
.B2(n_2),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_8),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_211),
.C(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_9),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_9),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_233),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_9),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_186),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_0),
.Y(n_261)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_228),
.C(n_232),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_253),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_223),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_258),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_203),
.B1(n_191),
.B2(n_205),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_261),
.B(n_214),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_246),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_195),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_225),
.B1(n_227),
.B2(n_217),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_227),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_255),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_208),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_259),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_202),
.B1(n_208),
.B2(n_185),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_199),
.CI(n_196),
.CON(n_258),
.SN(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_213),
.B(n_193),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_196),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_214),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_268),
.C(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_238),
.C(n_225),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_230),
.C(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_279),
.C(n_250),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_10),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_240),
.B1(n_245),
.B2(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_241),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_272),
.B1(n_275),
.B2(n_277),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_267),
.A2(n_245),
.B(n_244),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_276),
.B(n_258),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_263),
.A2(n_245),
.B1(n_248),
.B2(n_258),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_243),
.B1(n_279),
.B2(n_247),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_250),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_299),
.B(n_12),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_303),
.B(n_304),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_275),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_273),
.C(n_12),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_14),
.B1(n_15),
.B2(n_3),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_273),
.B(n_11),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_287),
.B(n_293),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_311),
.B(n_317),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_6),
.B(n_7),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_301),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_295),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_298),
.B1(n_296),
.B2(n_15),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g322 ( 
.A1(n_314),
.A2(n_296),
.B(n_15),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_323),
.B(n_310),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_3),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

NAND2x1_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_311),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_324),
.A2(n_3),
.B(n_4),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_328),
.B(n_321),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_325),
.Y(n_332)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_332),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_330),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_321),
.CI(n_4),
.CON(n_336),
.SN(n_336)
);


endmodule