module fake_jpeg_13578_n_418 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_418);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_418;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_57),
.Y(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_59),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_16),
.C(n_15),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_60),
.A2(n_107),
.B(n_2),
.C(n_9),
.Y(n_159)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_63),
.Y(n_168)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_12),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_65),
.B(n_71),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_12),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_68),
.B(n_94),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_73),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_12),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_79),
.Y(n_147)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_45),
.Y(n_79)
);

INVx11_ASAP7_75t_SL g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_81),
.Y(n_177)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_82),
.B(n_83),
.Y(n_175)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_11),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_100),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_92),
.Y(n_145)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_93),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_10),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_97),
.B(n_99),
.Y(n_148)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_10),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_101),
.B(n_104),
.Y(n_151)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_103),
.Y(n_157)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_0),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_106),
.B1(n_112),
.B2(n_28),
.Y(n_119)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_26),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_26),
.B(n_1),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_153)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_58),
.A2(n_41),
.B1(n_35),
.B2(n_28),
.Y(n_120)
);

OAI22x1_ASAP7_75t_L g206 ( 
.A1(n_120),
.A2(n_123),
.B1(n_133),
.B2(n_141),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_35),
.B1(n_41),
.B2(n_53),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_121),
.A2(n_125),
.B1(n_128),
.B2(n_130),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_58),
.A2(n_35),
.B1(n_52),
.B2(n_50),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_60),
.A2(n_53),
.B1(n_50),
.B2(n_31),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_62),
.A2(n_53),
.B1(n_50),
.B2(n_31),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_31),
.B1(n_27),
.B2(n_52),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_129),
.A2(n_160),
.A3(n_177),
.B1(n_158),
.B2(n_170),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_27),
.B1(n_47),
.B2(n_34),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_63),
.A2(n_27),
.B1(n_32),
.B2(n_38),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_131),
.A2(n_139),
.B1(n_149),
.B2(n_154),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_25),
.B1(n_47),
.B2(n_34),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_100),
.A2(n_33),
.B1(n_38),
.B2(n_32),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_138),
.A2(n_160),
.B1(n_171),
.B2(n_134),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_66),
.A2(n_33),
.B1(n_36),
.B2(n_17),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_70),
.A2(n_36),
.B1(n_44),
.B2(n_39),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_87),
.A2(n_44),
.B1(n_39),
.B2(n_49),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_146),
.A2(n_156),
.B1(n_165),
.B2(n_166),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_67),
.A2(n_49),
.B1(n_6),
.B2(n_7),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_72),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_87),
.A2(n_39),
.B1(n_6),
.B2(n_9),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_89),
.A2(n_9),
.B1(n_39),
.B2(n_96),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_74),
.A2(n_86),
.B1(n_76),
.B2(n_98),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_172),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_61),
.B1(n_78),
.B2(n_93),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_91),
.A2(n_106),
.B1(n_112),
.B2(n_80),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_91),
.A2(n_112),
.B1(n_92),
.B2(n_85),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_92),
.A2(n_59),
.B1(n_82),
.B2(n_81),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_100),
.A2(n_60),
.B1(n_88),
.B2(n_89),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_75),
.A2(n_67),
.B1(n_66),
.B2(n_72),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_137),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_179),
.B(n_183),
.C(n_188),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_180),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_181),
.B(n_185),
.Y(n_253)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_182),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_137),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_184),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_132),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_186),
.B(n_190),
.Y(n_266)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_152),
.C(n_153),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_151),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_191),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_122),
.B(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_194),
.B(n_195),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_115),
.Y(n_195)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_113),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_197),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_153),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_213),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_115),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_199),
.B(n_202),
.Y(n_275)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_127),
.B(n_118),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_210),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_205),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_130),
.B(n_138),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_216),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_129),
.A2(n_155),
.B(n_163),
.C(n_118),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_208),
.A2(n_219),
.B(n_197),
.C(n_210),
.Y(n_261)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_144),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_142),
.B(n_129),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_142),
.B(n_129),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_189),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_221),
.B1(n_231),
.B2(n_213),
.Y(n_243)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_224),
.Y(n_245)
);

BUFx8_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

CKINVDCx12_ASAP7_75t_R g247 ( 
.A(n_218),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_144),
.B(n_124),
.C(n_126),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g220 ( 
.A1(n_158),
.A2(n_176),
.B1(n_169),
.B2(n_164),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_208),
.B(n_214),
.Y(n_242)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_117),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_126),
.B1(n_134),
.B2(n_135),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_117),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_227),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_136),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_229),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_135),
.B(n_136),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_143),
.B(n_150),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_233),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_143),
.A2(n_138),
.B1(n_160),
.B2(n_171),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_150),
.B(n_137),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_228),
.Y(n_267)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_116),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_192),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_181),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_246),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_SL g283 ( 
.A1(n_239),
.A2(n_242),
.B(n_248),
.C(n_257),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_249),
.B1(n_256),
.B2(n_269),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_243),
.Y(n_286)
);

AND2x6_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_232),
.Y(n_246)
);

OAI22x1_ASAP7_75t_SL g248 ( 
.A1(n_205),
.A2(n_215),
.B1(n_206),
.B2(n_178),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_214),
.A2(n_179),
.B1(n_183),
.B2(n_178),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_179),
.A2(n_183),
.B1(n_211),
.B2(n_226),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_207),
.B(n_206),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_192),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_249),
.Y(n_291)
);

AO21x1_ASAP7_75t_SL g278 ( 
.A1(n_261),
.A2(n_196),
.B(n_218),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_277),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_268),
.B(n_260),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_187),
.A2(n_191),
.B1(n_216),
.B2(n_225),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_222),
.A2(n_209),
.B1(n_184),
.B2(n_193),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_274),
.A2(n_260),
.B1(n_257),
.B2(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_180),
.B(n_203),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_278),
.A2(n_251),
.B(n_254),
.C(n_272),
.Y(n_319)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_245),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_282),
.B(n_292),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_201),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_285),
.C(n_288),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_241),
.B(n_218),
.C(n_201),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_302),
.B(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_291),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_238),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_294),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_265),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_237),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_297),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_298),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_299),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_246),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_300),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_266),
.B(n_271),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_262),
.B(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_242),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_239),
.A2(n_261),
.B1(n_258),
.B2(n_235),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_239),
.B1(n_247),
.B2(n_235),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_251),
.B(n_272),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_269),
.B1(n_255),
.B2(n_273),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_322),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_290),
.A2(n_255),
.B1(n_273),
.B2(n_263),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_321),
.B1(n_324),
.B2(n_326),
.Y(n_341)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_286),
.A2(n_273),
.B1(n_263),
.B2(n_236),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_294),
.A2(n_263),
.B1(n_251),
.B2(n_254),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_290),
.A2(n_305),
.B1(n_300),
.B2(n_281),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_279),
.B1(n_278),
.B2(n_283),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_283),
.B(n_296),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_333),
.A2(n_310),
.B(n_323),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_289),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_334),
.B(n_343),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_328),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_348),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_317),
.B(n_293),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_285),
.C(n_288),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_287),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_345),
.B(n_346),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_303),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_315),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_314),
.B(n_298),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_351),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_331),
.B(n_284),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_331),
.C(n_336),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_329),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_327),
.C(n_283),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_361),
.B(n_320),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_326),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_319),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_352),
.A2(n_311),
.B(n_283),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_338),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_349),
.A2(n_324),
.B1(n_321),
.B2(n_316),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_366),
.A2(n_341),
.B1(n_312),
.B2(n_322),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_341),
.A2(n_323),
.B1(n_327),
.B2(n_313),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_367),
.A2(n_338),
.B1(n_337),
.B2(n_333),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_357),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_376),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_374),
.Y(n_389)
);

OAI322xp33_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_334),
.A3(n_345),
.B1(n_348),
.B2(n_344),
.C1(n_346),
.C2(n_335),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_375),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_363),
.C(n_365),
.Y(n_392)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_356),
.Y(n_373)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

OAI322xp33_ASAP7_75t_L g375 ( 
.A1(n_358),
.A2(n_315),
.A3(n_342),
.B1(n_340),
.B2(n_339),
.C1(n_337),
.C2(n_319),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_320),
.C(n_330),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_361),
.C(n_362),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_381),
.Y(n_383)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_380),
.B(n_365),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_355),
.B(n_351),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_382),
.B(n_364),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_384),
.B(n_385),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_377),
.B(n_367),
.C(n_354),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_392),
.Y(n_393)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_390),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_389),
.A2(n_379),
.B(n_370),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_395),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_388),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_364),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_400),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_389),
.A2(n_379),
.B(n_374),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_399),
.A2(n_381),
.B(n_383),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_368),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_372),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_394),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_393),
.B(n_383),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_403),
.B(n_406),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_396),
.A2(n_391),
.B1(n_380),
.B2(n_373),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_405),
.A2(n_396),
.B1(n_359),
.B2(n_360),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_407),
.B(n_409),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_399),
.C(n_378),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_410),
.A2(n_404),
.B(n_366),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_404),
.C(n_402),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_408),
.C(n_410),
.Y(n_414)
);

INVxp33_ASAP7_75t_L g415 ( 
.A(n_413),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_414),
.B(n_412),
.C(n_368),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_415),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_417),
.B(n_360),
.Y(n_418)
);


endmodule