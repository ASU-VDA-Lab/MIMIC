module real_jpeg_23656_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_114;
wire n_49;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_262;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_216;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_20),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_34),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_1),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_1),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_20),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_46),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_27),
.B1(n_46),
.B2(n_66),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_20),
.B1(n_24),
.B2(n_30),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_6),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_6),
.A2(n_30),
.B1(n_54),
.B2(n_55),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_6),
.B(n_20),
.C(n_23),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_6),
.B(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_38),
.C(n_40),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_52),
.C(n_55),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_6),
.B(n_44),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_6),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_6),
.B(n_118),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_10),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_269),
.B(n_272),
.Y(n_11)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_72),
.B(n_268),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_70),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_14),
.B(n_70),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_60),
.C(n_62),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_15),
.A2(n_16),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_31),
.C(n_47),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_17),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_17),
.A2(n_81),
.B1(n_97),
.B2(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_17),
.B(n_114),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_17),
.A2(n_81),
.B1(n_113),
.B2(n_114),
.Y(n_136)
);

AOI211xp5_ASAP7_75t_L g158 ( 
.A1(n_17),
.A2(n_127),
.B(n_130),
.C(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_17),
.A2(n_81),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_17),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_17),
.A2(n_81),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_17),
.A2(n_95),
.B(n_98),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_29),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_18),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_19),
.A2(n_25),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_19),
.A2(n_25),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_19),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_20),
.A2(n_24),
.B1(n_38),
.B2(n_42),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_20),
.B(n_190),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_27),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_31),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_32)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_36),
.A2(n_37),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_40),
.B(n_201),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_47),
.A2(n_48),
.B1(n_84),
.B2(n_256),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_81),
.C(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_57),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_55),
.B(n_211),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_62),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_61),
.B(n_86),
.Y(n_114)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_70),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_70),
.B(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_71),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_88),
.B(n_267),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_74),
.B(n_77),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.C(n_83),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_113),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_83),
.B(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_84),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI31xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_248),
.A3(n_259),
.B(n_264),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_149),
.B(n_247),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_132),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_91),
.B(n_132),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_121),
.B1(n_122),
.B2(n_131),
.Y(n_91)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_111),
.B2(n_112),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_94),
.B(n_111),
.C(n_121),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_109),
.B2(n_110),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_98),
.B1(n_105),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_102),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_101),
.B(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_125),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_104),
.Y(n_212)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_115),
.B(n_120),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_157),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_113),
.A2(n_114),
.B1(n_127),
.B2(n_157),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_113),
.A2(n_114),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_162),
.C(n_177),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_114),
.A2(n_127),
.B(n_159),
.C(n_222),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_120),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_120),
.A2(n_253),
.B1(n_257),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_128),
.B(n_129),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_124),
.A2(n_127),
.B1(n_157),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_124),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_143),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_127),
.B(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_127),
.A2(n_157),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_127),
.A2(n_157),
.B1(n_199),
.B2(n_200),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_127),
.A2(n_157),
.B1(n_187),
.B2(n_228),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_128),
.A2(n_129),
.B(n_161),
.Y(n_239)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_141),
.B(n_148),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.C(n_140),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_133),
.A2(n_134),
.B1(n_138),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_136),
.B1(n_161),
.B2(n_168),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_142),
.Y(n_236)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_138),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_140),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_241),
.B(n_246),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_180),
.B(n_232),
.C(n_240),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_170),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_152),
.B(n_170),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_169),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_155),
.B(n_158),
.C(n_169),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_184),
.C(n_187),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_163),
.C(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_163),
.B1(n_177),
.B2(n_178),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_163),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_162),
.A2(n_163),
.B1(n_188),
.B2(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_163),
.B(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_172),
.A2(n_173),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_231),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_194),
.B(n_230),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_183),
.B(n_191),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_224),
.B(n_229),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_218),
.B(n_223),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_207),
.B(n_217),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_202),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_220),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_237),
.C(n_239),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_245),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_252),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.C(n_258),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_261),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_263),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);


endmodule