module fake_jpeg_28878_n_369 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_369);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_369;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx3_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_50),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_64),
.Y(n_90)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_68),
.Y(n_110)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_39),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_24),
.B1(n_45),
.B2(n_33),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_96),
.A2(n_68),
.B1(n_33),
.B2(n_26),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_31),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_106),
.Y(n_133)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_54),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_44),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_38),
.Y(n_135)
);

OR2x2_ASAP7_75t_SL g106 ( 
.A(n_51),
.B(n_32),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_56),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_116),
.A2(n_119),
.B1(n_123),
.B2(n_110),
.Y(n_164)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_71),
.B1(n_47),
.B2(n_45),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_22),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_136),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_24),
.B1(n_33),
.B2(n_45),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_126),
.A2(n_110),
.B1(n_107),
.B2(n_78),
.Y(n_160)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_135),
.Y(n_165)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_22),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_41),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_44),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_27),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_106),
.B1(n_136),
.B2(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_153),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_75),
.B1(n_102),
.B2(n_101),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_101),
.B1(n_115),
.B2(n_83),
.Y(n_171)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_88),
.A3(n_89),
.B1(n_68),
.B2(n_39),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_161),
.Y(n_174)
);

AOI22x1_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_32),
.B1(n_107),
.B2(n_78),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_75),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_131),
.B(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_27),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_38),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_173),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_179),
.B1(n_122),
.B2(n_83),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_158),
.B(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_102),
.B1(n_84),
.B2(n_80),
.Y(n_179)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_151),
.B(n_127),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_180),
.A2(n_182),
.B(n_132),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_117),
.B(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_183),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_146),
.B1(n_153),
.B2(n_149),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_200),
.B1(n_201),
.B2(n_179),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_202),
.B(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_203),
.Y(n_212)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_199),
.B1(n_173),
.B2(n_157),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_150),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_154),
.B1(n_157),
.B2(n_113),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_185),
.B1(n_174),
.B2(n_182),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_144),
.B1(n_114),
.B2(n_125),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_165),
.B(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_162),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_178),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_206),
.A2(n_210),
.B1(n_225),
.B2(n_226),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_177),
.C(n_182),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_202),
.C(n_188),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_214),
.B(n_191),
.Y(n_242)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_179),
.B1(n_171),
.B2(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_219),
.Y(n_229)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_194),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_221),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_176),
.B1(n_183),
.B2(n_184),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_223),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_162),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_158),
.B1(n_147),
.B2(n_156),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_147),
.B1(n_156),
.B2(n_159),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_222),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_212),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_201),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_210),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_34),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_239),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_216),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_199),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_32),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_240),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_191),
.C(n_189),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_246),
.C(n_211),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_197),
.C(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_262),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_237),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_252),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_218),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_214),
.B(n_209),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_214),
.B(n_209),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_255),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_213),
.B1(n_217),
.B2(n_226),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_256),
.A2(n_129),
.B1(n_114),
.B2(n_125),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_266),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_271),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_236),
.B(n_227),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_137),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_34),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_265),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_217),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_269),
.B1(n_240),
.B2(n_244),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_234),
.B(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_267),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_238),
.Y(n_269)
);

NOR2x1_ASAP7_75t_R g272 ( 
.A(n_270),
.B(n_265),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_272),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_247),
.B1(n_241),
.B2(n_238),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_274),
.A2(n_290),
.B1(n_293),
.B2(n_273),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_260),
.A2(n_247),
.B1(n_246),
.B2(n_163),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_289),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_139),
.C(n_142),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_291),
.C(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_253),
.B1(n_256),
.B2(n_264),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_46),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_142),
.B1(n_118),
.B2(n_40),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_112),
.C(n_104),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_104),
.C(n_112),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_36),
.B1(n_29),
.B2(n_46),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_261),
.B(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_271),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_297),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_286),
.B1(n_47),
.B2(n_24),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_270),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_309),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_267),
.B(n_42),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_300),
.B(n_306),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_40),
.C(n_29),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_304),
.C(n_307),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_32),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_272),
.A2(n_42),
.B(n_37),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_36),
.C(n_23),
.Y(n_307)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_21),
.C(n_20),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_19),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_283),
.B1(n_288),
.B2(n_279),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_303),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_292),
.C(n_283),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_315),
.B(n_319),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_318),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_41),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_286),
.C(n_37),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_286),
.C(n_23),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_322),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_305),
.A2(n_19),
.B(n_18),
.Y(n_321)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_321),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_0),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_334),
.Y(n_339)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_323),
.A2(n_301),
.B(n_303),
.Y(n_326)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_326),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_296),
.B1(n_307),
.B2(n_304),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_330),
.A2(n_329),
.B1(n_6),
.B2(n_7),
.Y(n_346)
);

NOR2x1_ASAP7_75t_SL g332 ( 
.A(n_319),
.B(n_295),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_332),
.A2(n_336),
.B(n_1),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_312),
.A2(n_138),
.B(n_120),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_315),
.A2(n_138),
.B(n_120),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_311),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_320),
.A2(n_91),
.B(n_2),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_324),
.C(n_311),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_340),
.Y(n_351)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_338),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_324),
.C(n_4),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_327),
.Y(n_341)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_341),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_1),
.C(n_4),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_344),
.C(n_7),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_331),
.A2(n_4),
.B(n_5),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_347),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g348 ( 
.A1(n_341),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_348),
.A2(n_339),
.B(n_12),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_355),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_8),
.C(n_9),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_345),
.C(n_347),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_356),
.B(n_360),
.Y(n_363)
);

AO21x1_ASAP7_75t_L g362 ( 
.A1(n_357),
.A2(n_358),
.B(n_354),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_350),
.A2(n_10),
.B(n_12),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_13),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_359),
.B(n_352),
.Y(n_361)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_361),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g364 ( 
.A1(n_362),
.A2(n_353),
.B(n_348),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_364),
.A2(n_363),
.B(n_360),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_365),
.B(n_14),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_368),
.A2(n_16),
.B1(n_17),
.B2(n_228),
.Y(n_369)
);


endmodule