module real_jpeg_23886_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_0),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_0),
.B(n_48),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_0),
.B(n_46),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_0),
.B(n_51),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_0),
.B(n_32),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_0),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_0),
.B(n_66),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_0),
.B(n_89),
.Y(n_258)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_2),
.B(n_46),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_66),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_2),
.B(n_48),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_2),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_2),
.B(n_32),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_89),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_4),
.B(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_4),
.B(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_4),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_32),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_4),
.B(n_51),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_4),
.B(n_48),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_32),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_6),
.B(n_51),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_6),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_6),
.B(n_48),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_6),
.B(n_46),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_6),
.B(n_66),
.Y(n_292)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_8),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_8),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_8),
.B(n_17),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_8),
.B(n_32),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_8),
.B(n_51),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_17),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_9),
.B(n_32),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_9),
.B(n_51),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_51),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_12),
.B(n_48),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_12),
.B(n_32),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_12),
.B(n_17),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_12),
.B(n_46),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_12),
.B(n_66),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_14),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_14),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_14),
.B(n_48),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_14),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_46),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_15),
.B(n_46),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_51),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_15),
.B(n_66),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_15),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_16),
.B(n_51),
.Y(n_82)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_17),
.Y(n_178)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_17),
.Y(n_223)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_152),
.CON(n_18),
.SN(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_21),
.B(n_77),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_54),
.C(n_71),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_44),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_23),
.B(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_29),
.C(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_26),
.B(n_60),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_29),
.A2(n_37),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_29),
.B(n_79),
.C(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_30),
.B(n_61),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_34),
.A2(n_36),
.B1(n_39),
.B2(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_35),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_39),
.C(n_40),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_38),
.B(n_44),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_39),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_40),
.A2(n_41),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_44),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.CI(n_50),
.CON(n_44),
.SN(n_44)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_47),
.C(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_51),
.Y(n_218)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_71),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_56),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.C(n_62),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_62),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_69),
.B1(n_75),
.B2(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_74),
.C(n_76),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_70),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_84),
.C(n_85),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_81),
.A2(n_82),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g331 ( 
.A(n_85),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.CI(n_88),
.CON(n_85),
.SN(n_85)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_87),
.C(n_88),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_90),
.B(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_104),
.C(n_108),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_91),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_100),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_92),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_94),
.B(n_100),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_97),
.B(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_104),
.B(n_108),
.Y(n_325)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_121),
.C(n_122),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_109),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_119),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_110),
.B(n_119),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_115),
.B(n_301),
.Y(n_300)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_121),
.B(n_122),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_138),
.B2(n_139),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_134),
.B2(n_135),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_327),
.C(n_328),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_317),
.C(n_318),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_303),
.C(n_304),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_280),
.C(n_281),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_248),
.C(n_249),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_228),
.C(n_229),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_188),
.C(n_200),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_173),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_161),
.B(n_168),
.C(n_173),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_163),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_169),
.B(n_171),
.C(n_172),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_181),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_174),
.B(n_182),
.C(n_183),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_187),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_199),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_192),
.A2(n_193),
.B1(n_199),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_224),
.C(n_225),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.C(n_214),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.C(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_242),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_243),
.C(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_238),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_237),
.C(n_238),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_233),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_236),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_238),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.CI(n_241),
.CON(n_238),
.SN(n_238)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_243),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.CI(n_246),
.CON(n_243),
.SN(n_243)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_264),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_253),
.C(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_259),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_260),
.C(n_263),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_255),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.CI(n_258),
.CON(n_255),
.SN(n_255)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_257),
.C(n_258),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_272),
.C(n_278),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_272),
.B1(n_278),
.B2(n_279),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_267),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_270),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_270),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_299),
.C(n_300),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_295),
.B2(n_302),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_296),
.C(n_297),
.Y(n_303)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_286),
.C(n_288),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_293),
.C(n_294),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_315),
.B2(n_316),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.C(n_315),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_321),
.C(n_326),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_324),
.B2(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);


endmodule