module fake_jpeg_590_n_125 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_16),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_41),
.B1(n_37),
.B2(n_39),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_35),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_41),
.B(n_43),
.C(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_66),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_67),
.B(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_81),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_6),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_23),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_51),
.C(n_14),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_51),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_17),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_22),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_100),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_76),
.C(n_80),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_106),
.C(n_94),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_8),
.B1(n_11),
.B2(n_15),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_7),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_105),
.A2(n_94),
.B(n_9),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_111),
.C(n_112),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_110),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_91),
.B1(n_9),
.B2(n_10),
.Y(n_109)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_102),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_106),
.C(n_101),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_119),
.B1(n_115),
.B2(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_98),
.C(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_114),
.C(n_98),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_28),
.Y(n_125)
);


endmodule