module fake_jpeg_8715_n_208 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_50),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_64),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_60),
.B1(n_62),
.B2(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_34),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_34),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_27),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_28),
.C(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_19),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_28),
.B1(n_38),
.B2(n_19),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_72),
.B(n_95),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_94),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_38),
.B1(n_30),
.B2(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_76),
.Y(n_108)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_84),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_37),
.B1(n_40),
.B2(n_45),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_81),
.B1(n_89),
.B2(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_1),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_80),
.Y(n_110)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_92),
.B1(n_61),
.B2(n_55),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_24),
.B1(n_27),
.B2(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_30),
.B1(n_23),
.B2(n_29),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_36),
.C(n_43),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_29),
.B(n_36),
.C(n_23),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_52),
.B(n_48),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_118),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_102),
.B(n_104),
.Y(n_132)
);

OR2x6_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_40),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_36),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_52),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_47),
.B1(n_37),
.B2(n_40),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_47),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_43),
.B1(n_24),
.B2(n_29),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_43),
.B1(n_36),
.B2(n_15),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_127),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_79),
.C(n_82),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_142),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_138),
.B(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_73),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_76),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_84),
.B1(n_96),
.B2(n_90),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_141),
.B1(n_111),
.B2(n_78),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_75),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_120),
.B1(n_110),
.B2(n_105),
.C(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_77),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_14),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_104),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_104),
.B1(n_115),
.B2(n_99),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_78),
.C(n_88),
.Y(n_142)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_102),
.B1(n_115),
.B2(n_113),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_149),
.B(n_3),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_130),
.Y(n_167)
);

OAI211xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_158),
.B(n_133),
.C(n_3),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_155),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_141),
.B(n_136),
.Y(n_149)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_78),
.B1(n_119),
.B2(n_100),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_131),
.B1(n_130),
.B2(n_5),
.Y(n_166)
);

NOR4xp25_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_12),
.C(n_11),
.D(n_4),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_119),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_123),
.C(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_162),
.Y(n_181)
);

XOR2x2_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_132),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_161),
.B(n_167),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_164),
.C(n_168),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_138),
.C(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_2),
.C(n_3),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_2),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_159),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_143),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_5),
.C(n_6),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_173),
.C(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_175),
.B(n_178),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_177),
.Y(n_189)
);

OAI321xp33_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_143),
.A3(n_149),
.B1(n_147),
.B2(n_145),
.C(n_144),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_179),
.A2(n_167),
.B1(n_144),
.B2(n_165),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_7),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_188),
.B1(n_180),
.B2(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_163),
.C(n_164),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_187),
.C(n_176),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_148),
.C(n_168),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_157),
.B1(n_152),
.B2(n_155),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_172),
.B(n_8),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_176),
.C(n_9),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_186),
.C(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_8),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_195),
.B(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_9),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_198),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_194),
.B(n_192),
.Y(n_202)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_202),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_204),
.B(n_9),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_205),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);


endmodule