module real_aes_3422_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_235;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_962;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_860;
wire n_781;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_936;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_947;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_639;
wire n_151;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g129 ( .A(n_0), .B(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_1), .Y(n_176) );
OA22x2_ASAP7_75t_L g117 ( .A1(n_2), .A2(n_118), .B1(n_119), .B2(n_120), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_2), .Y(n_118) );
O2A1O1Ixp33_ASAP7_75t_SL g202 ( .A1(n_3), .A2(n_171), .B(n_203), .C(n_204), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g142 ( .A1(n_4), .A2(n_84), .B1(n_137), .B2(n_143), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_5), .A2(n_32), .B1(n_594), .B2(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
INVx1_ASAP7_75t_L g543 ( .A(n_6), .Y(n_543) );
INVx1_ASAP7_75t_L g936 ( .A(n_6), .Y(n_936) );
NAND3xp33_ASAP7_75t_SL g961 ( .A(n_6), .B(n_962), .C(n_963), .Y(n_961) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_7), .Y(n_951) );
OAI22x1_ASAP7_75t_R g524 ( .A1(n_8), .A2(n_83), .B1(n_525), .B2(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g526 ( .A(n_8), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_9), .A2(n_91), .B1(n_636), .B2(n_637), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g940 ( .A1(n_10), .A2(n_59), .B1(n_941), .B2(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g942 ( .A(n_10), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_11), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_12), .A2(n_71), .B1(n_143), .B2(n_158), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_13), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_14), .A2(n_33), .B1(n_581), .B2(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g566 ( .A(n_15), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_16), .A2(n_64), .B1(n_137), .B2(n_177), .Y(n_239) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_17), .A2(n_70), .B(n_133), .Y(n_132) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_17), .A2(n_70), .B(n_133), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_18), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_19), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g564 ( .A(n_20), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_21), .B(n_180), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_22), .Y(n_269) );
BUFx3_ASAP7_75t_L g534 ( .A(n_23), .Y(n_534) );
BUFx8_ASAP7_75t_SL g956 ( .A(n_23), .Y(n_956) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_24), .A2(n_144), .B(n_209), .C(n_210), .Y(n_208) );
OAI22xp33_ASAP7_75t_SL g136 ( .A1(n_25), .A2(n_49), .B1(n_137), .B2(n_138), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_26), .A2(n_31), .B1(n_138), .B2(n_154), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_L g588 ( .A1(n_27), .A2(n_589), .B(n_592), .C(n_595), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_28), .B(n_576), .Y(n_575) );
O2A1O1Ixp5_ASAP7_75t_L g220 ( .A1(n_29), .A2(n_171), .B(n_221), .C(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g116 ( .A(n_30), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_30), .B(n_82), .Y(n_960) );
AND2x2_ASAP7_75t_L g963 ( .A(n_34), .B(n_964), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_35), .B(n_165), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_36), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_37), .A2(n_41), .B1(n_639), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_38), .A2(n_69), .B1(n_601), .B2(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_39), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g672 ( .A(n_40), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_42), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_43), .B(n_162), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_44), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_45), .A2(n_144), .B(n_562), .C(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g709 ( .A(n_46), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_47), .A2(n_939), .B1(n_940), .B2(n_943), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_47), .Y(n_943) );
INVx2_ASAP7_75t_L g603 ( .A(n_48), .Y(n_603) );
INVx1_ASAP7_75t_L g133 ( .A(n_50), .Y(n_133) );
AND2x4_ASAP7_75t_L g146 ( .A(n_51), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g214 ( .A(n_51), .B(n_147), .Y(n_214) );
INVx2_ASAP7_75t_L g665 ( .A(n_52), .Y(n_665) );
INVxp67_ASAP7_75t_SL g199 ( .A(n_53), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_53), .B(n_165), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_53), .A2(n_68), .B1(n_165), .B2(n_300), .Y(n_299) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_54), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_55), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_56), .Y(n_230) );
INVx2_ASAP7_75t_L g197 ( .A(n_57), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_58), .A2(n_171), .B(n_271), .C(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g941 ( .A(n_59), .Y(n_941) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_60), .Y(n_173) );
INVx1_ASAP7_75t_SL g593 ( .A(n_61), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_62), .B(n_180), .Y(n_179) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_63), .A2(n_79), .B1(n_157), .B2(n_159), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_65), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_66), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_67), .A2(n_104), .B1(n_957), .B2(n_965), .Y(n_103) );
NAND2xp33_ASAP7_75t_R g243 ( .A(n_68), .B(n_189), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_72), .A2(n_144), .B(n_594), .C(n_668), .Y(n_667) );
OR2x6_ASAP7_75t_L g113 ( .A(n_73), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g962 ( .A(n_73), .Y(n_962) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_74), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g695 ( .A(n_75), .Y(n_695) );
INVx1_ASAP7_75t_L g705 ( .A(n_76), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_77), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_78), .B(n_581), .Y(n_580) );
NOR2xp67_ASAP7_75t_L g558 ( .A(n_80), .B(n_221), .Y(n_558) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_81), .A2(n_171), .B(n_662), .C(n_664), .Y(n_661) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_81), .A2(n_171), .B(n_662), .C(n_664), .Y(n_688) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
INVx1_ASAP7_75t_L g525 ( .A(n_83), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_85), .A2(n_95), .B1(n_625), .B2(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g964 ( .A(n_86), .Y(n_964) );
BUFx5_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
INVx1_ASAP7_75t_L g155 ( .A(n_87), .Y(n_155) );
INVx2_ASAP7_75t_L g216 ( .A(n_88), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_89), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g275 ( .A(n_90), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_92), .Y(n_211) );
INVx2_ASAP7_75t_SL g147 ( .A(n_93), .Y(n_147) );
INVx1_ASAP7_75t_L g228 ( .A(n_94), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_96), .B(n_189), .Y(n_706) );
INVx1_ASAP7_75t_SL g656 ( .A(n_97), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_98), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g233 ( .A(n_99), .Y(n_233) );
AND2x2_ASAP7_75t_L g629 ( .A(n_100), .B(n_188), .Y(n_629) );
OAI21xp33_ASAP7_75t_SL g267 ( .A1(n_101), .A2(n_137), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_SL g602 ( .A(n_102), .Y(n_602) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_531), .B(n_535), .Y(n_104) );
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_117), .B(n_528), .Y(n_105) );
INVx3_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
BUFx8_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx10_ASAP7_75t_L g530 ( .A(n_109), .Y(n_530) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OR2x6_ASAP7_75t_L g935 ( .A(n_112), .B(n_936), .Y(n_935) );
INVx8_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g542 ( .A(n_113), .B(n_543), .Y(n_542) );
OR2x6_ASAP7_75t_L g954 ( .A(n_113), .B(n_543), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI22x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_524), .B2(n_527), .Y(n_120) );
INVx1_ASAP7_75t_L g538 ( .A(n_121), .Y(n_538) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g946 ( .A(n_122), .Y(n_946) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_415), .Y(n_122) );
NAND4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_312), .C(n_352), .D(n_386), .Y(n_123) );
AOI211xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_182), .B(n_244), .C(n_303), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_148), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_126), .A2(n_289), .B1(n_399), .B2(n_401), .Y(n_398) );
BUFx3_ASAP7_75t_L g412 ( .A(n_126), .Y(n_412) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g261 ( .A(n_127), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_127), .B(n_316), .Y(n_342) );
AND2x4_ASAP7_75t_L g384 ( .A(n_127), .B(n_306), .Y(n_384) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g289 ( .A(n_128), .Y(n_289) );
AND2x2_ASAP7_75t_L g309 ( .A(n_128), .B(n_306), .Y(n_309) );
INVx2_ASAP7_75t_L g327 ( .A(n_128), .Y(n_327) );
AND2x2_ASAP7_75t_L g337 ( .A(n_128), .B(n_262), .Y(n_337) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_128), .Y(n_369) );
NAND2xp33_ASAP7_75t_R g465 ( .A(n_128), .B(n_262), .Y(n_465) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_134), .Y(n_128) );
INVx2_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_130), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_131), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_131), .B(n_216), .Y(n_215) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx3_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
INVx2_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_141), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AOI22xp33_ASAP7_75t_SL g172 ( .A1(n_137), .A2(n_138), .B1(n_173), .B2(n_174), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_137), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_137), .A2(n_138), .B1(n_192), .B2(n_193), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_137), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_137), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_137), .B(n_269), .Y(n_268) );
NAND2xp33_ASAP7_75t_L g556 ( .A(n_137), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g576 ( .A(n_137), .Y(n_576) );
INVx2_ASAP7_75t_L g581 ( .A(n_137), .Y(n_581) );
INVx2_ASAP7_75t_L g627 ( .A(n_137), .Y(n_627) );
INVx2_ASAP7_75t_L g636 ( .A(n_137), .Y(n_636) );
INVx1_ASAP7_75t_L g663 ( .A(n_137), .Y(n_663) );
INVx2_ASAP7_75t_SL g159 ( .A(n_138), .Y(n_159) );
INVx2_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
INVx1_ASAP7_75t_L g579 ( .A(n_138), .Y(n_579) );
INVx2_ASAP7_75t_L g591 ( .A(n_138), .Y(n_591) );
INVx1_ASAP7_75t_L g698 ( .A(n_138), .Y(n_698) );
INVx6_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g143 ( .A(n_139), .Y(n_143) );
INVx2_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx3_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
INVx3_ASAP7_75t_L g144 ( .A(n_140), .Y(n_144) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
INVx4_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_140), .B(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g598 ( .A(n_140), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B(n_145), .Y(n_141) );
INVx2_ASAP7_75t_L g601 ( .A(n_143), .Y(n_601) );
INVx1_ASAP7_75t_L g700 ( .A(n_143), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g170 ( .A1(n_144), .A2(n_146), .B1(n_171), .B2(n_172), .C(n_175), .Y(n_170) );
INVx3_ASAP7_75t_L g622 ( .A(n_144), .Y(n_622) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
INVx1_ASAP7_75t_L g242 ( .A(n_146), .Y(n_242) );
INVx3_ASAP7_75t_L g583 ( .A(n_146), .Y(n_583) );
AND2x2_ASAP7_75t_L g628 ( .A(n_146), .B(n_161), .Y(n_628) );
INVx2_ASAP7_75t_L g366 ( .A(n_148), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_148), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
AND2x2_ASAP7_75t_L g520 ( .A(n_148), .B(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_166), .Y(n_148) );
OR2x2_ASAP7_75t_L g336 ( .A(n_149), .B(n_306), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_161), .B(n_163), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_151), .A2(n_164), .B(n_279), .Y(n_278) );
OA22x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B1(n_156), .B2(n_160), .Y(n_151) );
INVx4_ASAP7_75t_L g595 ( .A(n_152), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_154), .A2(n_177), .B1(n_196), .B2(n_197), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_154), .B(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_154), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g626 ( .A(n_154), .Y(n_626) );
INVx2_ASAP7_75t_L g639 ( .A(n_154), .Y(n_639) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g158 ( .A(n_155), .Y(n_158) );
INVx1_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
INVx3_ASAP7_75t_L g594 ( .A(n_157), .Y(n_594) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_161), .B(n_186), .Y(n_658) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_162), .B(n_242), .Y(n_604) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g632 ( .A(n_165), .Y(n_632) );
AND2x4_ASAP7_75t_L g326 ( .A(n_166), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_167), .B(n_262), .Y(n_290) );
INVx2_ASAP7_75t_L g371 ( .A(n_167), .Y(n_371) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B(n_179), .Y(n_167) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_168), .A2(n_170), .B(n_179), .Y(n_306) );
NOR2x1_ASAP7_75t_SL g553 ( .A(n_168), .B(n_213), .Y(n_553) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OR2x2_ASAP7_75t_L g198 ( .A(n_169), .B(n_199), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_171), .A2(n_191), .B1(n_194), .B2(n_195), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_171), .A2(n_194), .B1(n_239), .B2(n_240), .Y(n_238) );
INVx1_ASAP7_75t_L g255 ( .A(n_171), .Y(n_255) );
INVx1_ASAP7_75t_L g559 ( .A(n_171), .Y(n_559) );
INVx2_ASAP7_75t_SL g640 ( .A(n_171), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_171), .B(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_171), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g209 ( .A(n_177), .Y(n_209) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_177), .Y(n_562) );
INVx2_ASAP7_75t_L g621 ( .A(n_177), .Y(n_621) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_180), .B(n_242), .Y(n_241) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx3_ASAP7_75t_L g231 ( .A(n_181), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_181), .B(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_181), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_217), .Y(n_182) );
AND2x2_ASAP7_75t_L g311 ( .A(n_183), .B(n_256), .Y(n_311) );
INVx2_ASAP7_75t_SL g319 ( .A(n_183), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_183), .A2(n_321), .B1(n_328), .B2(n_333), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_183), .B(n_217), .Y(n_339) );
AND2x2_ASAP7_75t_L g395 ( .A(n_183), .B(n_390), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_183), .B(n_282), .Y(n_515) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_200), .Y(n_183) );
INVx1_ASAP7_75t_L g403 ( .A(n_184), .Y(n_403) );
AND2x2_ASAP7_75t_L g480 ( .A(n_184), .B(n_236), .Y(n_480) );
OAI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_190), .B(n_198), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_186), .B(n_634), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_187), .B(n_214), .Y(n_279) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
INVx1_ASAP7_75t_L g265 ( .A(n_189), .Y(n_265) );
INVx2_ASAP7_75t_L g301 ( .A(n_189), .Y(n_301) );
INVx1_ASAP7_75t_L g612 ( .A(n_189), .Y(n_612) );
INVx1_ASAP7_75t_L g253 ( .A(n_191), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_194), .A2(n_226), .B1(n_227), .B2(n_229), .Y(n_225) );
INVx2_ASAP7_75t_L g252 ( .A(n_194), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_SL g694 ( .A1(n_194), .A2(n_695), .B(n_696), .C(n_699), .Y(n_694) );
INVx1_ASAP7_75t_L g254 ( .A(n_195), .Y(n_254) );
AND2x2_ASAP7_75t_L g247 ( .A(n_200), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g285 ( .A(n_200), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_200), .B(n_218), .Y(n_302) );
INVx2_ASAP7_75t_L g332 ( .A(n_200), .Y(n_332) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_200), .Y(n_351) );
INVx1_ASAP7_75t_L g385 ( .A(n_200), .Y(n_385) );
OR2x2_ASAP7_75t_L g431 ( .A(n_200), .B(n_248), .Y(n_431) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_200), .Y(n_448) );
AO31x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_207), .A3(n_212), .B(n_215), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_205), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_209), .A2(n_600), .B1(n_602), .B2(n_603), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g219 ( .A(n_213), .B(n_220), .C(n_225), .Y(n_219) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_213), .A2(n_252), .B1(n_253), .B2(n_254), .C(n_255), .Y(n_251) );
NOR4xp25_ASAP7_75t_L g687 ( .A(n_213), .B(n_606), .C(n_667), .D(n_688), .Y(n_687) );
INVx4_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g264 ( .A(n_214), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g361 ( .A(n_217), .B(n_247), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_217), .B(n_284), .Y(n_372) );
AND2x4_ASAP7_75t_L g429 ( .A(n_217), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_235), .Y(n_217) );
INVx2_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
AND2x2_ASAP7_75t_L g331 ( .A(n_218), .B(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_R g349 ( .A(n_218), .Y(n_349) );
INVx2_ASAP7_75t_L g391 ( .A(n_218), .Y(n_391) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_218), .Y(n_408) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_231), .B(n_232), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g226 ( .A(n_222), .Y(n_226) );
INVx1_ASAP7_75t_L g271 ( .A(n_222), .Y(n_271) );
INVx2_ASAP7_75t_L g574 ( .A(n_222), .Y(n_574) );
INVx2_ASAP7_75t_L g637 ( .A(n_222), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_231), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g570 ( .A(n_231), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
AND2x2_ASAP7_75t_L g390 ( .A(n_236), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
AND2x2_ASAP7_75t_L g298 ( .A(n_237), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_241), .Y(n_237) );
OAI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_259), .B1(n_280), .B2(n_286), .C(n_291), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_256), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_247), .B(n_349), .Y(n_427) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_247), .Y(n_490) );
AND2x2_ASAP7_75t_L g284 ( .A(n_248), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_248), .B(n_257), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_248), .B(n_438), .Y(n_503) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
AND2x2_ASAP7_75t_L g297 ( .A(n_250), .B(n_298), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_252), .A2(n_267), .B(n_270), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_252), .A2(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g433 ( .A(n_256), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g493 ( .A(n_256), .B(n_364), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_256), .B(n_350), .Y(n_523) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OR2x2_ASAP7_75t_L g457 ( .A(n_257), .B(n_316), .Y(n_457) );
AND2x2_ASAP7_75t_L g378 ( .A(n_258), .B(n_332), .Y(n_378) );
INVx1_ASAP7_75t_SL g400 ( .A(n_258), .Y(n_400) );
INVx1_ASAP7_75t_L g439 ( .A(n_258), .Y(n_439) );
BUFx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_260), .B(n_382), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_276), .Y(n_260) );
INVx2_ASAP7_75t_L g293 ( .A(n_261), .Y(n_293) );
INVx2_ASAP7_75t_L g316 ( .A(n_262), .Y(n_316) );
INVx2_ASAP7_75t_L g325 ( .A(n_262), .Y(n_325) );
INVx1_ASAP7_75t_L g365 ( .A(n_262), .Y(n_365) );
AND2x2_ASAP7_75t_L g405 ( .A(n_262), .B(n_371), .Y(n_405) );
OR2x2_ASAP7_75t_L g476 ( .A(n_262), .B(n_327), .Y(n_476) );
BUFx2_ASAP7_75t_L g483 ( .A(n_262), .Y(n_483) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AOI21x1_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .B(n_274), .Y(n_263) );
AND2x4_ASAP7_75t_L g383 ( .A(n_276), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_276), .B(n_340), .Y(n_396) );
INVx3_ASAP7_75t_L g406 ( .A(n_276), .Y(n_406) );
AND2x2_ASAP7_75t_L g440 ( .A(n_276), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g517 ( .A(n_276), .B(n_337), .Y(n_517) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g307 ( .A(n_277), .Y(n_307) );
AND2x2_ASAP7_75t_L g317 ( .A(n_277), .B(n_306), .Y(n_317) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g345 ( .A(n_278), .Y(n_345) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_281), .B(n_383), .Y(n_443) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
OR2x2_ASAP7_75t_L g318 ( .A(n_282), .B(n_319), .Y(n_318) );
NOR4xp25_ASAP7_75t_L g381 ( .A(n_282), .B(n_358), .C(n_382), .D(n_385), .Y(n_381) );
OR2x2_ASAP7_75t_L g468 ( .A(n_282), .B(n_469), .Y(n_468) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g508 ( .A(n_285), .B(n_447), .Y(n_508) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_288), .B(n_344), .Y(n_343) );
NOR2xp67_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g450 ( .A(n_289), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
O2A1O1Ixp33_ASAP7_75t_SL g353 ( .A1(n_292), .A2(n_354), .B(n_356), .C(n_360), .Y(n_353) );
INVx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g461 ( .A(n_293), .B(n_335), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g471 ( .A1(n_294), .A2(n_472), .B(n_474), .Y(n_471) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_302), .Y(n_295) );
OR2x2_ASAP7_75t_L g329 ( .A(n_296), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g458 ( .A(n_296), .Y(n_458) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g414 ( .A(n_297), .B(n_391), .Y(n_414) );
INVx1_ASAP7_75t_L g447 ( .A(n_297), .Y(n_447) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g606 ( .A(n_301), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_301), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g499 ( .A(n_302), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_308), .B(n_310), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI32xp33_ASAP7_75t_L g338 ( .A1(n_305), .A2(n_339), .A3(n_340), .B1(n_343), .B2(n_346), .Y(n_338) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g478 ( .A(n_308), .Y(n_478) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g441 ( .A(n_309), .B(n_325), .Y(n_441) );
OAI322xp33_ASAP7_75t_L g518 ( .A1(n_310), .A2(n_371), .A3(n_376), .B1(n_473), .B2(n_483), .C1(n_519), .C2(n_522), .Y(n_518) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_338), .Y(n_312) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B(n_320), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx2_ASAP7_75t_L g496 ( .A(n_323), .Y(n_496) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g359 ( .A(n_325), .Y(n_359) );
AND2x2_ASAP7_75t_L g464 ( .A(n_325), .B(n_345), .Y(n_464) );
AND2x2_ASAP7_75t_L g504 ( .A(n_326), .B(n_406), .Y(n_504) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g479 ( .A(n_331), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g389 ( .A(n_332), .Y(n_389) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g355 ( .A(n_336), .Y(n_355) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g376 ( .A(n_342), .B(n_345), .Y(n_376) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_345), .B(n_369), .Y(n_495) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g436 ( .A(n_351), .B(n_437), .Y(n_436) );
NOR4xp25_ASAP7_75t_L g352 ( .A(n_353), .B(n_362), .C(n_373), .D(n_381), .Y(n_352) );
INVx2_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_357), .A2(n_424), .B1(n_425), .B2(n_428), .C(n_432), .Y(n_423) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_359), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B(n_372), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_365), .B(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_378), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g502 ( .A(n_378), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g469 ( .A(n_380), .B(n_389), .Y(n_469) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g419 ( .A(n_384), .B(n_406), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_384), .B(n_406), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_384), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_384), .B(n_483), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g501 ( .A(n_384), .B(n_463), .Y(n_501) );
INVx1_ASAP7_75t_SL g509 ( .A(n_384), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_385), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g434 ( .A(n_385), .Y(n_434) );
INVx1_ASAP7_75t_L g491 ( .A(n_385), .Y(n_491) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_392), .B(n_393), .C(n_409), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g486 ( .A(n_390), .Y(n_486) );
INVx1_ASAP7_75t_L g438 ( .A(n_391), .Y(n_438) );
OAI21xp33_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_396), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_398), .B(n_404), .C(n_406), .D(n_407), .Y(n_397) );
OR2x2_ASAP7_75t_L g401 ( .A(n_400), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g449 ( .A(n_405), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g475 ( .A(n_406), .B(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g473 ( .A(n_407), .B(n_431), .Y(n_473) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .C(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g489 ( .A(n_410), .Y(n_489) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_412), .B(n_467), .Y(n_466) );
AOI21xp33_ASAP7_75t_SL g462 ( .A1(n_413), .A2(n_463), .B(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_451), .C(n_505), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B(n_423), .C(n_442), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g459 ( .A(n_427), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_428), .A2(n_507), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g485 ( .A(n_431), .B(n_486), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B(n_440), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_435), .A2(n_501), .B1(n_502), .B2(n_504), .Y(n_500) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_449), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_470), .C(n_487), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_466), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_458), .B1(n_459), .B2(n_460), .C(n_462), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g512 ( .A(n_469), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_477), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g521 ( .A(n_476), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_481), .B2(n_484), .Y(n_477) );
AND2x4_ASAP7_75t_L g498 ( .A(n_480), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_492), .B1(n_494), .B2(n_497), .C(n_500), .Y(n_487) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .C(n_518), .Y(n_505) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_513), .B(n_516), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVxp67_ASAP7_75t_SL g527 ( .A(n_524), .Y(n_527) );
NAND2xp33_ASAP7_75t_SL g948 ( .A(n_528), .B(n_949), .Y(n_948) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_944), .B(n_955), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_937), .Y(n_536) );
OAI22x1_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_544), .B2(n_932), .Y(n_537) );
INVx4_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx8_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g947 ( .A(n_542), .Y(n_947) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_545), .A2(n_935), .B1(n_946), .B2(n_947), .Y(n_945) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_822), .Y(n_545) );
NOR4xp75_ASAP7_75t_SL g546 ( .A(n_547), .B(n_740), .C(n_786), .D(n_806), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_711), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_607), .B(n_613), .C(n_673), .Y(n_548) );
AOI222xp33_ASAP7_75t_L g887 ( .A1(n_549), .A2(n_854), .B1(n_888), .B2(n_891), .C1(n_895), .C2(n_901), .Y(n_887) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_567), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g675 ( .A(n_551), .B(n_585), .Y(n_675) );
INVx1_ASAP7_75t_L g723 ( .A(n_551), .Y(n_723) );
INVx1_ASAP7_75t_L g852 ( .A(n_551), .Y(n_852) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g691 ( .A(n_552), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g714 ( .A(n_552), .Y(n_714) );
OR2x2_ASAP7_75t_L g746 ( .A(n_552), .B(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g789 ( .A(n_552), .B(n_692), .Y(n_789) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_552), .Y(n_796) );
AND2x2_ASAP7_75t_L g856 ( .A(n_552), .B(n_747), .Y(n_856) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .A3(n_560), .B(n_565), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B(n_559), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_559), .A2(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVxp67_ASAP7_75t_L g751 ( .A(n_567), .Y(n_751) );
INVx1_ASAP7_75t_L g931 ( .A(n_567), .Y(n_931) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_585), .Y(n_567) );
AND2x2_ASAP7_75t_L g676 ( .A(n_568), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g798 ( .A(n_568), .B(n_693), .Y(n_798) );
INVx2_ASAP7_75t_L g803 ( .A(n_568), .Y(n_803) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI21x1_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B(n_584), .Y(n_569) );
OAI21x1_ASAP7_75t_L g710 ( .A1(n_570), .A2(n_583), .B(n_706), .Y(n_710) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_571), .A2(n_584), .B(n_611), .Y(n_610) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_577), .B(n_582), .Y(n_571) );
INVx1_ASAP7_75t_L g650 ( .A(n_574), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_576), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_582), .B(n_632), .Y(n_654) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g769 ( .A(n_585), .B(n_610), .Y(n_769) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g609 ( .A(n_586), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_586), .B(n_852), .Y(n_851) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g677 ( .A(n_587), .Y(n_677) );
INVx1_ASAP7_75t_L g736 ( .A(n_587), .Y(n_736) );
OA21x2_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_596), .B(n_605), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_595), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_595), .B(n_649), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B(n_604), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_597), .A2(n_635), .B1(n_638), .B2(n_640), .Y(n_634) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_601), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_601), .B(n_669), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g843 ( .A1(n_607), .A2(n_844), .B(n_845), .Y(n_843) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g774 ( .A(n_608), .B(n_691), .Y(n_774) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g715 ( .A(n_609), .Y(n_715) );
AND2x2_ASAP7_75t_L g724 ( .A(n_610), .B(n_693), .Y(n_724) );
BUFx2_ASAP7_75t_L g821 ( .A(n_610), .Y(n_821) );
OR2x2_ASAP7_75t_L g866 ( .A(n_610), .B(n_746), .Y(n_866) );
OA21x2_ASAP7_75t_L g682 ( .A1(n_611), .A2(n_642), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_612), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_643), .Y(n_614) );
INVx1_ASAP7_75t_L g863 ( .A(n_615), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_630), .Y(n_615) );
AND2x4_ASAP7_75t_L g685 ( .A(n_616), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g719 ( .A(n_616), .B(n_657), .Y(n_719) );
BUFx2_ASAP7_75t_SL g727 ( .A(n_616), .Y(n_727) );
INVx1_ASAP7_75t_L g739 ( .A(n_616), .Y(n_739) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2x1_ASAP7_75t_L g758 ( .A(n_617), .B(n_718), .Y(n_758) );
INVx2_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g777 ( .A(n_618), .Y(n_777) );
AO31x2_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_623), .A3(n_628), .B(n_629), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_622), .A2(n_652), .B(n_654), .Y(n_651) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g703 ( .A(n_627), .Y(n_703) );
AND2x2_ASAP7_75t_L g805 ( .A(n_630), .B(n_734), .Y(n_805) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g717 ( .A(n_631), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g842 ( .A(n_631), .B(n_645), .Y(n_842) );
AOI21x1_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_641), .Y(n_631) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NOR2x1_ASAP7_75t_L g825 ( .A(n_643), .B(n_826), .Y(n_825) );
OR2x2_ASAP7_75t_L g880 ( .A(n_643), .B(n_727), .Y(n_880) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_644), .B(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_L g783 ( .A(n_644), .B(n_727), .Y(n_783) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_657), .Y(n_644) );
AND2x2_ASAP7_75t_L g729 ( .A(n_645), .B(n_682), .Y(n_729) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g734 ( .A(n_646), .Y(n_734) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g718 ( .A(n_647), .Y(n_718) );
AOI21x1_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_655), .Y(n_647) );
NOR2x1_ASAP7_75t_L g864 ( .A(n_657), .B(n_718), .Y(n_864) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B(n_670), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_666), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g686 ( .A(n_671), .B(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_678), .B1(n_684), .B2(n_689), .Y(n_673) );
NOR2xp33_ASAP7_75t_SL g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_675), .B(n_785), .Y(n_922) );
AND2x2_ASAP7_75t_L g690 ( .A(n_676), .B(n_691), .Y(n_690) );
NAND2x1_ASAP7_75t_SL g808 ( .A(n_676), .B(n_796), .Y(n_808) );
INVx2_ASAP7_75t_SL g745 ( .A(n_677), .Y(n_745) );
AND2x2_ASAP7_75t_L g878 ( .A(n_677), .B(n_692), .Y(n_878) );
BUFx2_ASAP7_75t_L g925 ( .A(n_677), .Y(n_925) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_679), .A2(n_817), .B(n_818), .C(n_820), .Y(n_816) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2x1p5_ASAP7_75t_L g757 ( .A(n_681), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g773 ( .A(n_681), .Y(n_773) );
INVx2_ASAP7_75t_L g898 ( .A(n_681), .Y(n_898) );
INVx1_ASAP7_75t_L g902 ( .A(n_681), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_681), .B(n_892), .Y(n_915) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g765 ( .A(n_682), .Y(n_765) );
INVx1_ASAP7_75t_L g827 ( .A(n_682), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_682), .B(n_777), .Y(n_847) );
OR2x2_ASAP7_75t_L g889 ( .A(n_684), .B(n_890), .Y(n_889) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AND2x4_ASAP7_75t_L g761 ( .A(n_685), .B(n_717), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_685), .B(n_812), .Y(n_811) );
AND2x4_ASAP7_75t_L g871 ( .A(n_685), .B(n_841), .Y(n_871) );
AND2x2_ASAP7_75t_L g906 ( .A(n_685), .B(n_733), .Y(n_906) );
INVx1_ASAP7_75t_L g755 ( .A(n_686), .Y(n_755) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_686), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g776 ( .A(n_686), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_686), .B(n_920), .Y(n_919) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g844 ( .A(n_691), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_692), .B(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_701), .B(n_710), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_694), .A2(n_701), .B(n_710), .Y(n_747) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_697), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND3x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .C(n_707), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_716), .B1(n_720), .B2(n_725), .C(n_730), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_713), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx2_ASAP7_75t_SL g768 ( .A(n_714), .Y(n_768) );
AND2x4_ASAP7_75t_L g833 ( .A(n_714), .B(n_724), .Y(n_833) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_714), .Y(n_892) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
AND2x2_ASAP7_75t_L g794 ( .A(n_717), .B(n_727), .Y(n_794) );
AND2x2_ASAP7_75t_L g924 ( .A(n_717), .B(n_925), .Y(n_924) );
AND2x6_ASAP7_75t_SL g928 ( .A(n_717), .B(n_815), .Y(n_928) );
INVx1_ASAP7_75t_L g819 ( .A(n_718), .Y(n_819) );
AND2x2_ASAP7_75t_L g772 ( .A(n_719), .B(n_773), .Y(n_772) );
AND2x4_ASAP7_75t_L g840 ( .A(n_719), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g927 ( .A(n_719), .Y(n_927) );
NOR4xp25_ASAP7_75t_L g730 ( .A(n_721), .B(n_731), .C(n_735), .D(n_737), .Y(n_730) );
INVx3_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g874 ( .A(n_722), .B(n_835), .Y(n_874) );
AND2x4_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_724), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g785 ( .A(n_724), .Y(n_785) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g775 ( .A(n_729), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g890 ( .A(n_729), .Y(n_890) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_732), .B(n_737), .Y(n_914) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g812 ( .A(n_734), .Y(n_812) );
INVx1_ASAP7_75t_L g920 ( .A(n_734), .Y(n_920) );
OR2x2_ASAP7_75t_L g845 ( .A(n_735), .B(n_789), .Y(n_845) );
AND2x2_ASAP7_75t_L g882 ( .A(n_735), .B(n_883), .Y(n_882) );
INVx2_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
BUFx2_ASAP7_75t_L g780 ( .A(n_736), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g926 ( .A1(n_737), .A2(n_746), .B1(n_750), .B2(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g804 ( .A(n_739), .B(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_741), .B(n_770), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_748), .B(n_752), .C(n_759), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
AND2x2_ASAP7_75t_L g839 ( .A(n_744), .B(n_798), .Y(n_839) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g797 ( .A(n_745), .B(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_745), .Y(n_830) );
INVx1_ASAP7_75t_L g858 ( .A(n_745), .Y(n_858) );
OR2x2_ASAP7_75t_L g930 ( .A(n_746), .B(n_931), .Y(n_930) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_747), .Y(n_750) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx2_ASAP7_75t_L g817 ( .A(n_750), .Y(n_817) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
AND2x2_ASAP7_75t_L g782 ( .A(n_754), .B(n_757), .Y(n_782) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_755), .B(n_815), .Y(n_838) );
AND2x2_ASAP7_75t_L g911 ( .A(n_755), .B(n_812), .Y(n_911) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g762 ( .A(n_758), .B(n_763), .Y(n_762) );
AOI21xp33_ASAP7_75t_SL g759 ( .A1(n_760), .A2(n_762), .B(n_766), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_760), .A2(n_847), .B1(n_848), .B2(n_853), .Y(n_846) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g855 ( .A1(n_761), .A2(n_856), .B1(n_857), .B2(n_861), .C(n_865), .Y(n_855) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g814 ( .A(n_764), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
OR2x2_ASAP7_75t_L g801 ( .A(n_768), .B(n_802), .Y(n_801) );
OR2x6_ASAP7_75t_L g859 ( .A(n_768), .B(n_860), .Y(n_859) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_769), .Y(n_869) );
INVx1_ASAP7_75t_L g894 ( .A(n_769), .Y(n_894) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_781), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B1(n_775), .B2(n_778), .Y(n_771) );
INVx1_ASAP7_75t_L g831 ( .A(n_772), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_776), .B(n_812), .Y(n_829) );
AND2x2_ASAP7_75t_L g901 ( .A(n_776), .B(n_902), .Y(n_901) );
BUFx3_ASAP7_75t_L g815 ( .A(n_777), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_778), .A2(n_825), .B(n_828), .Y(n_824) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B(n_784), .Y(n_781) );
INVx1_ASAP7_75t_L g791 ( .A(n_782), .Y(n_791) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_799), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .B1(n_792), .B2(n_795), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_788), .A2(n_901), .B1(n_906), .B2(n_907), .Y(n_905) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI21xp5_ASAP7_75t_SL g799 ( .A1(n_795), .A2(n_800), .B(n_804), .Y(n_799) );
AND2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx2_ASAP7_75t_L g850 ( .A(n_798), .Y(n_850) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g883 ( .A(n_802), .Y(n_883) );
BUFx2_ASAP7_75t_SL g860 ( .A(n_803), .Y(n_860) );
INVx1_ASAP7_75t_L g877 ( .A(n_803), .Y(n_877) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_809), .B(n_816), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g810 ( .A(n_811), .B(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g818 ( .A(n_814), .B(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_815), .B(n_864), .Y(n_900) );
INVx1_ASAP7_75t_L g907 ( .A(n_817), .Y(n_907) );
INVxp67_ASAP7_75t_L g836 ( .A(n_819), .Y(n_836) );
AOI21xp33_ASAP7_75t_L g913 ( .A1(n_820), .A2(n_914), .B(n_915), .Y(n_913) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_821), .A2(n_910), .B(n_912), .Y(n_909) );
NOR3xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_872), .C(n_903), .Y(n_822) );
NAND3xp33_ASAP7_75t_SL g823 ( .A(n_824), .B(n_834), .C(n_855), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2x1_ASAP7_75t_L g885 ( .A(n_827), .B(n_886), .Y(n_885) );
O2A1O1Ixp33_ASAP7_75t_SL g828 ( .A1(n_829), .A2(n_830), .B(n_831), .C(n_832), .Y(n_828) );
INVx1_ASAP7_75t_L g904 ( .A(n_830), .Y(n_904) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_839), .B1(n_840), .B2(n_843), .C(n_846), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g917 ( .A(n_847), .Y(n_917) );
INVx2_ASAP7_75t_SL g848 ( .A(n_849), .Y(n_848) );
NOR2x1_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
INVx1_ASAP7_75t_L g854 ( .A(n_850), .Y(n_854) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_L g868 ( .A(n_856), .Y(n_868) );
NOR2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_866), .A2(n_867), .B(n_870), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NAND3xp33_ASAP7_75t_L g872 ( .A(n_873), .B(n_881), .C(n_887), .Y(n_872) );
NOR2x1_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
NOR2x1_ASAP7_75t_L g875 ( .A(n_876), .B(n_879), .Y(n_875) );
NAND2x1p5_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g912 ( .A(n_878), .Y(n_912) );
BUFx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g886 ( .A(n_880), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_884), .Y(n_881) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
AND2x4_ASAP7_75t_L g895 ( .A(n_896), .B(n_899), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
OAI211xp5_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_905), .B(n_908), .C(n_923), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_913), .B1(n_916), .B2(n_921), .Y(n_908) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
AND2x2_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVxp33_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g923 ( .A1(n_924), .A2(n_926), .B1(n_928), .B2(n_929), .Y(n_923) );
INVxp67_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
BUFx12f_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
CKINVDCx11_ASAP7_75t_R g933 ( .A(n_934), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
AOI21xp33_ASAP7_75t_L g944 ( .A1(n_938), .A2(n_945), .B(n_948), .Y(n_944) );
INVxp67_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
BUFx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
BUFx3_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g955 ( .A(n_956), .Y(n_955) );
BUFx4_ASAP7_75t_SL g957 ( .A(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
BUFx2_ASAP7_75t_L g967 ( .A(n_959), .Y(n_967) );
OR2x2_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .Y(n_959) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_SL g966 ( .A(n_967), .Y(n_966) );
endmodule