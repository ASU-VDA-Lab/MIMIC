module fake_jpeg_11543_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_29),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_71),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_35),
.B1(n_20),
.B2(n_37),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_97),
.B(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_85),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_16),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_86),
.B(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_16),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_90),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_43),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_101),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_35),
.B1(n_27),
.B2(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_38),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_107),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_27),
.B1(n_37),
.B2(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_30),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_39),
.B1(n_36),
.B2(n_27),
.Y(n_111)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_104),
.B1(n_99),
.B2(n_66),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_137),
.B1(n_101),
.B2(n_68),
.Y(n_149)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_18),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_122),
.B(n_127),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_39),
.B1(n_36),
.B2(n_18),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_96),
.B1(n_87),
.B2(n_63),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_65),
.A2(n_24),
.B(n_21),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_122),
.C(n_115),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_0),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_69),
.A2(n_39),
.B1(n_17),
.B2(n_9),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_144),
.Y(n_178)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_142),
.Y(n_170)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_161),
.B1(n_173),
.B2(n_135),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_72),
.B(n_68),
.C(n_94),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_165),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_133),
.A2(n_68),
.B1(n_100),
.B2(n_66),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_141),
.C(n_120),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_124),
.C(n_129),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

BUFx12_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_113),
.B(n_103),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_177),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_128),
.A2(n_87),
.B1(n_103),
.B2(n_93),
.Y(n_173)
);

AO21x2_ASAP7_75t_L g174 ( 
.A1(n_111),
.A2(n_63),
.B(n_106),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_174),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_214)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_118),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_127),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_110),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_174),
.B1(n_150),
.B2(n_152),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_188),
.B1(n_199),
.B2(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_190),
.B(n_205),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_198),
.Y(n_221)
);

AOI21x1_ASAP7_75t_SL g194 ( 
.A1(n_178),
.A2(n_135),
.B(n_121),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_201),
.B(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_121),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_174),
.A2(n_81),
.B1(n_82),
.B2(n_74),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_142),
.B(n_114),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_74),
.B1(n_82),
.B2(n_81),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_168),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_150),
.A2(n_135),
.B1(n_114),
.B2(n_140),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_168),
.C(n_176),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_136),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_126),
.C(n_12),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_166),
.C(n_4),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_160),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_148),
.B1(n_171),
.B2(n_166),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_1),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_216),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_2),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_3),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_217),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_149),
.B1(n_146),
.B2(n_151),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_223),
.A2(n_240),
.B1(n_244),
.B2(n_214),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_148),
.B1(n_171),
.B2(n_151),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_238),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_235),
.C(n_207),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_230),
.B(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_162),
.B1(n_4),
.B2(n_5),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_184),
.B(n_194),
.Y(n_255)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_191),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_190),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_237),
.B(n_203),
.Y(n_264)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_162),
.B(n_13),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_206),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_243),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_3),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_SL g244 ( 
.A1(n_201),
.A2(n_184),
.B(n_192),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_221),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_246),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_223),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_216),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_258),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_192),
.Y(n_261)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_217),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_215),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_235),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_278),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_273),
.C(n_257),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_227),
.C(n_192),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_222),
.B1(n_245),
.B2(n_236),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_276),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_245),
.B1(n_241),
.B2(n_233),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_280),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_243),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_231),
.B1(n_229),
.B2(n_220),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_232),
.B(n_197),
.Y(n_280)
);

OA22x2_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_238),
.B1(n_210),
.B2(n_200),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_283),
.A2(n_256),
.B1(n_267),
.B2(n_260),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_254),
.B1(n_263),
.B2(n_262),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_247),
.B1(n_263),
.B2(n_265),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_297),
.C(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_266),
.B1(n_256),
.B2(n_265),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_295),
.B1(n_300),
.B2(n_275),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_261),
.C(n_253),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_299),
.C(n_286),
.Y(n_301)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_280),
.B(n_261),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_255),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_301),
.B(n_312),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_255),
.C(n_268),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_303),
.B(n_228),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_307),
.C(n_289),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_270),
.Y(n_307)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_264),
.B1(n_259),
.B2(n_284),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_311),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_282),
.C(n_274),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_320),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_288),
.B1(n_287),
.B2(n_290),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_305),
.B1(n_302),
.B2(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_310),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_283),
.C(n_296),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_323),
.Y(n_331)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_267),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_304),
.C(n_283),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_317),
.B1(n_321),
.B2(n_316),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_329),
.B(n_326),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_324),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.C(n_330),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_332),
.B(n_331),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_320),
.B(n_313),
.C(n_260),
.Y(n_337)
);

OAI321xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_249),
.A3(n_248),
.B1(n_259),
.B2(n_202),
.C(n_218),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_248),
.B(n_249),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_196),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_202),
.Y(n_341)
);


endmodule