module fake_jpeg_12790_n_86 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_28),
.B2(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_28),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_5),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_31),
.B1(n_36),
.B2(n_33),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_5),
.B(n_6),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_4),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_15),
.B(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_14),
.C(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_6),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_7),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_8),
.B(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_59),
.B1(n_10),
.B2(n_19),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_59),
.B1(n_13),
.B2(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_78),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_69),
.B(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_76),
.B1(n_79),
.B2(n_66),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_74),
.Y(n_85)
);

AOI221xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.C(n_27),
.Y(n_86)
);


endmodule