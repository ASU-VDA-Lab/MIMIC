module real_jpeg_6129_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_0),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_0),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_0),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_0),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_0),
.B(n_160),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_0),
.B(n_342),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_0),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_0),
.B(n_438),
.Y(n_437)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_2),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_2),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_2),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_3),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_3),
.B(n_35),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_3),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_3),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_3),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_3),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_4),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_4),
.B(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_4),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_4),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_4),
.B(n_356),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_4),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_5),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_5),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_5),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_5),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_5),
.B(n_200),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_5),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_5),
.B(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_6),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_6),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_6),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_6),
.B(n_227),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_6),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_6),
.B(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_6),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_6),
.B(n_53),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_7),
.Y(n_489)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_8),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g300 ( 
.A(n_9),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_9),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_9),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_9),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_9),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_9),
.B(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_10),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_10),
.Y(n_448)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_12),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_12),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_12),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_13),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_13),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g366 ( 
.A(n_13),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_13),
.B(n_447),
.Y(n_446)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_15),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_15),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_15),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_15),
.B(n_227),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_15),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_15),
.B(n_397),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_15),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_15),
.B(n_488),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_16),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_16),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_16),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_16),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_16),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_16),
.B(n_150),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_16),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_16),
.B(n_414),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_17),
.Y(n_549)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_19),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_19),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_19),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_19),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_19),
.B(n_227),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_19),
.B(n_37),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_544),
.B(n_547),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_80),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_46),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_61),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_40),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_28),
.B(n_390),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_29),
.B(n_165),
.Y(n_451)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_30),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_50),
.C(n_57),
.Y(n_77)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_42),
.Y(n_480)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_42),
.Y(n_505)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_43),
.Y(n_152)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_43),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_45),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_76),
.C(n_78),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_47),
.B(n_534),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_62),
.C(n_66),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_48),
.A2(n_49),
.B1(n_530),
.B2(n_531),
.Y(n_529)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_54),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_67),
.C(n_71),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_56),
.A2(n_57),
.B1(n_71),
.B2(n_490),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_60),
.Y(n_162)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_60),
.Y(n_263)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_60),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_62),
.B(n_66),
.Y(n_531)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_67),
.A2(n_68),
.B1(n_492),
.B2(n_493),
.Y(n_491)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_71),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_71),
.A2(n_445),
.B1(n_446),
.B2(n_490),
.Y(n_509)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_73),
.Y(n_231)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_74),
.Y(n_260)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_74),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_74),
.Y(n_401)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_74),
.Y(n_459)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_535),
.Y(n_534)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_78),
.Y(n_535)
);

AO21x1_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_463),
.B(n_537),
.Y(n_81)
);

OAI21x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_424),
.B(n_462),
.Y(n_82)
);

AOI21x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_377),
.B(n_423),
.Y(n_83)
);

OAI21x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_328),
.B(n_376),
.Y(n_84)
);

AOI21x1_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_290),
.B(n_327),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_211),
.B(n_289),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_191),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_88),
.B(n_191),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_133),
.B2(n_190),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_89),
.B(n_134),
.C(n_173),
.Y(n_326)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_113),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_91),
.B(n_114),
.C(n_132),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_105),
.C(n_109),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_92),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_99),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_93),
.A2(n_94),
.B1(n_99),
.B2(n_100),
.Y(n_196)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_98),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_98),
.Y(n_392)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_104),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_105),
.B(n_109),
.Y(n_210)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_107),
.Y(n_443)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_112),
.Y(n_320)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_112),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_121),
.B1(n_131),
.B2(n_132),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B(n_120),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.Y(n_120)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_120),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_120),
.B(n_295),
.C(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_122),
.B(n_124),
.C(n_127),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_173),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_146),
.C(n_163),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_193),
.Y(n_192)
);

BUFx24_ASAP7_75t_SL g552 ( 
.A(n_135),
.Y(n_552)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_139),
.CI(n_143),
.CON(n_135),
.SN(n_135)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_139),
.C(n_143),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_142),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_145),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_147),
.B1(n_163),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.C(n_158),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_148),
.A2(n_149),
.B1(n_158),
.B2(n_159),
.Y(n_282)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_152),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_153),
.B(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g454 ( 
.A(n_161),
.Y(n_454)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_165),
.B(n_472),
.Y(n_471)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_168),
.Y(n_304)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_187),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_174),
.B(n_188),
.C(n_189),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_175),
.B(n_182),
.C(n_185),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_209),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_192),
.B(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_209),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.C(n_202),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_196),
.B(n_197),
.Y(n_275)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_202),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_284),
.B(n_288),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_269),
.B(n_283),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_251),
.B(n_268),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_240),
.B(n_250),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_223),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_223),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_219),
.Y(n_365)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_232),
.B2(n_233),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_228),
.C(n_232),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_238),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_245),
.B(n_249),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_244),
.Y(n_404)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_267),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_267),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_255),
.C(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_264),
.C(n_266),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx11_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_263),
.Y(n_398)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_272),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_279),
.C(n_280),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_326),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_291),
.B(n_326),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_308),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_294),
.C(n_308),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_305),
.B2(n_307),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_300),
.C(n_302),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_311),
.C(n_321),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_321),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_317),
.C(n_318),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_329),
.B(n_330),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_331),
.B(n_348),
.C(n_374),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_348),
.B1(n_374),
.B2(n_375),
.Y(n_332)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_336),
.B2(n_347),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_337),
.C(n_338),
.Y(n_379)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_336),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_346),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_340),
.B(n_341),
.C(n_346),
.Y(n_410)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_359),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_360),
.C(n_361),
.Y(n_408)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_349),
.Y(n_550)
);

FAx1_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_353),
.CI(n_355),
.CON(n_349),
.SN(n_349)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_350),
.B(n_353),
.C(n_355),
.Y(n_420)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_370),
.B2(n_371),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_366),
.B1(n_368),
.B2(n_369),
.Y(n_363)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_364),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_369),
.C(n_370),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_366),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_366),
.A2(n_369),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_369),
.B(n_384),
.C(n_389),
.Y(n_435)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_422),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_378),
.B(n_422),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_379),
.B(n_381),
.C(n_406),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_406),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_393),
.B2(n_405),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_382),
.B(n_394),
.C(n_395),
.Y(n_429)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_388),
.A2(n_389),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_388),
.B(n_442),
.C(n_445),
.Y(n_510)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_393),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_450),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_395),
.B(n_441),
.C(n_450),
.Y(n_469)
);

FAx1_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_399),
.CI(n_402),
.CON(n_395),
.SN(n_395)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_409),
.B2(n_421),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_410),
.C(n_411),
.Y(n_426)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_420),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_415),
.B1(n_418),
.B2(n_419),
.Y(n_412)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_413),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_415),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_418),
.C(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_415),
.A2(n_419),
.B1(n_437),
.B2(n_439),
.Y(n_436)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_435),
.C(n_439),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_420),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_461),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_461),
.Y(n_462)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_425),
.Y(n_553)
);

FAx1_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.CI(n_440),
.CON(n_425),
.SN(n_425)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_426),
.B(n_427),
.C(n_440),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_428),
.B(n_432),
.C(n_434),
.Y(n_518)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_449),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_487),
.C(n_490),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_451),
.B(n_455),
.C(n_460),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_455),
.B1(n_456),
.B2(n_460),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_453),
.Y(n_460)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_522),
.C(n_532),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_519),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_466),
.A2(n_541),
.B(n_542),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_512),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_467),
.B(n_512),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_483),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_468),
.B(n_484),
.C(n_507),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.C(n_481),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_469),
.B(n_514),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_481),
.B1(n_482),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_474),
.C(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_507),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_496),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_491),
.B1(n_494),
.B2(n_495),
.Y(n_485)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_486),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_486),
.B(n_495),
.C(n_496),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_491),
.Y(n_495)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_497),
.B(n_500),
.C(n_506),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_500),
.B1(n_501),
.B2(n_506),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_499),
.Y(n_506)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.C(n_511),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_508),
.B(n_517),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_511),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_516),
.C(n_518),
.Y(n_512)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_513),
.B(n_516),
.CI(n_518),
.CON(n_520),
.SN(n_520)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_521),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_521),
.Y(n_541)
);

BUFx24_ASAP7_75t_SL g551 ( 
.A(n_520),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_540),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_525),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_527),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_528),
.C(n_529),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

A2O1A1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_532),
.A2(n_538),
.B(n_539),
.C(n_543),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_536),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_536),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

BUFx12f_ASAP7_75t_L g548 ( 
.A(n_545),
.Y(n_548)
);

INVx13_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_549),
.Y(n_547)
);


endmodule