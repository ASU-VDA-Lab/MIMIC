module fake_jpeg_28564_n_363 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_363);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_363;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_50),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_36),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_52),
.Y(n_95)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_19),
.B(n_14),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_11),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_54),
.B(n_24),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_58),
.Y(n_106)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_0),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_38),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_70),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_28),
.B(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_1),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_80),
.Y(n_121)
);

CKINVDCx9p33_ASAP7_75t_R g81 ( 
.A(n_30),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_81),
.Y(n_120)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_84),
.B1(n_32),
.B2(n_26),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_46),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_83),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_86),
.A2(n_112),
.B1(n_123),
.B2(n_63),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_91),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_49),
.A2(n_18),
.B1(n_16),
.B2(n_25),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_110),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_41),
.C(n_18),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_93),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_45),
.B(n_16),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_102),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_18),
.B1(n_39),
.B2(n_33),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_60),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_137),
.B1(n_24),
.B2(n_65),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_59),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

INVx2_ASAP7_75t_R g122 ( 
.A(n_57),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_130),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_55),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_124),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_26),
.C(n_25),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_138),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_44),
.B(n_26),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_51),
.B(n_25),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_66),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_134),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_69),
.A2(n_43),
.B1(n_42),
.B2(n_27),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_136),
.B1(n_4),
.B2(n_5),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_43),
.B1(n_42),
.B2(n_27),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_61),
.A2(n_43),
.B1(n_42),
.B2(n_27),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_67),
.B(n_24),
.C(n_2),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_2),
.Y(n_156)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_143),
.A2(n_155),
.B1(n_172),
.B2(n_174),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_95),
.A2(n_73),
.B1(n_62),
.B2(n_76),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_160),
.B1(n_161),
.B2(n_166),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_95),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

AOI22x1_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_78),
.B1(n_77),
.B2(n_3),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_150),
.A2(n_167),
.B1(n_175),
.B2(n_145),
.Y(n_206)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_101),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_154),
.B(n_156),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_122),
.B1(n_87),
.B2(n_90),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_6),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_169),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_128),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_92),
.B1(n_139),
.B2(n_89),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_176),
.B1(n_183),
.B2(n_184),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_106),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_171),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_118),
.A2(n_103),
.B1(n_96),
.B2(n_139),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_118),
.A2(n_103),
.B1(n_96),
.B2(n_117),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_133),
.A2(n_121),
.B1(n_109),
.B2(n_104),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_135),
.A2(n_136),
.B1(n_131),
.B2(n_104),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_107),
.B(n_94),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_132),
.Y(n_202)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_114),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_181),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_114),
.A2(n_99),
.B1(n_108),
.B2(n_129),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_182),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_127),
.A2(n_131),
.B1(n_108),
.B2(n_129),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_127),
.A2(n_99),
.B1(n_94),
.B2(n_111),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_111),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_186),
.Y(n_190)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_113),
.B(n_132),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_197),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_113),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_199),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_159),
.B(n_113),
.Y(n_197)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_132),
.A3(n_164),
.B1(n_151),
.B2(n_142),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_218),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_151),
.A2(n_177),
.B(n_150),
.C(n_152),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_206),
.A2(n_210),
.B1(n_217),
.B2(n_191),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_157),
.B(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_213),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_143),
.A2(n_165),
.B1(n_151),
.B2(n_175),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_178),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_156),
.C(n_158),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_216),
.B(n_193),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_170),
.C(n_154),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_147),
.B1(n_150),
.B2(n_141),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_141),
.B(n_166),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_146),
.B(n_163),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_195),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_162),
.B(n_171),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_189),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_181),
.B(n_180),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_228),
.B(n_246),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_227),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_197),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_173),
.B(n_186),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_240),
.Y(n_272)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_183),
.B1(n_179),
.B2(n_153),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_237),
.Y(n_260)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx6_ASAP7_75t_SL g237 ( 
.A(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_241),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_185),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_243),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_149),
.B1(n_194),
.B2(n_189),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_254),
.B1(n_211),
.B2(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_248),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_204),
.B1(n_216),
.B2(n_214),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_213),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_249),
.B(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_194),
.B(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_252),
.B1(n_220),
.B2(n_215),
.Y(n_262)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_205),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_212),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_191),
.A2(n_206),
.B1(n_224),
.B2(n_196),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_275),
.B1(n_232),
.B2(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_238),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_215),
.B1(n_222),
.B2(n_220),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_261),
.A2(n_240),
.B1(n_252),
.B2(n_245),
.Y(n_299)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_221),
.C(n_211),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_266),
.C(n_271),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_267),
.B1(n_276),
.B2(n_231),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_249),
.C(n_248),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_254),
.A2(n_242),
.B1(n_250),
.B2(n_234),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_231),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_243),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_235),
.B(n_233),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_242),
.A2(n_231),
.B1(n_227),
.B2(n_233),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_242),
.A2(n_247),
.B1(n_235),
.B2(n_231),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_225),
.A2(n_228),
.B(n_247),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_260),
.B(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_288),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_226),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_295),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_281),
.A2(n_257),
.B(n_269),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_258),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_291),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_237),
.B1(n_245),
.B2(n_236),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_284),
.A2(n_236),
.B1(n_273),
.B2(n_255),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_251),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_287),
.A2(n_289),
.B1(n_296),
.B2(n_299),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_256),
.B1(n_278),
.B2(n_261),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_232),
.C(n_230),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_264),
.C(n_268),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_263),
.B(n_278),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_265),
.B1(n_274),
.B2(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_260),
.Y(n_308)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_266),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_307),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_312),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_288),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_282),
.B(n_257),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_262),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_269),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_313),
.A2(n_284),
.B1(n_299),
.B2(n_296),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_255),
.C(n_297),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_298),
.C(n_297),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_319),
.C(n_323),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_292),
.B1(n_283),
.B2(n_291),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_318),
.A2(n_305),
.B1(n_304),
.B2(n_283),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_279),
.C(n_281),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_314),
.B1(n_315),
.B2(n_308),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_306),
.B(n_280),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_321),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_289),
.C(n_287),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_300),
.Y(n_324)
);

AOI21xp33_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_329),
.B(n_330),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_327),
.A2(n_301),
.B(n_300),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_285),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_316),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_336),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_309),
.B(n_314),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_318),
.B(n_323),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_335),
.A2(n_338),
.B1(n_340),
.B2(n_333),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_307),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_303),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_337),
.B(n_322),
.Y(n_345)
);

A2O1A1O1Ixp25_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_327),
.B(n_330),
.C(n_319),
.D(n_325),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_304),
.B1(n_286),
.B2(n_290),
.Y(n_340)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_342),
.B(n_340),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_339),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_345),
.Y(n_350)
);

AOI21xp33_ASAP7_75t_L g347 ( 
.A1(n_341),
.A2(n_326),
.B(n_331),
.Y(n_347)
);

NOR2x1_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_332),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_338),
.B1(n_337),
.B2(n_335),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_353),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_351),
.B(n_334),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_354),
.A2(n_351),
.B(n_334),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_350),
.B(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_353),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_359),
.A2(n_358),
.B(n_356),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_360),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_352),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_362),
.B(n_336),
.Y(n_363)
);


endmodule