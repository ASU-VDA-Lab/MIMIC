module fake_jpeg_27784_n_30 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_3),
.B(n_2),
.Y(n_9)
);

BUFx24_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_7),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_6),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_11),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_16),
.B1(n_15),
.B2(n_8),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_21),
.C(n_22),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_11),
.A2(n_12),
.B(n_14),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_10),
.B(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_10),
.Y(n_23)
);

OAI221xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.C(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_26),
.C(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);


endmodule