module fake_jpeg_11324_n_464 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_464);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_464;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_14),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_59),
.Y(n_98)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_6),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_49),
.B(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_51),
.Y(n_141)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_6),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_7),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_54),
.B(n_35),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_61),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_7),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_73),
.Y(n_113)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx6f_ASAP7_75t_SL g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_78),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_26),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_89),
.Y(n_128)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_16),
.B(n_5),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_27),
.Y(n_144)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_100),
.B(n_88),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_51),
.A2(n_21),
.B1(n_55),
.B2(n_46),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_102),
.A2(n_114),
.B1(n_148),
.B2(n_17),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_44),
.B1(n_45),
.B2(n_22),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_105),
.A2(n_112),
.B1(n_15),
.B2(n_35),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_68),
.A2(n_45),
.B1(n_24),
.B2(n_44),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_21),
.B1(n_46),
.B2(n_43),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_27),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_119),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_42),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_78),
.B(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_146),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_37),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_32),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_62),
.A2(n_43),
.B1(n_44),
.B2(n_24),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_155),
.A2(n_143),
.B1(n_130),
.B2(n_136),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_67),
.B1(n_69),
.B2(n_92),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_96),
.B1(n_143),
.B2(n_130),
.Y(n_198)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_176),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_163),
.B(n_171),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_98),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_173),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_116),
.A2(n_70),
.B1(n_48),
.B2(n_17),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_179),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_37),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_108),
.B(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_178),
.Y(n_215)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_87),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_186),
.B1(n_190),
.B2(n_122),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_29),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_57),
.B1(n_64),
.B2(n_71),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_193),
.B1(n_141),
.B2(n_117),
.Y(n_219)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

BUFx24_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_139),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_187),
.Y(n_206)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_102),
.A2(n_66),
.B1(n_52),
.B2(n_63),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_122),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_124),
.B(n_86),
.C(n_72),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_192),
.C(n_117),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_139),
.B(n_88),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_79),
.C(n_76),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_114),
.A2(n_24),
.B1(n_15),
.B2(n_43),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_123),
.B(n_32),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_17),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_198),
.A2(n_207),
.B1(n_213),
.B2(n_153),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_97),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_209),
.B(n_229),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_155),
.A2(n_115),
.B1(n_135),
.B2(n_149),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_131),
.B1(n_136),
.B2(n_135),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_214),
.A2(n_219),
.B1(n_159),
.B2(n_186),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_220),
.B(n_129),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_177),
.A2(n_140),
.B1(n_131),
.B2(n_147),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_161),
.B1(n_183),
.B2(n_185),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_157),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_230),
.A2(n_238),
.B1(n_241),
.B2(n_250),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_168),
.B1(n_192),
.B2(n_166),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_162),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_239),
.B(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_176),
.C(n_151),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_240),
.B(n_251),
.C(n_228),
.Y(n_279)
);

OAI22x1_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_170),
.B1(n_140),
.B2(n_134),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_170),
.B(n_97),
.C(n_134),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_198),
.A2(n_175),
.B1(n_115),
.B2(n_158),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_246),
.B1(n_257),
.B2(n_182),
.Y(n_261)
);

AND2x6_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_134),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_254),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_199),
.A2(n_167),
.B1(n_150),
.B2(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_180),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_253),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_201),
.A2(n_164),
.B1(n_156),
.B2(n_149),
.Y(n_250)
);

INVx11_ASAP7_75t_L g252 ( 
.A(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_252),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_152),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_206),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_211),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_200),
.B(n_84),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_147),
.B1(n_58),
.B2(n_74),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_206),
.B(n_223),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_206),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_279),
.C(n_283),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_212),
.B1(n_226),
.B2(n_205),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_267),
.A2(n_270),
.B1(n_284),
.B2(n_188),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_221),
.B(n_211),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_280),
.B(n_165),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_260),
.A2(n_205),
.B1(n_227),
.B2(n_202),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_230),
.A2(n_227),
.B1(n_202),
.B2(n_228),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_274),
.A2(n_290),
.B1(n_248),
.B2(n_234),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_231),
.A2(n_211),
.B(n_223),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_225),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_246),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_225),
.Y(n_283)
);

OAI22x1_ASAP7_75t_SL g284 ( 
.A1(n_237),
.A2(n_241),
.B1(n_242),
.B2(n_245),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_251),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_253),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_289),
.B(n_33),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_250),
.A2(n_203),
.B1(n_216),
.B2(n_196),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_263),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_295),
.Y(n_322)
);

AO22x1_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_243),
.B1(n_247),
.B2(n_244),
.Y(n_294)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_296),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_272),
.A2(n_257),
.B(n_233),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_297),
.B(n_305),
.Y(n_349)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_300),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_256),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_301),
.B(n_303),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_240),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_309),
.C(n_80),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_239),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_273),
.A2(n_265),
.B1(n_278),
.B2(n_272),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_304),
.A2(n_311),
.B1(n_315),
.B2(n_270),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_278),
.B(n_254),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_236),
.Y(n_306)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_267),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_307),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_255),
.C(n_252),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_310),
.A2(n_276),
.B(n_288),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_273),
.A2(n_203),
.B1(n_217),
.B2(n_216),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_217),
.Y(n_312)
);

OAI21xp33_ASAP7_75t_R g330 ( 
.A1(n_312),
.A2(n_282),
.B(n_276),
.Y(n_330)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_313),
.A2(n_274),
.B(n_268),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_265),
.A2(n_29),
.B1(n_204),
.B2(n_197),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_287),
.B(n_197),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_316),
.B(n_27),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_287),
.A2(n_204),
.B(n_154),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_320),
.B(n_280),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_261),
.A2(n_184),
.B1(n_40),
.B2(n_34),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_318),
.A2(n_271),
.B1(n_40),
.B2(n_34),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_262),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_286),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_321),
.A2(n_329),
.B1(n_330),
.B2(n_339),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_324),
.B(n_328),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_325),
.A2(n_331),
.B(n_317),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_345),
.Y(n_350)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_277),
.B(n_268),
.C(n_282),
.D(n_290),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_304),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_333),
.B(n_337),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_334),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_183),
.Y(n_337)
);

NOR3xp33_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_33),
.C(n_56),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_343),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_291),
.A2(n_307),
.B1(n_297),
.B2(n_311),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_291),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_341)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_341),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_10),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_342),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_346),
.Y(n_363)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_298),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_292),
.C(n_306),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_365),
.C(n_368),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_349),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_336),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_320),
.B(n_293),
.C(n_295),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_361),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_309),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_322),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_327),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_322),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_335),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_320),
.C(n_294),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_297),
.B1(n_299),
.B2(n_294),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_366),
.A2(n_370),
.B1(n_327),
.B2(n_338),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_313),
.C(n_310),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_369),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_332),
.A2(n_300),
.B1(n_314),
.B2(n_318),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_343),
.A2(n_314),
.B1(n_296),
.B2(n_27),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_344),
.B1(n_331),
.B2(n_335),
.Y(n_376)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_373),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_340),
.B(n_0),
.Y(n_374)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_374),
.Y(n_384)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_375),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_391),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_385),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_325),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_394),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_367),
.Y(n_386)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_368),
.A2(n_328),
.B(n_340),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_387),
.A2(n_352),
.B(n_362),
.Y(n_400)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_360),
.C(n_365),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_390),
.C(n_363),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_369),
.B(n_329),
.C(n_323),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_372),
.A2(n_321),
.B1(n_323),
.B2(n_341),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_392),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_395),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_366),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_334),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_358),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_408),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_400),
.A2(n_393),
.B(n_354),
.Y(n_423)
);

AOI321xp33_ASAP7_75t_L g402 ( 
.A1(n_378),
.A2(n_363),
.A3(n_353),
.B1(n_374),
.B2(n_373),
.C(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_402),
.Y(n_424)
);

BUFx24_ASAP7_75t_SL g403 ( 
.A(n_395),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_403),
.B(n_410),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_385),
.Y(n_414)
);

A2O1A1O1Ixp25_ASAP7_75t_L g408 ( 
.A1(n_378),
.A2(n_353),
.B(n_361),
.C(n_357),
.D(n_359),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_392),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_412),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_384),
.A2(n_359),
.B1(n_370),
.B2(n_361),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_390),
.A2(n_380),
.B1(n_394),
.B2(n_381),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_407),
.A2(n_380),
.B1(n_382),
.B2(n_379),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_413),
.A2(n_419),
.B1(n_427),
.B2(n_412),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_5),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_398),
.A2(n_387),
.B(n_381),
.Y(n_415)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_389),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_422),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_397),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_425),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_402),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_377),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_411),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_351),
.C(n_2),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_9),
.Y(n_426)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_426),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_408),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_424),
.A2(n_406),
.B1(n_405),
.B2(n_401),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_434),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_416),
.A2(n_401),
.B(n_411),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_435),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_431),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_432),
.A2(n_415),
.B1(n_420),
.B2(n_421),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_9),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_433),
.A2(n_425),
.B(n_423),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_420),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_427),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_441),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_428),
.B(n_414),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_437),
.B(n_417),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_422),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_444),
.B(n_5),
.C(n_11),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_446),
.A2(n_447),
.B1(n_448),
.B2(n_438),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_432),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_445),
.A2(n_433),
.B1(n_436),
.B2(n_438),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_450),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_451),
.A2(n_453),
.B(n_448),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_443),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_444),
.B(n_12),
.C(n_3),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_456),
.B(n_457),
.Y(n_459)
);

AOI322xp5_ASAP7_75t_L g458 ( 
.A1(n_455),
.A2(n_454),
.A3(n_441),
.B1(n_440),
.B2(n_443),
.C1(n_452),
.C2(n_453),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g460 ( 
.A1(n_458),
.A2(n_0),
.B(n_3),
.Y(n_460)
);

AOI322xp5_ASAP7_75t_L g461 ( 
.A1(n_460),
.A2(n_0),
.A3(n_3),
.B1(n_4),
.B2(n_103),
.C1(n_459),
.C2(n_312),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_0),
.Y(n_462)
);

BUFx24_ASAP7_75t_SL g463 ( 
.A(n_462),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_463),
.A2(n_4),
.B(n_103),
.Y(n_464)
);


endmodule