module fake_jpeg_18362_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_56),
.Y(n_64)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_48),
.B1(n_42),
.B2(n_38),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_48),
.B1(n_42),
.B2(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_49),
.B1(n_39),
.B2(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_82),
.B1(n_85),
.B2(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_60),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_83),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_3),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_49),
.B(n_50),
.C(n_21),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_14),
.B(n_27),
.C(n_26),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_61),
.B1(n_20),
.B2(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_16),
.B1(n_33),
.B2(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_83),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_15),
.B1(n_30),
.B2(n_28),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_92),
.B1(n_77),
.B2(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_80),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_35),
.CON(n_94),
.SN(n_94)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_82),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_89),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_100),
.B1(n_96),
.B2(n_99),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_101),
.B1(n_102),
.B2(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_92),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_94),
.B(n_92),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_95),
.B1(n_93),
.B2(n_13),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_10),
.B(n_11),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_19),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_24),
.B(n_25),
.Y(n_111)
);


endmodule