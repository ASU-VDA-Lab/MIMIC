module fake_jpeg_20223_n_215 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx2_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_14),
.B1(n_24),
.B2(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_15),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_15),
.B(n_29),
.C(n_21),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_44),
.A2(n_5),
.B(n_6),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_29),
.B1(n_21),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_2),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_31),
.A2(n_24),
.B1(n_14),
.B2(n_27),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_30),
.B1(n_3),
.B2(n_4),
.Y(n_77)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_15),
.B1(n_27),
.B2(n_23),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_45),
.B1(n_56),
.B2(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_69),
.B(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_22),
.B1(n_20),
.B2(n_13),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_16),
.B(n_25),
.C(n_22),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_20),
.B1(n_13),
.B2(n_25),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_85),
.B1(n_51),
.B2(n_63),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_30),
.C(n_4),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_83),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_5),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_93),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_7),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_63),
.Y(n_108)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_91),
.Y(n_107)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_7),
.B(n_8),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_8),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_95),
.C(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_10),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_11),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_62),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_114),
.B1(n_119),
.B2(n_85),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_113),
.B(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_72),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_123),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_55),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_62),
.B1(n_81),
.B2(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_144),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_76),
.B1(n_91),
.B2(n_98),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_100),
.B1(n_116),
.B2(n_76),
.Y(n_150)
);

BUFx12f_ASAP7_75t_SL g142 ( 
.A(n_99),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_113),
.B(n_107),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_76),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_67),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_67),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_156),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_161),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_133),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_116),
.B(n_113),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_159),
.B(n_133),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_105),
.B1(n_122),
.B2(n_102),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_124),
.C(n_104),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_145),
.C(n_138),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_142),
.B(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_174),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_155),
.B(n_147),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_170),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_166),
.B(n_176),
.Y(n_186)
);

AOI22x1_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_177),
.B1(n_149),
.B2(n_151),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_162),
.C(n_157),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_172),
.A2(n_178),
.B1(n_149),
.B2(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

AO221x1_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_146),
.B1(n_117),
.B2(n_128),
.C(n_135),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_148),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_132),
.C(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_182),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_153),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_189),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_169),
.B(n_186),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_160),
.C(n_130),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_165),
.C(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_140),
.B1(n_163),
.B2(n_139),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_175),
.B(n_168),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_197),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_187),
.A2(n_164),
.B(n_154),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_184),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_178),
.B(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_181),
.B1(n_179),
.B2(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_193),
.A2(n_131),
.B1(n_125),
.B2(n_120),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_194),
.A3(n_196),
.B1(n_139),
.B2(n_130),
.C1(n_136),
.C2(n_104),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_146),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_SL g210 ( 
.A(n_204),
.B(n_207),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_202),
.A2(n_196),
.B(n_102),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_199),
.B(n_198),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_200),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_209),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_206),
.B1(n_110),
.B2(n_89),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_212),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_75),
.B(n_110),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_90),
.Y(n_215)
);


endmodule