module fake_jpeg_7614_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_29),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_35),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx2_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_67),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_20),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_36),
.B(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_70),
.B(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_47),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_20),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_94),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_91),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_90),
.B1(n_95),
.B2(n_35),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_42),
.B1(n_33),
.B2(n_26),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_21),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_33),
.B1(n_26),
.B2(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_65),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_41),
.C(n_40),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_42),
.B1(n_64),
.B2(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_83),
.B1(n_80),
.B2(n_84),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_121),
.B1(n_124),
.B2(n_77),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_18),
.B1(n_55),
.B2(n_54),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_46),
.Y(n_147)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_126),
.B1(n_73),
.B2(n_92),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_64),
.B1(n_60),
.B2(n_54),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_78),
.B1(n_79),
.B2(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_55),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_60),
.B1(n_61),
.B2(n_25),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_52),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_72),
.A2(n_61),
.B1(n_32),
.B2(n_25),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

BUFx24_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_133),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_74),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_155),
.C(n_46),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_140),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_139),
.B1(n_113),
.B2(n_115),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_91),
.B(n_85),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_107),
.A3(n_19),
.B1(n_24),
.B2(n_46),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_81),
.B1(n_84),
.B2(n_98),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_142),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_28),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_83),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_110),
.A2(n_80),
.B1(n_32),
.B2(n_22),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_151),
.B1(n_153),
.B2(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_30),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_127),
.B1(n_112),
.B2(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_47),
.B1(n_45),
.B2(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_30),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_41),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_165),
.C(n_181),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_154),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_184),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_129),
.B(n_144),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_160),
.A2(n_166),
.B(n_164),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_152),
.B1(n_134),
.B2(n_140),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_130),
.B1(n_34),
.B2(n_31),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_125),
.B1(n_104),
.B2(n_107),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_167),
.B1(n_172),
.B2(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_104),
.B1(n_123),
.B2(n_103),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_103),
.B1(n_93),
.B2(n_99),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_14),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_141),
.B(n_153),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_182),
.B(n_147),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_45),
.B1(n_99),
.B2(n_117),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_46),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_75),
.B(n_19),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_24),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_0),
.C(n_1),
.Y(n_213)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_16),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_205),
.B(n_211),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_196),
.B1(n_198),
.B2(n_201),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_139),
.B1(n_148),
.B2(n_133),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_189),
.A2(n_194),
.B1(n_200),
.B2(n_170),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_142),
.B1(n_130),
.B2(n_117),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_168),
.B1(n_182),
.B2(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_199),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_183),
.A3(n_161),
.B1(n_177),
.B2(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_142),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_203),
.C(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_130),
.B1(n_34),
.B2(n_31),
.Y(n_194)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_180),
.B1(n_159),
.B2(n_158),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_19),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_24),
.Y(n_204)
);

AND2x4_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_34),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_31),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_207),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_22),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_213),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_30),
.B1(n_16),
.B2(n_15),
.Y(n_209)
);

OAI22x1_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_185),
.B1(n_175),
.B2(n_161),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_186),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_197),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_223),
.Y(n_249)
);

BUFx8_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_221),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_222),
.A2(n_230),
.B1(n_233),
.B2(n_239),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_229),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_187),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_227),
.B(n_234),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_229),
.B(n_238),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_168),
.B1(n_172),
.B2(n_170),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_191),
.B1(n_190),
.B2(n_192),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_197),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_189),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_206),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_207),
.B(n_184),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_213),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_210),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_214),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_194),
.B1(n_5),
.B2(n_6),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_261),
.B(n_223),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_195),
.C(n_193),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_258),
.C(n_263),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_253),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_195),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_203),
.C(n_204),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_15),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_241),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_260),
.A2(n_231),
.B1(n_222),
.B2(n_219),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_215),
.A2(n_4),
.B(n_5),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_218),
.B(n_6),
.C(n_7),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_270),
.B(n_262),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_224),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_216),
.B1(n_225),
.B2(n_233),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_273),
.B1(n_249),
.B2(n_264),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_251),
.B1(n_250),
.B2(n_257),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_215),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_279),
.C(n_281),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_259),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_225),
.C(n_226),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_245),
.B(n_264),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_247),
.B(n_230),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_284),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_290),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_281),
.C(n_7),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_243),
.B(n_245),
.Y(n_288)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_270),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_224),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_292),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_242),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_217),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_277),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_263),
.C(n_255),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_296),
.C(n_283),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_254),
.B1(n_240),
.B2(n_261),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_295),
.A2(n_278),
.B1(n_282),
.B2(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_221),
.C(n_256),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_221),
.B(n_7),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_297),
.A2(n_286),
.B(n_287),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_306),
.C(n_308),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_302),
.B1(n_303),
.B2(n_6),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_309),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_275),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_267),
.C(n_269),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_297),
.B(n_295),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_310),
.B(n_306),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_304),
.B(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_317),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_290),
.C(n_284),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_315),
.A2(n_318),
.B(n_319),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_285),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_10),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_8),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_8),
.B(n_9),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_8),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_10),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_300),
.B1(n_11),
.B2(n_12),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_316),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_312),
.A2(n_10),
.B(n_11),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_328),
.A2(n_11),
.B(n_12),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_330),
.A2(n_331),
.B(n_322),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_327),
.C(n_321),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_334),
.B(n_326),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_329),
.C(n_12),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_13),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_13),
.B(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_13),
.Y(n_339)
);


endmodule