module fake_netlist_1_8024_n_33 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_10), .B(n_0), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_12), .Y(n_17) );
O2A1O1Ixp33_ASAP7_75t_L g18 ( .A1(n_11), .A2(n_13), .B(n_9), .C(n_10), .Y(n_18) );
O2A1O1Ixp33_ASAP7_75t_L g19 ( .A1(n_14), .A2(n_1), .B(n_4), .C(n_5), .Y(n_19) );
NOR2xp33_ASAP7_75t_SL g20 ( .A(n_19), .B(n_14), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_17), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_21), .Y(n_24) );
INVx1_ASAP7_75t_SL g25 ( .A(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_22), .B1(n_20), .B2(n_12), .Y(n_27) );
OAI221xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_20), .B1(n_24), .B2(n_23), .C(n_25), .Y(n_28) );
O2A1O1Ixp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_18), .B(n_16), .C(n_25), .Y(n_29) );
INVx2_ASAP7_75t_SL g30 ( .A(n_29), .Y(n_30) );
INVx5_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_31), .B1(n_15), .B2(n_7), .Y(n_33) );
endmodule