module real_aes_2766_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_0), .B(n_152), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_1), .A2(n_134), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_2), .B(n_111), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_3), .A2(n_11), .B1(n_815), .B2(n_816), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_3), .Y(n_816) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_4), .B(n_142), .Y(n_198) );
INVx1_ASAP7_75t_L g139 ( .A(n_5), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_6), .B(n_142), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_7), .B(n_129), .Y(n_475) );
INVx1_ASAP7_75t_L g503 ( .A(n_8), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_9), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_10), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_11), .Y(n_815) );
NAND2xp33_ASAP7_75t_L g179 ( .A(n_12), .B(n_146), .Y(n_179) );
INVx2_ASAP7_75t_L g131 ( .A(n_13), .Y(n_131) );
AOI221x1_ASAP7_75t_L g221 ( .A1(n_14), .A2(n_26), .B1(n_134), .B2(n_152), .C(n_222), .Y(n_221) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_15), .B(n_110), .C(n_112), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g442 ( .A(n_15), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_16), .B(n_152), .Y(n_175) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_17), .A2(n_173), .B(n_174), .Y(n_172) );
INVx1_ASAP7_75t_L g484 ( .A(n_18), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_19), .B(n_165), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_20), .B(n_142), .Y(n_141) );
AO21x1_ASAP7_75t_L g193 ( .A1(n_21), .A2(n_152), .B(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g108 ( .A(n_22), .Y(n_108) );
INVx1_ASAP7_75t_L g482 ( .A(n_23), .Y(n_482) );
INVx1_ASAP7_75t_SL g468 ( .A(n_24), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_25), .B(n_153), .Y(n_562) );
NAND2x1_ASAP7_75t_L g207 ( .A(n_27), .B(n_142), .Y(n_207) );
AOI33xp33_ASAP7_75t_L g530 ( .A1(n_28), .A2(n_53), .A3(n_458), .B1(n_465), .B2(n_531), .B3(n_532), .Y(n_530) );
NAND2x1_ASAP7_75t_L g161 ( .A(n_29), .B(n_146), .Y(n_161) );
INVx1_ASAP7_75t_L g512 ( .A(n_30), .Y(n_512) );
OR2x2_ASAP7_75t_L g130 ( .A(n_31), .B(n_86), .Y(n_130) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_31), .A2(n_86), .B(n_131), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_32), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_33), .B(n_146), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_34), .B(n_142), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_35), .B(n_146), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_36), .A2(n_134), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g135 ( .A(n_37), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g150 ( .A(n_37), .B(n_139), .Y(n_150) );
INVx1_ASAP7_75t_L g464 ( .A(n_37), .Y(n_464) );
INVxp67_ASAP7_75t_L g112 ( .A(n_38), .Y(n_112) );
OR2x6_ASAP7_75t_L g443 ( .A(n_38), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_39), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_40), .B(n_152), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_41), .B(n_456), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_42), .A2(n_129), .B1(n_169), .B2(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_43), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_44), .B(n_153), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_45), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_46), .B(n_146), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_47), .B(n_173), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_48), .B(n_153), .Y(n_504) );
INVxp33_ASAP7_75t_L g821 ( .A(n_49), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_50), .A2(n_134), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_51), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_52), .B(n_146), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_54), .B(n_153), .Y(n_542) );
INVx1_ASAP7_75t_L g138 ( .A(n_55), .Y(n_138) );
INVx1_ASAP7_75t_L g148 ( .A(n_55), .Y(n_148) );
AND2x2_ASAP7_75t_L g543 ( .A(n_56), .B(n_165), .Y(n_543) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_57), .A2(n_75), .B1(n_456), .B2(n_462), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_58), .B(n_456), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_59), .B(n_142), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_60), .B(n_169), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_61), .Y(n_806) );
AOI21xp5_ASAP7_75t_SL g492 ( .A1(n_62), .A2(n_462), .B(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_63), .A2(n_134), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g478 ( .A(n_64), .Y(n_478) );
AO21x1_ASAP7_75t_L g195 ( .A1(n_65), .A2(n_134), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_66), .B(n_152), .Y(n_183) );
INVx1_ASAP7_75t_L g541 ( .A(n_67), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_68), .B(n_152), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_69), .A2(n_462), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g244 ( .A(n_70), .B(n_166), .Y(n_244) );
INVx1_ASAP7_75t_L g136 ( .A(n_71), .Y(n_136) );
INVx1_ASAP7_75t_L g144 ( .A(n_71), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_72), .A2(n_97), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_72), .Y(n_116) );
AND2x2_ASAP7_75t_L g167 ( .A(n_73), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_74), .B(n_456), .Y(n_533) );
AND2x2_ASAP7_75t_L g471 ( .A(n_76), .B(n_168), .Y(n_471) );
INVx1_ASAP7_75t_L g479 ( .A(n_77), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_78), .A2(n_462), .B(n_467), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_79), .A2(n_462), .B(n_525), .C(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_80), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g445 ( .A(n_80), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_81), .B(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g181 ( .A(n_82), .B(n_168), .Y(n_181) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_83), .B(n_168), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_84), .A2(n_462), .B1(n_528), .B2(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g194 ( .A(n_85), .B(n_129), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_87), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g211 ( .A(n_88), .B(n_168), .Y(n_211) );
INVx1_ASAP7_75t_L g494 ( .A(n_89), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_90), .A2(n_115), .B1(n_787), .B2(n_791), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_91), .B(n_142), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_92), .A2(n_134), .B(n_140), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_93), .B(n_146), .Y(n_223) );
AND2x2_ASAP7_75t_L g534 ( .A(n_94), .B(n_168), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_95), .B(n_142), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_96), .A2(n_510), .B(n_511), .C(n_513), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_97), .Y(n_117) );
BUFx2_ASAP7_75t_L g798 ( .A(n_98), .Y(n_798) );
BUFx2_ASAP7_75t_SL g811 ( .A(n_98), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_99), .A2(n_134), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_100), .B(n_153), .Y(n_495) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_113), .B(n_820), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g822 ( .A(n_105), .Y(n_822) );
INVx3_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_109), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_108), .B(n_445), .Y(n_444) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_795), .B(n_807), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B(n_786), .Y(n_114) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_438), .B1(n_446), .B2(n_784), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g813 ( .A1(n_120), .A2(n_121), .B1(n_814), .B2(n_817), .Y(n_813) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_121), .A2(n_447), .B1(n_788), .B2(n_789), .Y(n_787) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_336), .Y(n_121) );
NAND3xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_248), .C(n_303), .Y(n_122) );
AOI221xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_188), .B1(n_212), .B2(n_216), .C(n_226), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_171), .Y(n_124) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_125), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g247 ( .A(n_125), .Y(n_247) );
AND2x2_ASAP7_75t_L g292 ( .A(n_125), .B(n_229), .Y(n_292) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_156), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g280 ( .A(n_127), .Y(n_280) );
INVx1_ASAP7_75t_L g290 ( .A(n_127), .Y(n_290) );
AO21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B(n_154), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_128), .B(n_155), .Y(n_154) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_128), .A2(n_132), .B(n_154), .Y(n_254) );
INVx1_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_129), .A2(n_175), .B(n_176), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_129), .B(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_129), .B(n_149), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_129), .A2(n_492), .B(n_496), .Y(n_491) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_130), .B(n_131), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_151), .Y(n_132) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
BUFx3_ASAP7_75t_L g460 ( .A(n_135), .Y(n_460) );
AND2x6_ASAP7_75t_L g146 ( .A(n_136), .B(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g466 ( .A(n_136), .Y(n_466) );
AND2x4_ASAP7_75t_L g462 ( .A(n_137), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x4_ASAP7_75t_L g142 ( .A(n_138), .B(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g458 ( .A(n_138), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_139), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B(n_149), .Y(n_140) );
INVxp67_ASAP7_75t_L g485 ( .A(n_142), .Y(n_485) );
AND2x4_ASAP7_75t_L g153 ( .A(n_143), .B(n_147), .Y(n_153) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVxp67_ASAP7_75t_L g483 ( .A(n_146), .Y(n_483) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_149), .A2(n_161), .B(n_162), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_149), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_149), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_149), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_149), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_149), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_149), .A2(n_241), .B(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g467 ( .A1(n_149), .A2(n_468), .B(n_469), .C(n_470), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_149), .A2(n_469), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_149), .A2(n_469), .B(n_503), .C(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g528 ( .A(n_149), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_149), .A2(n_469), .B(n_541), .C(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_149), .A2(n_562), .B(n_563), .Y(n_561) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g152 ( .A(n_150), .B(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_150), .Y(n_513) );
INVx1_ASAP7_75t_L g480 ( .A(n_153), .Y(n_480) );
OR2x2_ASAP7_75t_L g269 ( .A(n_156), .B(n_172), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_156), .B(n_215), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_156), .B(n_180), .Y(n_313) );
INVx2_ASAP7_75t_L g322 ( .A(n_156), .Y(n_322) );
AND2x2_ASAP7_75t_L g343 ( .A(n_156), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g427 ( .A(n_156), .B(n_246), .Y(n_427) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g255 ( .A(n_157), .B(n_180), .Y(n_255) );
AND2x2_ASAP7_75t_L g388 ( .A(n_157), .B(n_215), .Y(n_388) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_157), .Y(n_414) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_164), .B(n_167), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_163), .Y(n_158) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_164), .A2(n_454), .B(n_471), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_165), .A2(n_183), .B(n_184), .Y(n_182) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_165), .A2(n_221), .B(n_225), .Y(n_220) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_165), .A2(n_221), .B(n_225), .Y(n_232) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx3_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_168), .A2(n_210), .B1(n_509), .B2(n_514), .Y(n_508) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_169), .B(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx4f_ASAP7_75t_L g173 ( .A(n_170), .Y(n_173) );
AND2x4_ASAP7_75t_L g342 ( .A(n_171), .B(n_343), .Y(n_342) );
AOI321xp33_ASAP7_75t_L g356 ( .A1(n_171), .A2(n_285), .A3(n_286), .B1(n_318), .B2(n_357), .C(n_360), .Y(n_356) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_180), .Y(n_171) );
BUFx3_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
INVx2_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_172), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g279 ( .A(n_172), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g312 ( .A(n_172), .Y(n_312) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_173), .A2(n_501), .B(n_505), .Y(n_500) );
INVx2_ASAP7_75t_SL g525 ( .A(n_173), .Y(n_525) );
INVx5_ASAP7_75t_L g215 ( .A(n_180), .Y(n_215) );
NOR2x1_ASAP7_75t_SL g264 ( .A(n_180), .B(n_254), .Y(n_264) );
BUFx2_ASAP7_75t_L g359 ( .A(n_180), .Y(n_359) );
OR2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVxp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_201), .Y(n_189) );
NOR2xp33_ASAP7_75t_SL g257 ( .A(n_190), .B(n_258), .Y(n_257) );
NOR4xp25_ASAP7_75t_L g360 ( .A(n_190), .B(n_354), .C(n_358), .D(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g398 ( .A(n_190), .Y(n_398) );
AND2x2_ASAP7_75t_L g432 ( .A(n_190), .B(n_372), .Y(n_432) );
BUFx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g233 ( .A(n_191), .Y(n_233) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g287 ( .A(n_192), .Y(n_287) );
OAI21x1_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_195), .B(n_199), .Y(n_192) );
INVx1_ASAP7_75t_L g200 ( .A(n_194), .Y(n_200) );
AOI33xp33_ASAP7_75t_L g428 ( .A1(n_201), .A2(n_230), .A3(n_261), .B1(n_277), .B2(n_383), .B3(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g218 ( .A(n_202), .B(n_219), .Y(n_218) );
AND2x4_ASAP7_75t_L g228 ( .A(n_202), .B(n_229), .Y(n_228) );
BUFx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g235 ( .A(n_203), .Y(n_235) );
INVxp67_ASAP7_75t_L g316 ( .A(n_203), .Y(n_316) );
AND2x2_ASAP7_75t_L g372 ( .A(n_203), .B(n_237), .Y(n_372) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_203) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_210), .A2(n_238), .B(n_244), .Y(n_237) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_210), .A2(n_238), .B(n_244), .Y(n_273) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_210), .A2(n_537), .B(n_543), .Y(n_536) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_210), .A2(n_537), .B(n_543), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_212), .A2(n_394), .B(n_395), .Y(n_393) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g381 ( .A(n_213), .B(n_255), .Y(n_381) );
AND3x2_ASAP7_75t_L g383 ( .A(n_213), .B(n_267), .C(n_322), .Y(n_383) );
INVx3_ASAP7_75t_SL g335 ( .A(n_214), .Y(n_335) );
INVx4_ASAP7_75t_L g229 ( .A(n_215), .Y(n_229) );
AND2x2_ASAP7_75t_L g267 ( .A(n_215), .B(n_254), .Y(n_267) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g261 ( .A(n_219), .Y(n_261) );
AND2x4_ASAP7_75t_L g286 ( .A(n_219), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g349 ( .A(n_219), .B(n_237), .Y(n_349) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g319 ( .A(n_220), .Y(n_319) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_220), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_R g226 ( .A1(n_227), .A2(n_230), .B(n_234), .C(n_245), .Y(n_226) );
CKINVDCx16_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g278 ( .A(n_229), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_229), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_229), .B(n_246), .Y(n_407) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g389 ( .A(n_231), .B(n_379), .Y(n_389) );
AND2x2_ASAP7_75t_SL g231 ( .A(n_232), .B(n_233), .Y(n_231) );
AND2x2_ASAP7_75t_L g236 ( .A(n_232), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g258 ( .A(n_232), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g274 ( .A(n_232), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g307 ( .A(n_232), .B(n_287), .Y(n_307) );
AND2x4_ASAP7_75t_L g272 ( .A(n_233), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g296 ( .A(n_233), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g334 ( .A(n_233), .B(n_259), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g262 ( .A(n_235), .B(n_259), .Y(n_262) );
AND2x2_ASAP7_75t_L g277 ( .A(n_235), .B(n_237), .Y(n_277) );
BUFx2_ASAP7_75t_L g333 ( .A(n_235), .Y(n_333) );
AND2x2_ASAP7_75t_L g347 ( .A(n_235), .B(n_258), .Y(n_347) );
INVx2_ASAP7_75t_L g259 ( .A(n_237), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_239), .B(n_243), .Y(n_238) );
OAI22xp33_ASAP7_75t_L g295 ( .A1(n_245), .A2(n_296), .B1(n_298), .B2(n_302), .Y(n_295) );
INVx2_ASAP7_75t_SL g326 ( .A(n_245), .Y(n_326) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g301 ( .A(n_246), .B(n_254), .Y(n_301) );
INVx1_ASAP7_75t_L g408 ( .A(n_247), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_281), .C(n_295), .Y(n_248) );
OAI221xp5_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_256), .B1(n_260), .B2(n_263), .C(n_265), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVxp67_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g309 ( .A(n_253), .Y(n_309) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_253), .Y(n_437) );
INVx1_ASAP7_75t_L g400 ( .A(n_255), .Y(n_400) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_255), .B(n_279), .Y(n_410) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_259), .B(n_287), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OR2x2_ASAP7_75t_L g293 ( .A(n_261), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g371 ( .A(n_261), .Y(n_371) );
AND2x2_ASAP7_75t_L g306 ( .A(n_262), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g352 ( .A(n_264), .B(n_312), .Y(n_352) );
AND2x2_ASAP7_75t_L g429 ( .A(n_264), .B(n_427), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_270), .B1(n_277), .B2(n_278), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g288 ( .A(n_269), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx2_ASAP7_75t_L g294 ( .A(n_272), .Y(n_294) );
AND2x4_ASAP7_75t_L g318 ( .A(n_272), .B(n_319), .Y(n_318) );
OAI21xp33_ASAP7_75t_SL g348 ( .A1(n_272), .A2(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g375 ( .A(n_272), .B(n_333), .Y(n_375) );
INVx2_ASAP7_75t_L g297 ( .A(n_273), .Y(n_297) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
INVx1_ASAP7_75t_SL g354 ( .A(n_274), .Y(n_354) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx2_ASAP7_75t_L g285 ( .A(n_276), .Y(n_285) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_276), .B(n_297), .Y(n_379) );
AND2x2_ASAP7_75t_L g376 ( .A(n_279), .B(n_322), .Y(n_376) );
AND2x2_ASAP7_75t_L g402 ( .A(n_279), .B(n_388), .Y(n_402) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_280), .Y(n_324) );
INVx1_ASAP7_75t_L g344 ( .A(n_280), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_288), .B1(n_291), .B2(n_293), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_286), .B(n_297), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_286), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g425 ( .A(n_286), .Y(n_425) );
INVx2_ASAP7_75t_SL g350 ( .A(n_288), .Y(n_350) );
AND2x2_ASAP7_75t_L g362 ( .A(n_290), .B(n_322), .Y(n_362) );
INVx2_ASAP7_75t_L g368 ( .A(n_290), .Y(n_368) );
INVxp33_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g327 ( .A(n_293), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_296), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g418 ( .A(n_296), .Y(n_418) );
INVx1_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_299), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g357 ( .A(n_301), .B(n_358), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_301), .A2(n_431), .B1(n_432), .B2(n_433), .Y(n_430) );
NOR3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_325), .C(n_328), .Y(n_303) );
OAI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_308), .B1(n_310), .B2(n_314), .C(n_317), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g423 ( .A(n_308), .Y(n_423) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g392 ( .A(n_309), .B(n_358), .Y(n_392) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g323 ( .A(n_312), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g394 ( .A(n_314), .Y(n_394) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g391 ( .A(n_315), .Y(n_391) );
INVx1_ASAP7_75t_L g397 ( .A(n_316), .Y(n_397) );
OR2x2_ASAP7_75t_L g420 ( .A(n_316), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_SL g329 ( .A(n_319), .Y(n_329) );
AND2x2_ASAP7_75t_L g399 ( .A(n_319), .B(n_379), .Y(n_399) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_319), .B(n_332), .Y(n_431) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g436 ( .A(n_322), .Y(n_436) );
INVx1_ASAP7_75t_L g386 ( .A(n_324), .Y(n_386) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B(n_331), .C(n_335), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_329), .B(n_379), .Y(n_403) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_332), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AND2x2_ASAP7_75t_L g340 ( .A(n_334), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g421 ( .A(n_334), .Y(n_421) );
NAND4xp75_ASAP7_75t_L g336 ( .A(n_337), .B(n_393), .C(n_409), .D(n_430), .Y(n_336) );
NOR3x1_ASAP7_75t_L g337 ( .A(n_338), .B(n_355), .C(n_377), .Y(n_337) );
NAND4xp75_ASAP7_75t_L g338 ( .A(n_339), .B(n_345), .C(n_348), .D(n_351), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_340), .B(n_342), .Y(n_339) );
AND2x2_ASAP7_75t_L g390 ( .A(n_341), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g415 ( .A(n_342), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_SL g404 ( .A(n_347), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_363), .Y(n_355) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_359), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_369), .B(n_373), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI322xp33_ASAP7_75t_L g395 ( .A1(n_367), .A2(n_396), .A3(n_400), .B1(n_401), .B2(n_403), .C1(n_404), .C2(n_405), .Y(n_395) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_368), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_371), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_372), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_382), .C(n_384), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .B1(n_390), .B2(n_392), .Y(n_384) );
NOR2xp33_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .Y(n_385) );
INVx2_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_399), .Y(n_396) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_402), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_406), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g412 ( .A(n_407), .B(n_413), .Y(n_412) );
O2A1O1Ixp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_416), .C(n_419), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_422), .B1(n_424), .B2(n_426), .C(n_428), .Y(n_419) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx4_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
CKINVDCx6p67_ASAP7_75t_R g788 ( .A(n_439), .Y(n_788) );
INVx3_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
AND2x6_ASAP7_75t_SL g441 ( .A(n_442), .B(n_443), .Y(n_441) );
OR2x6_ASAP7_75t_SL g784 ( .A(n_442), .B(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g794 ( .A(n_442), .B(n_443), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_442), .B(n_785), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_443), .Y(n_785) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR3x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_649), .C(n_720), .Y(n_447) );
NAND3x1_ASAP7_75t_SL g448 ( .A(n_449), .B(n_576), .C(n_598), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_566), .Y(n_449) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_497), .B1(n_544), .B2(n_548), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_451), .A2(n_752), .B1(n_753), .B2(n_755), .Y(n_751) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_472), .Y(n_451) );
AND2x2_ASAP7_75t_L g567 ( .A(n_452), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_452), .B(n_614), .Y(n_633) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g551 ( .A(n_453), .Y(n_551) );
AND2x2_ASAP7_75t_L g601 ( .A(n_453), .B(n_474), .Y(n_601) );
INVx1_ASAP7_75t_L g640 ( .A(n_453), .Y(n_640) );
OR2x2_ASAP7_75t_L g677 ( .A(n_453), .B(n_489), .Y(n_677) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_453), .Y(n_689) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_453), .Y(n_713) );
AND2x2_ASAP7_75t_L g770 ( .A(n_453), .B(n_597), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_461), .Y(n_454) );
INVx1_ASAP7_75t_L g521 ( .A(n_456), .Y(n_521) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_460), .Y(n_456) );
INVx1_ASAP7_75t_L g557 ( .A(n_457), .Y(n_557) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OR2x6_ASAP7_75t_L g469 ( .A(n_458), .B(n_466), .Y(n_469) );
INVxp33_ASAP7_75t_L g531 ( .A(n_458), .Y(n_531) );
INVx1_ASAP7_75t_L g558 ( .A(n_460), .Y(n_558) );
INVxp67_ASAP7_75t_L g519 ( .A(n_462), .Y(n_519) );
NOR2x1p5_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_469), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_477) );
INVxp67_ASAP7_75t_L g510 ( .A(n_469), .Y(n_510) );
INVx2_ASAP7_75t_L g564 ( .A(n_469), .Y(n_564) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_487), .Y(n_472) );
INVx1_ASAP7_75t_L g645 ( .A(n_473), .Y(n_645) );
AND2x2_ASAP7_75t_L g671 ( .A(n_473), .B(n_489), .Y(n_671) );
NAND2x1_ASAP7_75t_L g687 ( .A(n_473), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g568 ( .A(n_474), .B(n_554), .Y(n_568) );
INVx3_ASAP7_75t_L g597 ( .A(n_474), .Y(n_597) );
NOR2x1_ASAP7_75t_SL g716 ( .A(n_474), .B(n_489), .Y(n_716) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_481), .B(n_486), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_480), .B(n_512), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_484), .B2(n_485), .Y(n_481) );
NOR2x1_ASAP7_75t_L g624 ( .A(n_487), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g595 ( .A(n_488), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx4_ASAP7_75t_L g565 ( .A(n_489), .Y(n_565) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_489), .Y(n_610) );
AND2x2_ASAP7_75t_L g682 ( .A(n_489), .B(n_554), .Y(n_682) );
AND2x4_ASAP7_75t_L g699 ( .A(n_489), .B(n_643), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_489), .B(n_641), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_489), .B(n_550), .Y(n_775) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_497), .A2(n_592), .B1(n_663), .B2(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_522), .Y(n_497) );
INVx2_ASAP7_75t_L g665 ( .A(n_498), .Y(n_665) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_506), .Y(n_498) );
BUFx3_ASAP7_75t_L g655 ( .A(n_499), .Y(n_655) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_500), .B(n_524), .Y(n_547) );
INVx2_ASAP7_75t_L g571 ( .A(n_500), .Y(n_571) );
INVx1_ASAP7_75t_L g583 ( .A(n_500), .Y(n_583) );
AND2x4_ASAP7_75t_L g590 ( .A(n_500), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g607 ( .A(n_500), .B(n_507), .Y(n_607) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_500), .Y(n_621) );
INVxp67_ASAP7_75t_L g629 ( .A(n_500), .Y(n_629) );
AND2x2_ASAP7_75t_L g658 ( .A(n_506), .B(n_574), .Y(n_658) );
AND2x2_ASAP7_75t_L g674 ( .A(n_506), .B(n_575), .Y(n_674) );
NOR2xp67_ASAP7_75t_L g761 ( .A(n_506), .B(n_574), .Y(n_761) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g570 ( .A(n_507), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g581 ( .A(n_507), .Y(n_581) );
INVx1_ASAP7_75t_L g594 ( .A(n_507), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_507), .B(n_536), .Y(n_631) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_515), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_519), .B1(n_520), .B2(n_521), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g754 ( .A(n_522), .Y(n_754) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_535), .Y(n_522) );
AND2x2_ASAP7_75t_L g628 ( .A(n_523), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g657 ( .A(n_523), .Y(n_657) );
AND2x2_ASAP7_75t_L g759 ( .A(n_523), .B(n_574), .Y(n_759) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_524), .B(n_536), .Y(n_619) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B(n_534), .Y(n_524) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_525), .A2(n_526), .B(n_534), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_527), .B(n_533), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_L g545 ( .A(n_535), .Y(n_545) );
NAND2x1p5_ASAP7_75t_L g734 ( .A(n_535), .B(n_655), .Y(n_734) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_536), .Y(n_648) );
AND2x2_ASAP7_75t_L g675 ( .A(n_536), .B(n_621), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AND2x2_ASAP7_75t_L g589 ( .A(n_545), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g605 ( .A(n_545), .Y(n_605) );
AND2x2_ASAP7_75t_L g693 ( .A(n_545), .B(n_570), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_545), .B(n_713), .Y(n_718) );
AND2x2_ASAP7_75t_L g728 ( .A(n_545), .B(n_607), .Y(n_728) );
OR2x2_ASAP7_75t_L g765 ( .A(n_545), .B(n_665), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_546), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g725 ( .A(n_546), .B(n_581), .Y(n_725) );
AND2x2_ASAP7_75t_L g741 ( .A(n_546), .B(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g735 ( .A(n_547), .B(n_631), .Y(n_735) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_L g617 ( .A(n_549), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_549), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g715 ( .A(n_549), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_549), .B(n_596), .Y(n_740) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_550), .Y(n_587) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_551), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_552), .A2(n_585), .B1(n_603), .B2(n_606), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_552), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_SL g719 ( .A(n_552), .Y(n_719) );
AND2x4_ASAP7_75t_SL g552 ( .A(n_553), .B(n_565), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g596 ( .A(n_554), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
INVx1_ASAP7_75t_L g643 ( .A(n_554), .Y(n_643) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .C(n_559), .Y(n_556) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_565), .Y(n_585) );
AND2x4_ASAP7_75t_L g642 ( .A(n_565), .B(n_643), .Y(n_642) );
NOR2x1_ASAP7_75t_L g703 ( .A(n_565), .B(n_672), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g667 ( .A(n_567), .B(n_610), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_567), .A2(n_748), .B(n_749), .Y(n_747) );
INVx2_ASAP7_75t_L g625 ( .A(n_568), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_569), .A2(n_679), .B1(n_683), .B2(n_686), .Y(n_678) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_570), .Y(n_636) );
AND2x2_ASAP7_75t_L g646 ( .A(n_570), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g685 ( .A(n_570), .Y(n_685) );
NAND2x1_ASAP7_75t_SL g710 ( .A(n_570), .B(n_579), .Y(n_710) );
AND2x2_ASAP7_75t_L g606 ( .A(n_572), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2x1_ASAP7_75t_L g582 ( .A(n_574), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g579 ( .A(n_575), .Y(n_579) );
INVx2_ASAP7_75t_L g591 ( .A(n_575), .Y(n_591) );
AOI21xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_584), .B(n_588), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_579), .B(n_773), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_580), .A2(n_669), .B1(n_673), .B2(n_676), .Y(n_668) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
BUFx2_ASAP7_75t_L g773 ( .A(n_581), .Y(n_773) );
INVx1_ASAP7_75t_SL g780 ( .A(n_581), .Y(n_780) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_582), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OA21x2_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_592), .B(n_595), .Y(n_588) );
AND2x2_ASAP7_75t_L g592 ( .A(n_590), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g634 ( .A(n_590), .B(n_630), .Y(n_634) );
AND2x2_ASAP7_75t_L g749 ( .A(n_590), .B(n_647), .Y(n_749) );
AND2x2_ASAP7_75t_L g752 ( .A(n_590), .B(n_658), .Y(n_752) );
AND2x4_ASAP7_75t_L g760 ( .A(n_590), .B(n_761), .Y(n_760) );
OAI21xp33_ASAP7_75t_L g714 ( .A1(n_592), .A2(n_715), .B(n_717), .Y(n_714) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g742 ( .A(n_594), .Y(n_742) );
AND2x2_ASAP7_75t_L g758 ( .A(n_594), .B(n_759), .Y(n_758) );
INVx4_ASAP7_75t_L g672 ( .A(n_596), .Y(n_672) );
INVx1_ASAP7_75t_L g641 ( .A(n_597), .Y(n_641) );
AND2x2_ASAP7_75t_L g663 ( .A(n_597), .B(n_616), .Y(n_663) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_622), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B(n_608), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g609 ( .A(n_601), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_SL g762 ( .A(n_601), .B(n_614), .Y(n_762) );
AND2x2_ASAP7_75t_L g783 ( .A(n_601), .B(n_699), .Y(n_783) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g709 ( .A(n_606), .Y(n_709) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_611), .B(n_618), .Y(n_608) );
OR2x6_ASAP7_75t_L g661 ( .A(n_610), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_617), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
OR2x2_ASAP7_75t_L g684 ( .A(n_619), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g781 ( .A(n_619), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_620), .B(n_754), .Y(n_753) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_635), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B1(n_632), .B2(n_634), .Y(n_623) );
OR2x2_ASAP7_75t_L g695 ( .A(n_625), .B(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_627), .Y(n_652) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g701 ( .A(n_630), .Y(n_701) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_644), .B2(n_646), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
AND2x4_ASAP7_75t_SL g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g644 ( .A(n_642), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g705 ( .A(n_645), .B(n_699), .Y(n_705) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_650), .B(n_690), .Y(n_649) );
NOR2xp67_ASAP7_75t_L g650 ( .A(n_651), .B(n_664), .Y(n_650) );
AOI21xp33_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_659), .Y(n_651) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp33_ASAP7_75t_SL g729 ( .A1(n_661), .A2(n_730), .B1(n_732), .B2(n_735), .Y(n_729) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_662), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g712 ( .A(n_663), .B(n_713), .Y(n_712) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B(n_668), .C(n_678), .Y(n_664) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp33_ASAP7_75t_SL g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVxp33_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g681 ( .A(n_672), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_673), .A2(n_693), .B1(n_694), .B2(n_697), .C(n_700), .Y(n_692) );
AND2x4_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g733 ( .A(n_674), .Y(n_733) );
INVx2_ASAP7_75t_SL g731 ( .A(n_677), .Y(n_731) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2x1_ASAP7_75t_L g730 ( .A(n_681), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g727 ( .A(n_687), .Y(n_727) );
INVx1_ASAP7_75t_L g756 ( .A(n_688), .Y(n_756) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_706), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_704), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g745 ( .A(n_696), .Y(n_745) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g766 ( .A(n_699), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g771 ( .A(n_699), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVxp33_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g724 ( .A(n_703), .Y(n_724) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_711), .B(n_714), .Y(n_706) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g767 ( .A(n_713), .Y(n_767) );
AND2x2_ASAP7_75t_L g755 ( .A(n_716), .B(n_756), .Y(n_755) );
NOR2xp33_ASAP7_75t_R g717 ( .A(n_718), .B(n_719), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_736), .C(n_763), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_729), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_726), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
OR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_750), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_738), .B(n_747), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_739), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_746), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_751), .B(n_757), .Y(n_750) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_760), .B(n_762), .Y(n_757) );
INVx1_ASAP7_75t_L g776 ( .A(n_760), .Y(n_776) );
AOI211xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_766), .B(n_768), .C(n_777), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_772), .B1(n_774), .B2(n_776), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_782), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
INVxp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
CKINVDCx11_ASAP7_75t_R g790 ( .A(n_784), .Y(n_790) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_799), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
INVxp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_800), .A2(n_813), .B(n_818), .Y(n_812) );
NOR2xp33_ASAP7_75t_SL g800 ( .A(n_801), .B(n_806), .Y(n_800) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
BUFx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_804), .Y(n_803) );
BUFx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
BUFx2_ASAP7_75t_L g819 ( .A(n_805), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_808), .B(n_812), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
CKINVDCx11_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
CKINVDCx8_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_814), .Y(n_817) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
endmodule