module fake_aes_1103_n_698 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_698);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_698;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_599;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g78 ( .A(n_17), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_61), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_28), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_13), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_9), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_58), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
BUFx2_ASAP7_75t_SL g85 ( .A(n_53), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_75), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_38), .Y(n_87) );
INVx2_ASAP7_75t_SL g88 ( .A(n_14), .Y(n_88) );
INVxp67_ASAP7_75t_L g89 ( .A(n_6), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_60), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_36), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_18), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_12), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_62), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_71), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_20), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_17), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_57), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_41), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_18), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_32), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_67), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_76), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_33), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_7), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_45), .Y(n_109) );
INVxp33_ASAP7_75t_L g110 ( .A(n_56), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_49), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_27), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_5), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_74), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_29), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_19), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_11), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_30), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_66), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_46), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_48), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_12), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_24), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_86), .Y(n_126) );
NOR2xp33_ASAP7_75t_R g127 ( .A(n_105), .B(n_31), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_118), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
NAND2x1_ASAP7_75t_L g133 ( .A(n_82), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_119), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_80), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_100), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_87), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_87), .A2(n_125), .B(n_91), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_89), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_84), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_91), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_86), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_84), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_92), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_109), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_95), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_96), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_102), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_86), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_96), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_117), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_93), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_101), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_101), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_85), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_125), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_103), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_108), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_85), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_132), .B(n_93), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_132), .B(n_94), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_151), .B(n_103), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
INVxp67_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_131), .B(n_110), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_158), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_137), .B(n_94), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
AOI22x1_ASAP7_75t_L g180 ( .A1(n_129), .A2(n_111), .B1(n_123), .B2(n_122), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_146), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_162), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_129), .B(n_124), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_166), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_149), .Y(n_185) );
NAND2x1_ASAP7_75t_L g186 ( .A(n_130), .B(n_111), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_130), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g192 ( .A(n_128), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_134), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_134), .B(n_104), .Y(n_195) );
AND2x6_ASAP7_75t_L g196 ( .A(n_135), .B(n_106), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_141), .B(n_145), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_141), .B(n_121), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_145), .B(n_124), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_148), .B(n_97), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_153), .B(n_123), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_153), .B(n_97), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
INVx4_ASAP7_75t_SL g206 ( .A(n_160), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
NAND3xp33_ASAP7_75t_L g208 ( .A(n_157), .B(n_99), .C(n_113), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_161), .B(n_122), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_161), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_164), .B(n_160), .Y(n_211) );
AND2x6_ASAP7_75t_L g212 ( .A(n_164), .B(n_120), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_142), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_138), .B(n_120), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_133), .B(n_99), .C(n_113), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
INVxp33_ASAP7_75t_L g217 ( .A(n_133), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_163), .Y(n_219) );
INVx4_ASAP7_75t_L g220 ( .A(n_163), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_140), .B(n_150), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_163), .B(n_116), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g224 ( .A(n_165), .B(n_108), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_163), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_146), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_146), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_144), .A2(n_81), .B1(n_107), .B2(n_98), .Y(n_228) );
NAND3x1_ASAP7_75t_L g229 ( .A(n_165), .B(n_116), .C(n_112), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_211), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_178), .B(n_155), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_211), .Y(n_232) );
BUFx4f_ASAP7_75t_SL g233 ( .A(n_177), .Y(n_233) );
CKINVDCx11_ASAP7_75t_R g234 ( .A(n_192), .Y(n_234) );
NOR3xp33_ASAP7_75t_SL g235 ( .A(n_215), .B(n_214), .C(n_176), .Y(n_235) );
BUFx2_ASAP7_75t_SL g236 ( .A(n_171), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_213), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_187), .B(n_165), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_176), .B(n_165), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_173), .B(n_127), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_175), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_223), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_183), .B(n_106), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_207), .Y(n_245) );
NOR2x1_ASAP7_75t_L g246 ( .A(n_208), .B(n_159), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_167), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_223), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_173), .B(n_78), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_174), .B(n_90), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_174), .B(n_115), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_198), .B(n_114), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_224), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_196), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_178), .B(n_147), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_196), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_196), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_194), .A2(n_112), .B(n_163), .C(n_152), .Y(n_259) );
AND2x6_ASAP7_75t_L g260 ( .A(n_218), .B(n_156), .Y(n_260) );
BUFx12f_ASAP7_75t_L g261 ( .A(n_167), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_183), .B(n_156), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_200), .B(n_1), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_179), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_200), .B(n_156), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_214), .B(n_37), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_169), .B(n_152), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_169), .B(n_152), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_222), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_195), .B(n_2), .C(n_3), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_168), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_202), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_196), .Y(n_273) );
INVxp33_ASAP7_75t_L g274 ( .A(n_228), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_202), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_204), .B(n_139), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_204), .B(n_2), .Y(n_278) );
OR2x6_ASAP7_75t_L g279 ( .A(n_229), .B(n_139), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_184), .B(n_35), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_171), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_197), .B(n_139), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_182), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_185), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_195), .B(n_3), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_199), .B(n_4), .C(n_5), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_201), .B(n_126), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_205), .B(n_126), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_171), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_212), .Y(n_290) );
NOR3xp33_ASAP7_75t_SL g291 ( .A(n_199), .B(n_4), .C(n_6), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g292 ( .A(n_209), .B(n_8), .Y(n_292) );
OR2x6_ASAP7_75t_L g293 ( .A(n_186), .B(n_126), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_171), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_209), .B(n_8), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_273), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_261), .Y(n_297) );
OR2x6_ASAP7_75t_SL g298 ( .A(n_242), .B(n_217), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_289), .B(n_189), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_237), .Y(n_300) );
NOR2x1_ASAP7_75t_SL g301 ( .A(n_236), .B(n_210), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_263), .A2(n_295), .B1(n_285), .B2(n_244), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_283), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_273), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_244), .B(n_217), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_264), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_274), .B(n_203), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_264), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_273), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_284), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_245), .Y(n_315) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_242), .A2(n_180), .B1(n_190), .B2(n_203), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_263), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_239), .B(n_171), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_243), .A2(n_219), .B(n_225), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_230), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_269), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_263), .A2(n_188), .B1(n_220), .B2(n_216), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_233), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_248), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_247), .Y(n_327) );
AOI21xp33_ASAP7_75t_L g328 ( .A1(n_266), .A2(n_188), .B(n_220), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_285), .A2(n_212), .B1(n_216), .B2(n_221), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_234), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_230), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_231), .B(n_212), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_287), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_247), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_256), .B(n_9), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_256), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_289), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_239), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_250), .Y(n_339) );
INVx4_ASAP7_75t_L g340 ( .A(n_289), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_254), .B(n_212), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_288), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_232), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_243), .A2(n_193), .B(n_191), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_249), .A2(n_191), .B(n_226), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_343), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_336), .A2(n_246), .B1(n_285), .B2(n_295), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_343), .B(n_295), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_336), .A2(n_272), .B1(n_278), .B2(n_244), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_303), .A2(n_292), .B1(n_278), .B2(n_275), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_303), .A2(n_240), .B1(n_253), .B2(n_279), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_343), .B(n_232), .Y(n_352) );
AOI22xp33_ASAP7_75t_SL g353 ( .A1(n_318), .A2(n_236), .B1(n_254), .B2(n_279), .Y(n_353) );
OR2x6_ASAP7_75t_SL g354 ( .A(n_335), .B(n_298), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_300), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_300), .Y(n_356) );
AOI21x1_ASAP7_75t_L g357 ( .A1(n_345), .A2(n_262), .B(n_277), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_309), .A2(n_279), .B1(n_249), .B2(n_268), .Y(n_358) );
CKINVDCx9p33_ASAP7_75t_R g359 ( .A(n_297), .Y(n_359) );
INVxp67_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_313), .Y(n_361) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_318), .B(n_294), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_299), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_304), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_300), .A2(n_241), .B(n_294), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_322), .A2(n_279), .B1(n_267), .B2(n_251), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_304), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_322), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_331), .B(n_235), .Y(n_369) );
INVx4_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_316), .A2(n_259), .B(n_291), .Y(n_371) );
INVx4_ASAP7_75t_SL g372 ( .A(n_313), .Y(n_372) );
CKINVDCx11_ASAP7_75t_R g373 ( .A(n_330), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_331), .Y(n_374) );
NAND2xp33_ASAP7_75t_R g375 ( .A(n_297), .B(n_270), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_310), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g378 ( .A(n_364), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_368), .B(n_335), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_367), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_349), .B(n_339), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_368), .A2(n_324), .B1(n_310), .B2(n_323), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_357), .A2(n_344), .B(n_308), .Y(n_383) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_360), .A2(n_234), .B(n_286), .C(n_325), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_374), .A2(n_324), .B1(n_310), .B2(n_307), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_350), .A2(n_326), .B1(n_306), .B2(n_302), .C(n_314), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_357), .A2(n_308), .B(n_307), .Y(n_388) );
BUFx12f_ASAP7_75t_L g389 ( .A(n_373), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_375), .B(n_302), .C(n_238), .D(n_325), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_376), .B(n_311), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_363), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g393 ( .A1(n_347), .A2(n_332), .B1(n_329), .B2(n_314), .C(n_311), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_352), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g395 ( .A1(n_369), .A2(n_298), .B1(n_317), .B2(n_333), .C1(n_342), .C2(n_338), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_351), .A2(n_334), .B1(n_308), .B2(n_342), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_376), .B(n_317), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_374), .B(n_317), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_363), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_364), .B(n_338), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_351), .A2(n_334), .B1(n_333), .B2(n_342), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_350), .A2(n_341), .B1(n_319), .B2(n_333), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_395), .A2(n_371), .B1(n_362), .B2(n_358), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_397), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_397), .B(n_355), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_399), .Y(n_407) );
BUFx2_ASAP7_75t_L g408 ( .A(n_399), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_398), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_381), .A2(n_366), .B1(n_352), .B2(n_348), .C(n_252), .Y(n_410) );
OR2x6_ASAP7_75t_L g411 ( .A(n_399), .B(n_363), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_380), .Y(n_412) );
OAI211xp5_ASAP7_75t_SL g413 ( .A1(n_401), .A2(n_354), .B(n_359), .C(n_353), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_391), .B(n_355), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
NOR4xp25_ASAP7_75t_SL g416 ( .A(n_384), .B(n_371), .C(n_372), .D(n_328), .Y(n_416) );
OAI21xp5_ASAP7_75t_SL g417 ( .A1(n_395), .A2(n_341), .B(n_319), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_387), .B(n_265), .C(n_348), .D(n_280), .Y(n_418) );
OAI33xp33_ASAP7_75t_L g419 ( .A1(n_390), .A2(n_356), .A3(n_355), .B1(n_371), .B2(n_14), .B3(n_15), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_371), .B1(n_362), .B2(n_356), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_388), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_394), .A2(n_362), .B1(n_356), .B2(n_370), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_390), .A2(n_320), .B1(n_341), .B2(n_319), .C(n_365), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_370), .B1(n_341), .B2(n_319), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_379), .B(n_370), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_391), .B(n_370), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_382), .A2(n_327), .B1(n_299), .B2(n_340), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_398), .Y(n_429) );
OA21x2_ASAP7_75t_L g430 ( .A1(n_388), .A2(n_328), .B(n_271), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_393), .A2(n_327), .B1(n_271), .B2(n_255), .C(n_258), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_389), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_385), .A2(n_299), .B(n_260), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_403), .A2(n_327), .B1(n_340), .B2(n_337), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_386), .B(n_372), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_379), .B(n_293), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_386), .B(n_392), .Y(n_438) );
NAND4xp25_ASAP7_75t_SL g439 ( .A(n_382), .B(n_10), .C(n_11), .D(n_13), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_414), .B(n_392), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_414), .B(n_385), .Y(n_441) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_423), .B(n_340), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_436), .B(n_383), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_421), .Y(n_444) );
OAI33xp33_ASAP7_75t_L g445 ( .A1(n_412), .A2(n_396), .A3(n_400), .B1(n_16), .B2(n_19), .B3(n_20), .Y(n_445) );
NAND3xp33_ASAP7_75t_SL g446 ( .A(n_416), .B(n_389), .C(n_290), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_415), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_421), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_419), .A2(n_337), .B1(n_172), .B2(n_181), .C(n_226), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_406), .B(n_383), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_406), .B(n_372), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_432), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_405), .B(n_372), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_405), .B(n_372), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_417), .A2(n_337), .B1(n_294), .B2(n_257), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_415), .B(n_361), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_411), .Y(n_458) );
AOI322xp5_ASAP7_75t_L g459 ( .A1(n_433), .A2(n_10), .A3(n_15), .B1(n_16), .B2(n_21), .C1(n_22), .C2(n_23), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_409), .B(n_21), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_439), .A2(n_337), .B1(n_170), .B2(n_227), .C(n_181), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_438), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_427), .B(n_438), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_408), .Y(n_465) );
AND2x4_ASAP7_75t_SL g466 ( .A(n_411), .B(n_361), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_436), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_430), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_430), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_423), .B(n_361), .Y(n_470) );
OAI33xp33_ASAP7_75t_L g471 ( .A1(n_413), .A2(n_22), .A3(n_23), .B1(n_25), .B2(n_26), .B3(n_34), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_420), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_426), .B(n_361), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_430), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_427), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_407), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_404), .A2(n_293), .B1(n_321), .B2(n_296), .C(n_290), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_407), .B(n_361), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_411), .B(n_361), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_411), .B(n_301), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_411), .B(n_39), .Y(n_485) );
INVx2_ASAP7_75t_SL g486 ( .A(n_425), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_425), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_428), .Y(n_488) );
INVx5_ASAP7_75t_L g489 ( .A(n_434), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_416), .B(n_42), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_410), .B(n_301), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_449), .Y(n_492) );
NAND2xp33_ASAP7_75t_SL g493 ( .A(n_485), .B(n_433), .Y(n_493) );
NAND2xp33_ASAP7_75t_R g494 ( .A(n_460), .B(n_43), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_447), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_480), .B(n_437), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_461), .B(n_422), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g498 ( .A(n_459), .B(n_418), .C(n_424), .D(n_428), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_464), .B(n_418), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_451), .B(n_435), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_451), .B(n_44), .Y(n_502) );
NOR2xp33_ASAP7_75t_R g503 ( .A(n_442), .B(n_296), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_464), .B(n_47), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_478), .B(n_51), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_441), .B(n_52), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_461), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_459), .B(n_431), .C(n_257), .D(n_276), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_480), .B(n_260), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_465), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_474), .B(n_54), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_449), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_441), .B(n_55), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_460), .A2(n_276), .A3(n_258), .B(n_255), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_478), .B(n_59), .Y(n_518) );
NOR3x1_ASAP7_75t_L g519 ( .A(n_446), .B(n_63), .C(n_64), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_440), .B(n_65), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_467), .B(n_68), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_467), .B(n_69), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_449), .B(n_72), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_440), .B(n_73), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_453), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_474), .B(n_77), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_453), .B(n_206), .Y(n_527) );
NAND2xp33_ASAP7_75t_L g528 ( .A(n_485), .B(n_313), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_453), .Y(n_529) );
OAI322xp33_ASAP7_75t_L g530 ( .A1(n_472), .A2(n_170), .A3(n_172), .B1(n_181), .B2(n_227), .C1(n_226), .C2(n_191), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_479), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_460), .B(n_260), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_488), .B(n_293), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_458), .B(n_312), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_443), .B(n_206), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_473), .B(n_293), .Y(n_536) );
OAI21xp33_ASAP7_75t_SL g537 ( .A1(n_442), .A2(n_321), .B(n_296), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_479), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_457), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_458), .B(n_312), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_487), .B(n_260), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_443), .B(n_206), .Y(n_542) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_450), .B(n_170), .C(n_172), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_487), .B(n_260), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_443), .B(n_170), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_443), .B(n_172), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_444), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_486), .B(n_260), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_457), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_452), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_473), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_507), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_498), .A2(n_445), .B1(n_515), .B2(n_512), .C(n_500), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_539), .B(n_549), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_543), .A2(n_450), .B(n_442), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_495), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_538), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_499), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_497), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_497), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_551), .B(n_486), .Y(n_561) );
AOI32xp33_ASAP7_75t_L g562 ( .A1(n_493), .A2(n_462), .A3(n_484), .B1(n_458), .B2(n_486), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_510), .B(n_458), .Y(n_563) );
OAI32xp33_ASAP7_75t_L g564 ( .A1(n_494), .A2(n_493), .A3(n_537), .B1(n_538), .B2(n_526), .Y(n_564) );
AOI31xp33_ASAP7_75t_L g565 ( .A1(n_504), .A2(n_471), .A3(n_445), .B(n_462), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_531), .Y(n_566) );
OAI21xp33_ASAP7_75t_SL g567 ( .A1(n_511), .A2(n_526), .B(n_504), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_516), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_529), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_520), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_508), .A2(n_475), .B1(n_472), .B2(n_488), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_519), .B(n_481), .C(n_446), .D(n_475), .Y(n_572) );
OA22x2_ASAP7_75t_L g573 ( .A1(n_550), .A2(n_484), .B1(n_466), .B2(n_452), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_524), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_502), .Y(n_575) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_511), .A2(n_491), .B(n_481), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_492), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_492), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_513), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_513), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_525), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_505), .A2(n_491), .B1(n_489), .B2(n_484), .Y(n_582) );
AOI21xp33_ASAP7_75t_SL g583 ( .A1(n_502), .A2(n_484), .B(n_456), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g584 ( .A1(n_503), .A2(n_490), .B(n_470), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_496), .B(n_476), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_503), .A2(n_489), .B1(n_466), .B2(n_483), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_501), .B(n_454), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_501), .A2(n_471), .B1(n_476), .B2(n_470), .C(n_477), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_547), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_506), .B(n_454), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_545), .B(n_483), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g593 ( .A1(n_517), .A2(n_456), .B1(n_489), .B2(n_490), .C(n_477), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_506), .A2(n_468), .B1(n_469), .B2(n_477), .C(n_455), .Y(n_594) );
NAND2x1_ASAP7_75t_L g595 ( .A(n_523), .B(n_546), .Y(n_595) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_528), .B(n_455), .Y(n_596) );
AOI32xp33_ASAP7_75t_L g597 ( .A1(n_528), .A2(n_483), .A3(n_466), .B1(n_482), .B2(n_468), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_523), .Y(n_598) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_530), .B(n_482), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_547), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_545), .B(n_489), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_546), .B(n_489), .Y(n_602) );
NAND2x1_ASAP7_75t_SL g603 ( .A(n_518), .B(n_469), .Y(n_603) );
AOI21xp33_ASAP7_75t_L g604 ( .A1(n_521), .A2(n_469), .B(n_468), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_592), .B(n_489), .Y(n_605) );
XNOR2xp5_ASAP7_75t_L g606 ( .A(n_557), .B(n_514), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_577), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_567), .A2(n_514), .B1(n_532), .B2(n_518), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_570), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_553), .B(n_533), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_559), .B(n_533), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_588), .B(n_489), .Y(n_612) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_572), .B(n_522), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_564), .A2(n_534), .B(n_540), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_556), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_560), .B(n_548), .Y(n_617) );
NOR2x1_ASAP7_75t_L g618 ( .A(n_599), .B(n_522), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_571), .A2(n_509), .B1(n_544), .B2(n_541), .C(n_536), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_568), .B(n_540), .Y(n_620) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_566), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_554), .B(n_540), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_586), .B(n_534), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_552), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_573), .A2(n_534), .B1(n_535), .B2(n_542), .Y(n_625) );
INVx3_ASAP7_75t_SL g626 ( .A(n_573), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_558), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_569), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_586), .B(n_448), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_574), .A2(n_542), .B1(n_535), .B2(n_527), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_561), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_578), .Y(n_632) );
CKINVDCx14_ASAP7_75t_R g633 ( .A(n_598), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_579), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_589), .B(n_448), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_565), .A2(n_448), .B(n_444), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_580), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_562), .A2(n_444), .B1(n_527), .B2(n_296), .C(n_321), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_581), .Y(n_639) );
BUFx3_ASAP7_75t_L g640 ( .A(n_563), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_585), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_615), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_626), .A2(n_583), .B(n_584), .C(n_576), .Y(n_643) );
XNOR2x1_ASAP7_75t_L g644 ( .A(n_613), .B(n_596), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_610), .B(n_593), .C(n_576), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_616), .B(n_563), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_618), .A2(n_587), .B(n_597), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_614), .A2(n_555), .B(n_595), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_636), .B(n_594), .C(n_604), .Y(n_649) );
NAND4xp75_ASAP7_75t_L g650 ( .A(n_608), .B(n_604), .C(n_602), .D(n_601), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_615), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_633), .B(n_575), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_628), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_626), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_606), .A2(n_582), .B1(n_591), .B2(n_600), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_621), .A2(n_582), .B(n_590), .C(n_603), .Y(n_656) );
INVx3_ASAP7_75t_L g657 ( .A(n_640), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_628), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_631), .B(n_181), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_607), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_609), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_640), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g663 ( .A1(n_606), .A2(n_321), .B1(n_312), .B2(n_305), .C(n_226), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_633), .B(n_227), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_648), .A2(n_638), .B(n_625), .C(n_605), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_645), .B(n_635), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_642), .Y(n_667) );
AOI21xp33_ASAP7_75t_SL g668 ( .A1(n_644), .A2(n_620), .B(n_630), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g669 ( .A1(n_655), .A2(n_622), .A3(n_623), .B1(n_624), .B2(n_627), .C1(n_611), .C2(n_617), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_656), .A2(n_619), .B1(n_639), .B2(n_634), .C(n_641), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_643), .B(n_641), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_651), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_647), .A2(n_605), .B1(n_629), .B2(n_612), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_661), .B(n_612), .Y(n_674) );
INVx2_ASAP7_75t_SL g675 ( .A(n_662), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_654), .B(n_652), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_644), .A2(n_637), .B(n_632), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_654), .B(n_637), .Y(n_678) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_654), .A2(n_632), .B(n_607), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_657), .A2(n_305), .B(n_313), .C(n_258), .Y(n_680) );
AOI32xp33_ASAP7_75t_L g681 ( .A1(n_652), .A2(n_305), .A3(n_255), .B1(n_281), .B2(n_313), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_649), .B(n_227), .Y(n_682) );
AOI322xp5_ASAP7_75t_L g683 ( .A1(n_662), .A2(n_281), .A3(n_313), .B1(n_657), .B2(n_646), .C1(n_653), .C2(n_658), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_664), .A2(n_657), .B(n_663), .C(n_659), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_660), .Y(n_685) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_650), .B(n_664), .Y(n_686) );
OR3x2_ASAP7_75t_L g687 ( .A(n_686), .B(n_673), .C(n_665), .Y(n_687) );
AOI31xp33_ASAP7_75t_L g688 ( .A1(n_670), .A2(n_666), .A3(n_671), .B(n_676), .Y(n_688) );
NAND3xp33_ASAP7_75t_SL g689 ( .A(n_668), .B(n_683), .C(n_677), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_669), .A2(n_675), .B1(n_679), .B2(n_682), .C(n_674), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_687), .Y(n_691) );
AND2x2_ASAP7_75t_SL g692 ( .A(n_690), .B(n_678), .Y(n_692) );
AND3x2_ASAP7_75t_L g693 ( .A(n_688), .B(n_678), .C(n_667), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_691), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_693), .Y(n_695) );
INVx4_ASAP7_75t_L g696 ( .A(n_694), .Y(n_696) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_695), .A3(n_692), .B1(n_689), .B2(n_693), .C1(n_672), .C2(n_685), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_697), .A2(n_684), .B1(n_681), .B2(n_680), .C(n_660), .Y(n_698) );
endmodule