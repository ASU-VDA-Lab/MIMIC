module real_jpeg_6913_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

BUFx5_ASAP7_75t_L g313 ( 
.A(n_0),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_0),
.Y(n_321)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_1),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_1),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g442 ( 
.A(n_1),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_1),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_2),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_2),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_2),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_2),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_2),
.B(n_285),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_2),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_2),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_2),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_3),
.B(n_64),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_3),
.B(n_52),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_3),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_3),
.B(n_259),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_4),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g427 ( 
.A(n_4),
.Y(n_427)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_5),
.Y(n_511)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_6),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_6),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_7),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_7),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_7),
.B(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_7),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_7),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_7),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_7),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_7),
.B(n_467),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_8),
.B(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_8),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_8),
.B(n_235),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_8),
.B(n_429),
.Y(n_428)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_12),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_12),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_12),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_12),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_12),
.B(n_395),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_13),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_14),
.B(n_87),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_14),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_14),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_14),
.B(n_280),
.Y(n_305)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_14),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_14),
.B(n_129),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_15),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_15),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g374 ( 
.A(n_15),
.B(n_301),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_15),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_16),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_16),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_16),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_16),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_16),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_17),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_17),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_17),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_17),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_17),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_17),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_17),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_17),
.B(n_415),
.Y(n_414)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_19),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_19),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_19),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_19),
.B(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_19),
.B(n_423),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_510),
.B(n_512),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_173),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_172),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_148),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_148),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_112),
.C(n_124),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_25),
.B(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_80),
.C(n_94),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_26),
.B(n_498),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_43),
.C(n_59),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_27),
.B(n_43),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_28),
.B(n_37),
.C(n_42),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_29),
.B(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_31),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_42),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_35),
.Y(n_260)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_36),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_40),
.Y(n_246)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_40),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_40),
.Y(n_425)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_41),
.Y(n_217)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_41),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.C(n_54),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_44),
.B(n_54),
.Y(n_457)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_48),
.Y(n_135)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_48),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_49),
.B(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_53),
.Y(n_395)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_59),
.B(n_487),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_67),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_60),
.B(n_68),
.C(n_79),
.Y(n_122)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_65),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_66),
.Y(n_198)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_66),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_79),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_69),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_115),
.C(n_119),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_72),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_72),
.Y(n_339)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_97),
.C(n_101),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_73),
.A2(n_79),
.B1(n_97),
.B2(n_98),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_78),
.Y(n_297)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_78),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_80),
.A2(n_94),
.B1(n_95),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_80),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_86),
.C(n_89),
.Y(n_140)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.C(n_110),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_96),
.B(n_485),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_97),
.A2(n_98),
.B1(n_436),
.B2(n_439),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_97),
.B(n_436),
.C(n_440),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_100),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_101),
.B(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_104),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_485)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_110),
.A2(n_111),
.B1(n_466),
.B2(n_468),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_111),
.B(n_468),
.C(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_112),
.B(n_124),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_122),
.C(n_123),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_113),
.B(n_501),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_116),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_132),
.C(n_136),
.Y(n_169)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_122),
.B(n_123),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_139),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_137),
.B2(n_138),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_138),
.C(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_131),
.B2(n_136),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_133),
.B1(n_161),
.B2(n_166),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_144),
.C(n_147),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_142),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_167),
.B2(n_168),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_161),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_165),
.Y(n_397)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

AO21x1_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_490),
.B(n_507),
.Y(n_173)
);

OAI21x1_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_473),
.B(n_489),
.Y(n_174)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_446),
.B(n_472),
.Y(n_175)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_401),
.B(n_445),
.Y(n_176)
);

AOI21x1_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_364),
.B(n_400),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_290),
.B(n_363),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_273),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_180),
.B(n_273),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_224),
.B2(n_272),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_181),
.B(n_225),
.C(n_256),
.Y(n_399)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_201),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_183),
.B(n_202),
.C(n_223),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_195),
.C(n_199),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_184),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_185),
.A2(n_186),
.B1(n_191),
.B2(n_192),
.Y(n_278)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_194),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_195),
.B(n_199),
.Y(n_289)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_210),
.B1(n_222),
.B2(n_223),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_205),
.B(n_209),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.Y(n_209)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_209),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_209),
.B(n_369),
.C(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_210),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.CI(n_218),
.CON(n_210),
.SN(n_210)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_211),
.B(n_214),
.C(n_218),
.Y(n_398)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_256),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_238),
.C(n_249),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_231),
.C(n_234),
.Y(n_271)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_239),
.B1(n_249),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.C(n_247),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_240),
.A2(n_241),
.B1(n_247),
.B2(n_248),
.Y(n_356)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_242),
.B(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_246),
.Y(n_333)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_253),
.Y(n_270)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_269),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_257),
.B(n_270),
.C(n_271),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g379 ( 
.A(n_258),
.B(n_265),
.C(n_267),
.Y(n_379)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.C(n_288),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_274),
.B(n_361),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_277),
.B(n_288),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_279),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_281),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_282),
.B(n_284),
.Y(n_327)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_286),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_358),
.B(n_362),
.Y(n_290)
);

OA21x2_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_343),
.B(n_357),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_324),
.B(n_342),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_314),
.B(n_323),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_302),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_302),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_298),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_309),
.B2(n_310),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_306),
.C(n_309),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_312),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_318),
.B(n_322),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_341),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_341),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_328),
.C(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_336),
.C(n_340),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_337),
.B2(n_340),
.Y(n_334)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_346),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_353),
.C(n_354),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_360),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_399),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_399),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_381),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_368),
.C(n_381),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_370),
.B1(n_378),
.B2(n_380),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_374),
.C(n_375),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_375),
.B2(n_376),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_378),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_384),
.C(n_392),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_392),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_387),
.C(n_389),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

INVx6_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_398),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_396),
.C(n_398),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_403),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_404),
.B(n_420),
.C(n_443),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_406),
.A2(n_420),
.B1(n_443),
.B2(n_444),
.Y(n_405)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_406),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_409),
.B2(n_419),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_410),
.C(n_411),
.Y(n_448)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_409),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_418),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_413),
.B(n_414),
.C(n_418),
.Y(n_463)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_420),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_431),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_432),
.C(n_433),
.Y(n_461)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_421),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_426),
.CI(n_428),
.CON(n_421),
.SN(n_421)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_426),
.C(n_428),
.Y(n_469)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_440),
.B2(n_441),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_436),
.Y(n_439)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_471),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_471),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_450),
.C(n_459),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_459),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_452),
.B1(n_454),
.B2(n_458),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_455),
.C(n_456),
.Y(n_479)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_454),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_461),
.B1(n_462),
.B2(n_470),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_463),
.C(n_464),
.Y(n_475)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_469),
.Y(n_464)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_466),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_469),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_488),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_488),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_475),
.B(n_477),
.C(n_486),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_486),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_481),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_482),
.C(n_484),
.Y(n_502)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.Y(n_481)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_503),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_496),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_500),
.C(n_502),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_500),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_502),
.B(n_505),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_506),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_506),
.Y(n_508)
);

INVx8_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx13_ASAP7_75t_L g513 ( 
.A(n_511),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_514),
.Y(n_512)
);


endmodule