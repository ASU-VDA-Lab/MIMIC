module fake_jpeg_963_n_221 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_221);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_0),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_54),
.B1(n_60),
.B2(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_77),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_63),
.B1(n_57),
.B2(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_80),
.B1(n_57),
.B2(n_67),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_54),
.B1(n_73),
.B2(n_52),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_54),
.B1(n_73),
.B2(n_52),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_101),
.B1(n_72),
.B2(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_98),
.B(n_102),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_66),
.B1(n_62),
.B2(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_107),
.Y(n_126)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_69),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_110),
.Y(n_131)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_72),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_65),
.C(n_53),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_97),
.C(n_96),
.Y(n_121)
);

CKINVDCx12_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_7),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_95),
.B(n_94),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_134),
.B(n_3),
.Y(n_143)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_86),
.B(n_91),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_65),
.B(n_53),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_34),
.C(n_40),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_39),
.B1(n_38),
.B2(n_36),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_51),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_50),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_128),
.Y(n_146)
);

BUFx12f_ASAP7_75t_SL g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_4),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_65),
.B(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_138),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_143),
.B(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_53),
.B1(n_49),
.B2(n_48),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_145),
.B1(n_32),
.B2(n_29),
.Y(n_168)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_147),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_144),
.C(n_150),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_41),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_154),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_4),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_152),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_33),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_115),
.C(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_13),
.C(n_14),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_12),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_9),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

OAI22x1_ASAP7_75t_SL g159 ( 
.A1(n_151),
.A2(n_143),
.B1(n_140),
.B2(n_137),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_162),
.B1(n_168),
.B2(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

AO21x1_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_127),
.B(n_118),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_165),
.B(n_15),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_130),
.B1(n_129),
.B2(n_133),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_130),
.B(n_129),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_172),
.B(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_27),
.B(n_25),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_16),
.C(n_17),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_176),
.B(n_23),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_14),
.B(n_15),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_179),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_150),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_185),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_191),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_16),
.Y(n_188)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_189),
.B(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_167),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_159),
.B1(n_177),
.B2(n_173),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_195),
.B1(n_194),
.B2(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_161),
.B(n_165),
.C(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_171),
.C(n_170),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_200),
.C(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_181),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_171),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_205),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_206),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g213 ( 
.A(n_210),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_202),
.C(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_212),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_213),
.B(n_211),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_198),
.A3(n_203),
.B1(n_197),
.B2(n_212),
.C1(n_195),
.C2(n_182),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_17),
.A3(n_18),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_22),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_219),
.B(n_18),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_19),
.Y(n_221)
);


endmodule