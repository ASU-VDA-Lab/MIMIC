module real_jpeg_17775_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_535),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_0),
.B(n_536),
.Y(n_535)
);

AND2x2_ASAP7_75t_SL g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_1),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_1),
.B(n_58),
.Y(n_176)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_2),
.Y(n_315)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_2),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_3),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g450 ( 
.A(n_3),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_4),
.B(n_58),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_4),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_4),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_4),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_4),
.B(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_4),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_4),
.B(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_4),
.B(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_5),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_6),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_6),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_6),
.B(n_93),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_6),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_6),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_7),
.Y(n_174)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_7),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_7),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g459 ( 
.A(n_7),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_8),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_8),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_8),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_8),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_8),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_8),
.A2(n_9),
.B1(n_289),
.B2(n_294),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_9),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_9),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g308 ( 
.A(n_9),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_9),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_9),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_9),
.B(n_500),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_10),
.Y(n_136)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_10),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_10),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_10),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_11),
.B(n_110),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_11),
.B(n_214),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_11),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g313 ( 
.A(n_11),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_11),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_11),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_11),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_11),
.B(n_459),
.Y(n_458)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_12),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_12),
.Y(n_322)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_13),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_13),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_13),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_13),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_13),
.B(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_15),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_15),
.B(n_40),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_15),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_15),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_15),
.B(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_15),
.B(n_426),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_15),
.B(n_510),
.Y(n_509)
);

BUFx4f_ASAP7_75t_L g142 ( 
.A(n_16),
.Y(n_142)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_16),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g464 ( 
.A(n_16),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_16),
.Y(n_498)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_17),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_17),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_23),
.B(n_71),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_23),
.Y(n_537)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_38),
.CI(n_51),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.C(n_33),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_25),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_25),
.A2(n_26),
.B1(n_60),
.B2(n_61),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_25),
.B(n_164),
.C(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_25),
.A2(n_26),
.B1(n_235),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_60),
.C(n_65),
.Y(n_59)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_29),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_30),
.B(n_128),
.C(n_133),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_30),
.B(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_32),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_34),
.B1(n_44),
.B2(n_48),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_33),
.B(n_249),
.C(n_258),
.Y(n_248)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_35),
.A2(n_258),
.B1(n_259),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_35),
.Y(n_380)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_36),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_78),
.C(n_83),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_39),
.A2(n_49),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_44),
.B(n_139),
.C(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_44),
.B(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.C(n_59),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_60),
.A2(n_61),
.B1(n_103),
.B2(n_104),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_60),
.A2(n_61),
.B1(n_159),
.B2(n_160),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_103),
.C(n_108),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_61),
.B(n_160),
.C(n_296),
.Y(n_353)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2x1_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.C(n_96),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g119 ( 
.A(n_76),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_87),
.C(n_91),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_81),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_83),
.B(n_208),
.C(n_212),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_83),
.B(n_212),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_91),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_91),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_91),
.B(n_207),
.C(n_213),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_91),
.A2(n_92),
.B1(n_213),
.B2(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_92),
.B(n_176),
.Y(n_217)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_94),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_95),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.C(n_111),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_98),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_101),
.B(n_170),
.C(n_175),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_103),
.A2(n_104),
.B1(n_138),
.B2(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_103),
.A2(n_104),
.B1(n_308),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_138),
.C(n_143),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_104),
.B(n_308),
.C(n_310),
.Y(n_307)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_106),
.Y(n_351)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_107),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21x1_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_177),
.B(n_533),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_117),
.B(n_120),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_145),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.C(n_137),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_125),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_127),
.B(n_137),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_133),
.A2(n_164),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_136),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_139),
.B1(n_172),
.B2(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_139),
.B(n_255),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_139),
.B(n_360),
.Y(n_423)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_144),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_165),
.C(n_169),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_162),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_148),
.B(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_150),
.B(n_162),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.C(n_159),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_154),
.Y(n_311)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_154),
.Y(n_482)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AO22x1_ASAP7_75t_SL g216 ( 
.A1(n_170),
.A2(n_171),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_195),
.C(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_172),
.A2(n_173),
.B1(n_199),
.B2(n_200),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_172),
.B(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_173),
.B(n_430),
.Y(n_466)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_174),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_174),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_261),
.B(n_530),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_219),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_181),
.A2(n_531),
.B(n_532),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_182),
.B(n_184),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_206),
.C(n_216),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_191),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_204),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_192),
.B(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_194),
.B(n_204),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_196),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_196),
.B(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_199),
.A2(n_200),
.B1(n_303),
.B2(n_304),
.Y(n_327)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_200),
.B(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_201),
.Y(n_319)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_216),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

OR2x6_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_220),
.B(n_222),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.C(n_229),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_223),
.B(n_226),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_229),
.B(n_411),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_242),
.C(n_247),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_230),
.A2(n_231),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.C(n_239),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_232),
.B(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_234),
.A2(n_239),
.B1(n_240),
.B2(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_234),
.Y(n_388)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_235),
.Y(n_343)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_400)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_249),
.A2(n_250),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_251),
.A2(n_255),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_251),
.Y(n_359)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_252),
.Y(n_432)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_254),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_255),
.Y(n_360)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_257),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_260),
.Y(n_428)
);

NAND2x1_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_413),
.Y(n_261)
);

A2O1A1O1Ixp25_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_390),
.B(n_406),
.C(n_407),
.D(n_412),
.Y(n_262)
);

OAI21x1_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_366),
.B(n_389),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_337),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g529 ( 
.A(n_265),
.B(n_337),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_298),
.C(n_323),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_266),
.B(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_278),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_267),
.B(n_279),
.C(n_295),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.C(n_273),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_268),
.B(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_269),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_421)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_295),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_285),
.B(n_288),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_288),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_288),
.Y(n_363)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_298),
.A2(n_299),
.B1(n_323),
.B2(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_312),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_306),
.B2(n_307),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_301),
.B(n_307),
.C(n_312),
.Y(n_354)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_308),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_310),
.B(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_313),
.B(n_317),
.C(n_320),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_323),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.C(n_328),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_324),
.B(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_327),
.B(n_328),
.Y(n_419)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.C(n_335),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_329),
.B(n_335),
.Y(n_471)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_332),
.B(n_471),
.Y(n_470)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_355),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_356),
.C(n_365),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_354),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_344),
.Y(n_339)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_353),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_349),
.B1(n_350),
.B2(n_352),
.Y(n_345)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_346),
.Y(n_352)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_350),
.B(n_353),
.C(n_382),
.Y(n_381)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_352),
.Y(n_382)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_370),
.C(n_371),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_365),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_361),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_363),
.C(n_364),
.Y(n_375)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_362),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g528 ( 
.A(n_366),
.B(n_529),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_368),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_368),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_369),
.B(n_392),
.C(n_393),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_385),
.B2(n_386),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_373),
.Y(n_392)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_381),
.B1(n_383),
.B2(n_384),
.Y(n_376)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_381),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_396),
.C(n_397),
.Y(n_395)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_386),
.Y(n_393)
);

NAND4xp25_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_407),
.C(n_414),
.D(n_528),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_394),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_402),
.B1(n_404),
.B2(n_405),
.Y(n_398)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_399),
.Y(n_404)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_400),
.Y(n_401)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_402),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_404),
.C(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_408),
.B(n_410),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_436),
.B(n_527),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_433),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_416),
.B(n_433),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.C(n_422),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_417),
.A2(n_418),
.B1(n_524),
.B2(n_525),
.Y(n_523)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_420),
.B(n_422),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.C(n_429),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_423),
.A2(n_424),
.B1(n_425),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_423),
.Y(n_474)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_429),
.B(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_521),
.B(n_526),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_475),
.B(n_520),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_467),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_439),
.B(n_467),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_456),
.C(n_465),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g485 ( 
.A1(n_440),
.A2(n_441),
.B1(n_486),
.B2(n_488),
.Y(n_485)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_451),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_449),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_449),
.C(n_451),
.Y(n_469)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_456),
.A2(n_465),
.B1(n_466),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_456),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_460),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_457),
.A2(n_458),
.B1(n_460),
.B2(n_461),
.Y(n_478)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_464),
.Y(n_511)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_472),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_469),
.B(n_470),
.C(n_472),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_489),
.B(n_519),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_485),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g519 ( 
.A(n_477),
.B(n_485),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.C(n_483),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_502),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_479),
.A2(n_480),
.B1(n_483),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_483),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_486),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_490),
.A2(n_504),
.B(n_518),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_501),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_491),
.B(n_501),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_499),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_499),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_508),
.B(n_517),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_506),
.B(n_507),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_512),
.Y(n_508)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_522),
.B(n_523),
.Y(n_526)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);


endmodule