module fake_jpeg_8783_n_138 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_18),
.Y(n_52)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_29),
.B1(n_27),
.B2(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_22),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_24),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_19),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_34),
.B1(n_42),
.B2(n_48),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_54),
.A3(n_47),
.B1(n_51),
.B2(n_21),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_67),
.C(n_24),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_32),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_22),
.B(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_84),
.B1(n_59),
.B2(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_44),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_86),
.Y(n_95)
);

AOI21x1_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_15),
.B(n_35),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_72),
.B1(n_65),
.B2(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_23),
.B1(n_45),
.B2(n_42),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_1),
.Y(n_85)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_55),
.B(n_14),
.C(n_26),
.D(n_2),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_90),
.C(n_91),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_69),
.C(n_71),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_59),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_82),
.B(n_85),
.C(n_15),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_96),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_71),
.C(n_55),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_35),
.C(n_45),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_100),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_111),
.B(n_73),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_86),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_98),
.B1(n_76),
.B2(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_115),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_119),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_120),
.B(n_108),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_88),
.B1(n_76),
.B2(n_68),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_108),
.B1(n_15),
.B2(n_26),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_15),
.C(n_20),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_15),
.C(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_119),
.B(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_125),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_4),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.C1(n_11),
.C2(n_13),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_11),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_134),
.B(n_13),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_126),
.C(n_124),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.C(n_5),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_135),
.B(n_2),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_136),
.Y(n_138)
);


endmodule