module real_jpeg_7035_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_2),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_2),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_2),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_2),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_2),
.B(n_31),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_3),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_3),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_78),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_4),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_4),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_4),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_4),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_4),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_5),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_5),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_5),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_5),
.B(n_326),
.Y(n_325)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_6),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_8),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_8),
.B(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_11),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_12),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_12),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_12),
.B(n_93),
.Y(n_227)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_12),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_12),
.B(n_221),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_12),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_13),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_13),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_13),
.B(n_43),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_13),
.B(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_14),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_15),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_15),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_15),
.B(n_93),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_200),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_199),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_158),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_19),
.B(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.C(n_131),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_20),
.A2(n_21),
.B1(n_104),
.B2(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_64),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_22),
.B(n_65),
.C(n_85),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_53),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_23),
.B(n_53),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_30),
.C(n_34),
.Y(n_106)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_28),
.Y(n_168)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_29),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_29),
.Y(n_259)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_38),
.Y(n_192)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_38),
.Y(n_248)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_40),
.B(n_366),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.C(n_49),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_41),
.B(n_45),
.CI(n_49),
.CON(n_133),
.SN(n_133)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g213 ( 
.A(n_44),
.Y(n_213)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_52),
.Y(n_145)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_52),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.C(n_61),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_54),
.A2(n_163),
.B1(n_164),
.B2(n_169),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_54),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_54),
.A2(n_61),
.B1(n_163),
.B2(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_57),
.A2(n_344),
.B1(n_345),
.B2(n_347),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_57),
.Y(n_344)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_60),
.Y(n_218)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_60),
.Y(n_243)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_61),
.Y(n_346)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_63),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_85),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_74),
.C(n_81),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_66),
.B(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_66),
.A2(n_67),
.B(n_70),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_73),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_74),
.B(n_81),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_78),
.Y(n_289)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_79),
.Y(n_266)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_79),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_82),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_82),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_82),
.B(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_98),
.Y(n_85)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_86),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_96),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_87),
.A2(n_96),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_87),
.A2(n_155),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_91),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

OR2x2_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_110),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_126),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_96),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_99),
.B(n_101),
.C(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_104),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_120),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_106),
.B(n_107),
.C(n_120),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_119),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_196),
.C(n_197),
.Y(n_195)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_111),
.Y(n_331)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_123),
.A2(n_124),
.B1(n_135),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_135),
.C(n_138),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_125),
.C(n_129),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_127),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_125),
.A2(n_127),
.B1(n_233),
.B2(n_234),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_127),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_131),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_150),
.C(n_156),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_132),
.B(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.C(n_141),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_133),
.B(n_353),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_133),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_134),
.A2(n_141),
.B1(n_142),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_134),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_135),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_138),
.B(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_314)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_150),
.B(n_156),
.Y(n_362)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_155),
.B(n_245),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_158),
.Y(n_378)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_180),
.CI(n_198),
.CON(n_158),
.SN(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_172),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_170),
.B2(n_171),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_179),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_178),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_178),
.B(n_226),
.C(n_230),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_195),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_357),
.B(n_373),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_335),
.B(n_356),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_304),
.B(n_334),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_261),
.B(n_303),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_249),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_206),
.B(n_249),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_231),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_223),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_208),
.B(n_223),
.C(n_231),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.C(n_219),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_215),
.Y(n_251)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_219),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_232),
.B(n_318),
.C(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_260),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_260),
.B1(n_295),
.B2(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_297),
.B(n_302),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_282),
.B(n_296),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_271),
.B(n_281),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_279),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_279),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B(n_278),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_284),
.B1(n_290),
.B2(n_291),
.Y(n_283)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_292),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_285),
.A2(n_286),
.B(n_290),
.Y(n_298)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B(n_295),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_305),
.B(n_306),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_315),
.B2(n_316),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_317),
.C(n_320),
.Y(n_336)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_313),
.C(n_314),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_333),
.Y(n_320)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_329),
.B2(n_332),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_332),
.C(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

INVx4_ASAP7_75t_SL g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_337),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_350),
.B2(n_355),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_351),
.C(n_352),
.Y(n_367)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_343),
.C(n_348),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_348),
.B2(n_349),
.Y(n_341)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_342),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_350),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_368),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_367),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_367),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_364),
.C(n_365),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_368),
.A2(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_370),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);


endmodule