module fake_jpeg_717_n_599 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_599);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_599;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_1),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_57),
.Y(n_178)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_59),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_65),
.A2(n_46),
.B1(n_50),
.B2(n_44),
.Y(n_137)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_69),
.B(n_76),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_74),
.Y(n_174)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_17),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_114),
.Y(n_128)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_79),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_82),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_83),
.B(n_95),
.Y(n_193)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_88),
.Y(n_201)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_89),
.Y(n_209)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_24),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_94),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_18),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_96),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_98),
.Y(n_218)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_33),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_99),
.B(n_13),
.Y(n_214)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_100),
.Y(n_175)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_0),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_103),
.B(n_9),
.Y(n_206)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

BUFx12f_ASAP7_75t_SL g157 ( 
.A(n_105),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_110),
.Y(n_217)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_117),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_21),
.B(n_0),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_37),
.Y(n_116)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_34),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_29),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

INVx6_ASAP7_75t_SL g188 ( 
.A(n_125),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_130),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_133),
.B(n_147),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_137),
.A2(n_155),
.B1(n_194),
.B2(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_54),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_138),
.B(n_159),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_103),
.A2(n_50),
.B1(n_44),
.B2(n_47),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_143),
.A2(n_181),
.B1(n_182),
.B2(n_186),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_108),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_154),
.B(n_162),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_47),
.B1(n_46),
.B2(n_36),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_69),
.B(n_49),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_118),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_49),
.B1(n_36),
.B2(n_31),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_182),
.B1(n_181),
.B2(n_180),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_165),
.B(n_132),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_76),
.B(n_31),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_169),
.B(n_173),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_29),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_79),
.B(n_15),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_177),
.B(n_204),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_55),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_60),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_65),
.B(n_4),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_185),
.B(n_190),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_64),
.A2(n_72),
.B1(n_96),
.B2(n_70),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_92),
.B(n_4),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_74),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_191),
.A2(n_192),
.B1(n_174),
.B2(n_215),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_80),
.A2(n_88),
.B1(n_87),
.B2(n_82),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_119),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_121),
.B(n_9),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_196),
.A2(n_206),
.B(n_208),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_75),
.B(n_9),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_59),
.B(n_10),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_84),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_57),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_214),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_77),
.B(n_14),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_77),
.B(n_14),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_77),
.B(n_14),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_77),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_77),
.B(n_15),
.C(n_56),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_128),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_224),
.B(n_230),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_156),
.B(n_212),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_225),
.A2(n_250),
.B(n_276),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_155),
.A2(n_168),
.B1(n_216),
.B2(n_199),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_226),
.A2(n_238),
.B1(n_262),
.B2(n_269),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_142),
.B(n_198),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_228),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_126),
.B(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_229),
.Y(n_325)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_141),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_231),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_164),
.A2(n_193),
.B1(n_145),
.B2(n_197),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_232),
.B(n_240),
.Y(n_357)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_233),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_176),
.A2(n_203),
.B1(n_152),
.B2(n_209),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_234),
.A2(n_280),
.B1(n_270),
.B2(n_239),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_158),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_236),
.B(n_245),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_176),
.A2(n_203),
.B1(n_152),
.B2(n_209),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_237),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_163),
.B1(n_127),
.B2(n_136),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_139),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_242),
.Y(n_333)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_150),
.Y(n_243)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_175),
.B(n_129),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_126),
.A2(n_197),
.B(n_131),
.Y(n_250)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_251),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g252 ( 
.A1(n_167),
.A2(n_201),
.B1(n_195),
.B2(n_174),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_144),
.A2(n_184),
.B1(n_195),
.B2(n_200),
.Y(n_253)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_144),
.A2(n_184),
.B1(n_200),
.B2(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_265),
.Y(n_336)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_266),
.Y(n_346)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_187),
.B(n_161),
.CI(n_157),
.CON(n_267),
.SN(n_267)
);

OAI32xp33_ASAP7_75t_L g345 ( 
.A1(n_267),
.A2(n_307),
.A3(n_301),
.B1(n_229),
.B2(n_299),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_187),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_170),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_148),
.Y(n_270)
);

AO22x1_ASAP7_75t_L g271 ( 
.A1(n_134),
.A2(n_135),
.B1(n_145),
.B2(n_140),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_271),
.Y(n_353)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_140),
.Y(n_272)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_283),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_161),
.A2(n_170),
.B(n_218),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_218),
.A2(n_217),
.B1(n_183),
.B2(n_160),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_277),
.A2(n_281),
.B1(n_291),
.B2(n_304),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_151),
.A2(n_215),
.B1(n_166),
.B2(n_167),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_280),
.A2(n_294),
.B1(n_253),
.B2(n_234),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_183),
.A2(n_160),
.B1(n_151),
.B2(n_166),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_149),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_282),
.B(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_149),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_179),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_286),
.Y(n_340)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_202),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_157),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_288),
.Y(n_343)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_178),
.B(n_202),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_292),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_172),
.A2(n_178),
.B1(n_116),
.B2(n_37),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_172),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_187),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_293),
.B(n_308),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_185),
.A2(n_137),
.B1(n_192),
.B2(n_162),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_140),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_296),
.Y(n_359)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_146),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_165),
.B(n_156),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_300),
.C(n_279),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_185),
.A2(n_186),
.B1(n_155),
.B2(n_137),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_298),
.A2(n_302),
.B1(n_235),
.B2(n_225),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_165),
.B(n_156),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_188),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_307),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_155),
.A2(n_185),
.B1(n_143),
.B2(n_186),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_127),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_303),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_133),
.A2(n_116),
.B1(n_37),
.B2(n_99),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_214),
.A2(n_165),
.B(n_223),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_263),
.B(n_244),
.C(n_261),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_188),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_146),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_309),
.A2(n_330),
.B(n_311),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_240),
.B(n_306),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_311),
.B(n_317),
.C(n_318),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_236),
.B1(n_235),
.B2(n_245),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_314),
.A2(n_329),
.B1(n_335),
.B2(n_337),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_224),
.B(n_297),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_300),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_224),
.B(n_300),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_326),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_263),
.B(n_227),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_330),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_241),
.B(n_246),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_324),
.B(n_332),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_258),
.A2(n_248),
.B1(n_274),
.B2(n_305),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_328),
.A2(n_341),
.B(n_249),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_264),
.B(n_228),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_228),
.B(n_258),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_349),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_255),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_230),
.A2(n_294),
.B1(n_232),
.B2(n_281),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_278),
.A2(n_299),
.B1(n_285),
.B2(n_271),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_229),
.B(n_230),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_230),
.A2(n_252),
.B1(n_237),
.B2(n_271),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_350),
.A2(n_361),
.B1(n_273),
.B2(n_295),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_296),
.B(n_308),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_276),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_343),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_362),
.B(n_396),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_313),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_377),
.Y(n_413)
);

AO21x1_ASAP7_75t_L g411 ( 
.A1(n_367),
.A2(n_386),
.B(n_399),
.Y(n_411)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_368),
.Y(n_426)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_369),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_323),
.B(n_285),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_371),
.B(n_383),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_348),
.A2(n_338),
.B(n_353),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_378),
.B(n_403),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_381),
.Y(n_406)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_376),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_342),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_348),
.A2(n_250),
.B(n_278),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_321),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_380),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_359),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_312),
.B(n_260),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_257),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_247),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_385),
.B(n_391),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_267),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_312),
.B(n_314),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_387),
.B(n_402),
.Y(n_438)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_334),
.Y(n_388)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_388),
.Y(n_424)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_389),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_256),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_392),
.Y(n_427)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_393),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_394),
.A2(n_395),
.B1(n_397),
.B2(n_310),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_329),
.A2(n_272),
.B1(n_259),
.B2(n_267),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_284),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_337),
.A2(n_286),
.B1(n_288),
.B2(n_251),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_340),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_401),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_344),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_318),
.B(n_268),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_325),
.B(n_331),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_404),
.Y(n_431)
);

OA21x2_ASAP7_75t_L g405 ( 
.A1(n_372),
.A2(n_320),
.B(n_349),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g443 ( 
.A1(n_405),
.A2(n_373),
.B(n_386),
.C(n_403),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_357),
.C(n_319),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_433),
.Y(n_442)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_415),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_317),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_416),
.B(n_410),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_370),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_417),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_381),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_430),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_365),
.A2(n_320),
.B1(n_328),
.B2(n_335),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_373),
.B1(n_403),
.B2(n_402),
.Y(n_461)
);

AO22x1_ASAP7_75t_SL g430 ( 
.A1(n_365),
.A2(n_320),
.B1(n_350),
.B2(n_322),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_432),
.A2(n_377),
.B1(n_374),
.B2(n_386),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_364),
.B(n_309),
.C(n_326),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_315),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_435),
.B(n_419),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_353),
.B1(n_327),
.B2(n_361),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_436),
.A2(n_440),
.B1(n_397),
.B2(n_395),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_364),
.B(n_367),
.C(n_363),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_364),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_375),
.B(n_345),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_363),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_394),
.A2(n_327),
.B1(n_341),
.B2(n_354),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_384),
.Y(n_441)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_441),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_443),
.A2(n_477),
.B(n_414),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_379),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_444),
.B(n_447),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_445),
.A2(n_428),
.B1(n_436),
.B2(n_440),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_418),
.B(n_362),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_426),
.Y(n_448)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_448),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_411),
.A2(n_399),
.B(n_398),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_450),
.A2(n_451),
.B(n_462),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_425),
.A2(n_398),
.B(n_378),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_452),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_469),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_455),
.A2(n_458),
.B1(n_461),
.B2(n_438),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_421),
.B(n_400),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_456),
.B(n_465),
.Y(n_505)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_457),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_459),
.B(n_467),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_380),
.Y(n_460)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_411),
.A2(n_347),
.B(n_366),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_420),
.B(n_392),
.Y(n_463)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_412),
.B(n_354),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_388),
.Y(n_466)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_466),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_468),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_405),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_408),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_422),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_416),
.B(n_336),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_474),
.Y(n_481)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_423),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_478),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_336),
.C(n_346),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_433),
.B(n_346),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_441),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_425),
.A2(n_369),
.B(n_316),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_423),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_484),
.A2(n_477),
.B1(n_443),
.B2(n_462),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_485),
.Y(n_512)
);

NOR2x1_ASAP7_75t_R g486 ( 
.A(n_443),
.B(n_405),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_492),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_449),
.A2(n_406),
.B1(n_439),
.B2(n_438),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_488),
.A2(n_507),
.B1(n_478),
.B2(n_446),
.Y(n_513)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

INVxp33_ASAP7_75t_L g522 ( 
.A(n_494),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_496),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_430),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_430),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_454),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_463),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_503),
.Y(n_516)
);

A2O1A1O1Ixp25_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_434),
.B(n_427),
.C(n_424),
.D(n_429),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_460),
.Y(n_503)
);

A2O1A1O1Ixp25_ASAP7_75t_L g506 ( 
.A1(n_443),
.A2(n_449),
.B(n_461),
.C(n_451),
.D(n_467),
.Y(n_506)
);

INVxp33_ASAP7_75t_SL g521 ( 
.A(n_506),
.Y(n_521)
);

OAI22xp33_ASAP7_75t_L g507 ( 
.A1(n_458),
.A2(n_427),
.B1(n_424),
.B2(n_431),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_450),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_508),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_408),
.Y(n_509)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_509),
.Y(n_529)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_442),
.C(n_474),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_515),
.B(n_519),
.C(n_527),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_518),
.A2(n_510),
.B1(n_486),
.B2(n_479),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_442),
.C(n_472),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_528),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_473),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_524),
.B(n_531),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_470),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_525),
.B(n_482),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_481),
.B(n_446),
.C(n_457),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_481),
.B(n_452),
.Y(n_528)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_509),
.Y(n_530)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_530),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_496),
.B(n_429),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_497),
.B(n_431),
.C(n_351),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_532),
.B(n_504),
.C(n_483),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_489),
.B(n_414),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_534),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_393),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_489),
.B(n_382),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_479),
.Y(n_547)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_536),
.Y(n_549)
);

CKINVDCx14_ASAP7_75t_R g538 ( 
.A(n_516),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_538),
.B(n_539),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_514),
.B(n_505),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_533),
.Y(n_540)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_540),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_526),
.A2(n_484),
.B1(n_490),
.B2(n_493),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_544),
.A2(n_510),
.B1(n_521),
.B2(n_534),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_522),
.A2(n_487),
.B(n_494),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_545),
.A2(n_551),
.B(n_556),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_529),
.B(n_485),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_548),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_547),
.B(n_553),
.Y(n_559)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_522),
.A2(n_487),
.B(n_506),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_511),
.A2(n_490),
.B1(n_480),
.B2(n_493),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_519),
.B(n_507),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_554),
.B(n_520),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_555),
.B(n_557),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_550),
.Y(n_579)
);

NAND2x1p5_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_523),
.Y(n_562)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_562),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_564),
.A2(n_553),
.B1(n_537),
.B2(n_540),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_549),
.B(n_517),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_565),
.B(n_567),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_545),
.A2(n_532),
.B(n_531),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_566),
.A2(n_568),
.B(n_571),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_552),
.B(n_527),
.C(n_515),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_551),
.A2(n_535),
.B(n_528),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_557),
.B(n_524),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_569),
.B(n_552),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_556),
.A2(n_520),
.B(n_500),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_567),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_577),
.A2(n_581),
.B1(n_582),
.B2(n_566),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_563),
.Y(n_578)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_578),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_542),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_560),
.A2(n_541),
.B(n_548),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_580),
.A2(n_570),
.B(n_564),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_571),
.A2(n_546),
.B1(n_554),
.B2(n_547),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_561),
.A2(n_543),
.B1(n_542),
.B2(n_550),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_583),
.A2(n_589),
.B(n_573),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_584),
.B(n_586),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_575),
.B(n_572),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_587),
.B(n_588),
.C(n_574),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_578),
.A2(n_563),
.B(n_562),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_590),
.B(n_591),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_585),
.A2(n_574),
.B1(n_581),
.B2(n_559),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_593),
.B(n_589),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_595),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_596),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_597),
.B(n_592),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_598),
.A2(n_594),
.B(n_559),
.Y(n_599)
);


endmodule