module real_jpeg_15772_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_125),
.B1(n_128),
.B2(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_1),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_1),
.A2(n_63),
.B1(n_132),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_1),
.A2(n_132),
.B1(n_247),
.B2(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_1),
.A2(n_49),
.B1(n_132),
.B2(n_361),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_2),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_2),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_2),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_3),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_3),
.A2(n_148),
.B1(n_228),
.B2(n_232),
.Y(n_227)
);

AOI22x1_ASAP7_75t_SL g479 ( 
.A1(n_3),
.A2(n_148),
.B1(n_480),
.B2(n_484),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_3),
.A2(n_148),
.B1(n_184),
.B2(n_561),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_195),
.B1(n_196),
.B2(n_203),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_4),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_4),
.A2(n_149),
.B1(n_195),
.B2(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_4),
.A2(n_195),
.B1(n_407),
.B2(n_412),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_4),
.A2(n_184),
.B1(n_195),
.B2(n_526),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g443 ( 
.A1(n_5),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.Y(n_443)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_5),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_5),
.A2(n_446),
.B1(n_509),
.B2(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_6),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g470 ( 
.A(n_6),
.Y(n_470)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_7),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_7),
.Y(n_231)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_7),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_7),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g514 ( 
.A(n_7),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_8),
.A2(n_43),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_8),
.A2(n_43),
.B1(n_407),
.B2(n_523),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_9),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_9),
.A2(n_138),
.B1(n_328),
.B2(n_331),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_9),
.A2(n_138),
.B1(n_319),
.B2(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_9),
.A2(n_138),
.B1(n_423),
.B2(n_427),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_10),
.A2(n_434),
.B1(n_437),
.B2(n_438),
.Y(n_433)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_10),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_10),
.A2(n_437),
.B1(n_509),
.B2(n_510),
.Y(n_508)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_159),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g251 ( 
.A1(n_11),
.A2(n_102),
.A3(n_252),
.B1(n_256),
.B2(n_261),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_11),
.B(n_133),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_11),
.A2(n_28),
.B1(n_273),
.B2(n_360),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_11),
.A2(n_62),
.B1(n_381),
.B2(n_384),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_49),
.B1(n_56),
.B2(n_59),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_12),
.A2(n_59),
.B1(n_451),
.B2(n_455),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_12),
.A2(n_59),
.B1(n_484),
.B2(n_545),
.Y(n_544)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_13),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_14),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_14),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_14),
.A2(n_190),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_14),
.A2(n_190),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_14),
.A2(n_63),
.B1(n_190),
.B2(n_475),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g151 ( 
.A(n_16),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_17),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_534),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_500),
.B(n_532),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_400),
.B(n_497),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_275),
.B(n_399),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_237),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_24),
.B(n_237),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_169),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_90),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_26),
.B(n_90),
.C(n_169),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_60),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_27),
.B(n_60),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_37),
.B1(n_46),
.B2(n_48),
.Y(n_27)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_28),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_28),
.A2(n_314),
.B1(n_321),
.B2(n_322),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_28),
.A2(n_340),
.B1(n_360),
.B2(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_28),
.A2(n_48),
.B1(n_433),
.B2(n_469),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_28),
.A2(n_443),
.B(n_517),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_29),
.Y(n_321)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_31),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_35),
.Y(n_271)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_35),
.Y(n_436)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_36),
.Y(n_286)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_36),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_36),
.Y(n_445)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_38),
.A2(n_143),
.B1(n_152),
.B2(n_153),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_42),
.Y(n_213)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_46),
.Y(n_344)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_54),
.Y(n_440)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_55),
.Y(n_317)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_55),
.Y(n_343)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_77),
.B2(n_83),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_61),
.A2(n_62),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_62),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_62),
.B(n_293),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_62),
.A2(n_292),
.B(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_62),
.B(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_62),
.B(n_236),
.Y(n_370)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_71),
.Y(n_168)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_76),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_76),
.Y(n_418)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_84),
.A2(n_160),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_85),
.Y(n_527)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_86),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_142),
.C(n_158),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_91),
.B(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_123),
.B1(n_133),
.B2(n_134),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_92),
.A2(n_133),
.B1(n_134),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_92),
.A2(n_133),
.B1(n_542),
.B2(n_543),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_93),
.A2(n_124),
.B1(n_380),
.B2(n_386),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_93),
.A2(n_386),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_93),
.A2(n_386),
.B1(n_406),
.B2(n_479),
.Y(n_478)
);

OAI22x1_ASAP7_75t_SL g521 ( 
.A1(n_93),
.A2(n_386),
.B1(n_479),
.B2(n_522),
.Y(n_521)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_102),
.B(n_111),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_109),
.Y(n_260)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_109),
.Y(n_383)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_118),
.B2(n_121),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_113),
.Y(n_284)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_118),
.Y(n_294)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_120),
.Y(n_225)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_120),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_120),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_125),
.Y(n_523)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_128),
.Y(n_385)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_133),
.Y(n_386)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_142),
.B(n_158),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_143),
.A2(n_152),
.B1(n_268),
.B2(n_272),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_150),
.Y(n_320)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_151),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_152),
.A2(n_339),
.B1(n_344),
.B2(n_345),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_152),
.A2(n_432),
.B1(n_441),
.B2(n_442),
.Y(n_431)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_156),
.Y(n_274)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_171),
.B1(n_176),
.B2(n_182),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_159),
.A2(n_176),
.B1(n_182),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_159),
.Y(n_477)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_160),
.A2(n_473),
.B1(n_474),
.B2(n_525),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_160),
.A2(n_473),
.B1(n_525),
.B2(n_560),
.Y(n_559)
);

AOI22x1_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_164),
.B1(n_165),
.B2(n_167),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_186),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_170),
.B(n_187),
.C(n_193),
.Y(n_491)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g473 ( 
.A(n_176),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_185),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_188),
.Y(n_405)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_206),
.B1(n_226),
.B2(n_235),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_198),
.Y(n_509)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_202),
.Y(n_454)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_205),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g330 ( 
.A(n_205),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_206),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_206),
.A2(n_235),
.B1(n_304),
.B2(n_308),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_206),
.A2(n_235),
.B1(n_308),
.B2(n_327),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_206),
.A2(n_235),
.B1(n_244),
.B2(n_327),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_206),
.B(n_460),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g547 ( 
.A1(n_206),
.A2(n_235),
.B1(n_548),
.B2(n_549),
.Y(n_547)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_213),
.Y(n_355)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_224),
.Y(n_217)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_218),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_227),
.A2(n_236),
.B1(n_242),
.B2(n_461),
.Y(n_467)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_235),
.B(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_242),
.B1(n_243),
.B2(n_248),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_236),
.A2(n_242),
.B1(n_450),
.B2(n_508),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.C(n_249),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_238),
.A2(n_239),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_241),
.A2(n_249),
.B1(n_250),
.B2(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_241),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_266),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_251),
.A2(n_266),
.B1(n_267),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_251),
.Y(n_390)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_255),
.Y(n_458)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_392),
.B(n_398),
.Y(n_275)
);

AOI21x1_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_374),
.B(n_391),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_336),
.B(n_373),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_312),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_279),
.B(n_312),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_302),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_280),
.A2(n_302),
.B1(n_303),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_280),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_285),
.A3(n_287),
.B1(n_292),
.B2(n_295),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_323),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_313),
.B(n_325),
.C(n_335),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_314),
.Y(n_345)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_326),
.B2(n_335),
.Y(n_323)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_330),
.Y(n_462)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_348),
.B(n_372),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_346),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_343),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_365),
.B(n_371),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_359),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_356),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_370),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_370),
.Y(n_371)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_368),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_376),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_389),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_387),
.B2(n_388),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_388),
.C(n_389),
.Y(n_397)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_397),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_397),
.Y(n_398)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_486),
.B(n_492),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_401),
.B(n_486),
.C(n_499),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_429),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_402),
.B(n_430),
.C(n_465),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_419),
.C(n_420),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_404),
.B(n_420),
.Y(n_489)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_410),
.Y(n_485)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_410),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_419),
.B(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_422),
.A2(n_473),
.B1(n_474),
.B2(n_477),
.Y(n_472)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_465),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_447),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_431),
.A2(n_448),
.B(n_459),
.Y(n_528)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_459),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx5_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_458),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_471),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_466),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_468),
.Y(n_490)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_478),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_472),
.B(n_478),
.C(n_504),
.Y(n_503)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_490),
.C(n_491),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_487),
.A2(n_488),
.B1(n_495),
.B2(n_496),
.Y(n_494)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_490),
.B(n_491),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_494),
.Y(n_499)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_495),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_531),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g533 ( 
.A(n_502),
.B(n_531),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_505),
.Y(n_502)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_503),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_519),
.B1(n_529),
.B2(n_530),
.Y(n_505)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_506),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_506),
.B(n_530),
.C(n_565),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_507),
.A2(n_515),
.B1(n_516),
.B2(n_518),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_507),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_507),
.B(n_516),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_508),
.Y(n_548)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_515),
.A2(n_516),
.B1(n_558),
.B2(n_559),
.Y(n_557)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_519),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_528),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_528),
.C(n_538),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_524),
.Y(n_538)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_566),
.Y(n_534)
);

NOR2xp67_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_564),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_536),
.B(n_564),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_539),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_555),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_541),
.A2(n_547),
.B(n_554),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_547),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_556),
.A2(n_557),
.B1(n_562),
.B2(n_563),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_562),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);


endmodule