module fake_jpeg_941_n_139 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_14),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_0),
.C(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_13),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_49),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_1),
.B(n_2),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_25),
.B(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_4),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_28),
.A2(n_21),
.B1(n_6),
.B2(n_8),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_67),
.B1(n_46),
.B2(n_36),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_60),
.B1(n_59),
.B2(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_45),
.B1(n_30),
.B2(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_29),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_62),
.B1(n_76),
.B2(n_63),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_74),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_96),
.C(n_75),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_39),
.B1(n_41),
.B2(n_77),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_57),
.B(n_64),
.C(n_68),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_100)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_71),
.B(n_58),
.C(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_69),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_79),
.B(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_99),
.B1(n_107),
.B2(n_105),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_101),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_72),
.B1(n_82),
.B2(n_84),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_104),
.B1(n_87),
.B2(n_99),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_72),
.B1(n_90),
.B2(n_96),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_81),
.B(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_97),
.B(n_106),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_114),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_112),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_100),
.CON(n_111),
.SN(n_111)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_100),
.C(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_124),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_97),
.B(n_102),
.C(n_114),
.D(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_109),
.B1(n_117),
.B2(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_113),
.B1(n_102),
.B2(n_115),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_102),
.B1(n_124),
.B2(n_122),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_132),
.B(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_131),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_130),
.B(n_125),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_135),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_102),
.Y(n_139)
);


endmodule