module fake_jpeg_24066_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_31),
.B1(n_26),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_31),
.B1(n_21),
.B2(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_23),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_58),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_31),
.B1(n_21),
.B2(n_26),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_67),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_31),
.B1(n_21),
.B2(n_26),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_82),
.B1(n_20),
.B2(n_34),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_29),
.B1(n_46),
.B2(n_42),
.Y(n_90)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_70),
.Y(n_93)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_73),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_34),
.C(n_16),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_84),
.C(n_16),
.Y(n_109)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_28),
.B1(n_20),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_78),
.B1(n_49),
.B2(n_42),
.Y(n_103)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_28),
.B1(n_20),
.B2(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NAND2x1p5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_19),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_95),
.B(n_73),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_110),
.B1(n_63),
.B2(n_83),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_16),
.B(n_23),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_18),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_15),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_111),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_63),
.B1(n_81),
.B2(n_75),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_112),
.B1(n_113),
.B2(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_61),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_74),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_33),
.B1(n_32),
.B2(n_28),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_32),
.B1(n_33),
.B2(n_18),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_127),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_99),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_117),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_120),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_119),
.A2(n_114),
.B1(n_96),
.B2(n_107),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_126),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_122),
.C(n_138),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_30),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_111),
.B1(n_87),
.B2(n_100),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_131),
.B(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_30),
.B1(n_17),
.B2(n_25),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_114),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_135),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_30),
.B1(n_17),
.B2(n_25),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_17),
.B1(n_22),
.B2(n_48),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_24),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_38),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_142),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_22),
.Y(n_142)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_148),
.Y(n_194)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_108),
.B(n_89),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_162),
.B(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_152),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_171),
.C(n_172),
.Y(n_188)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_89),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_91),
.Y(n_159)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_164),
.B1(n_170),
.B2(n_173),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_91),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_66),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_159),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_158),
.B1(n_157),
.B2(n_165),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_140),
.C(n_117),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_92),
.C(n_104),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_88),
.B1(n_100),
.B2(n_104),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_116),
.B(n_106),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_176),
.A2(n_181),
.B(n_198),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_197),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_115),
.B1(n_134),
.B2(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_189),
.B1(n_199),
.B2(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_106),
.B1(n_107),
.B2(n_66),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_186),
.B1(n_200),
.B2(n_146),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_0),
.B(n_1),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_185),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_38),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_48),
.B1(n_56),
.B2(n_60),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_48),
.B1(n_24),
.B2(n_15),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_151),
.B1(n_148),
.B2(n_27),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_40),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_193),
.C(n_195),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_40),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_40),
.C(n_39),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_144),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_0),
.B(n_1),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_24),
.B1(n_27),
.B2(n_15),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_15),
.B1(n_27),
.B2(n_2),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_143),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_206),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_39),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_39),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_38),
.C(n_37),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_175),
.B(n_143),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_211),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_207),
.B(n_150),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_213),
.B(n_229),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_184),
.B(n_151),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_193),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_187),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_226),
.B1(n_227),
.B2(n_205),
.Y(n_242)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_231),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_195),
.B1(n_206),
.B2(n_178),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_188),
.A2(n_199),
.B1(n_192),
.B2(n_202),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_8),
.B(n_14),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_185),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_238),
.Y(n_268)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_245),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_217),
.B1(n_227),
.B2(n_208),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_181),
.C(n_204),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_223),
.C(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_0),
.Y(n_244)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_231),
.B1(n_211),
.B2(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_250),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_221),
.A2(n_3),
.B(n_4),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_251),
.B(n_11),
.Y(n_262)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_212),
.A2(n_9),
.B(n_13),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_257),
.A2(n_258),
.B1(n_262),
.B2(n_246),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_245),
.B(n_209),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_263),
.C(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_230),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_226),
.B1(n_218),
.B2(n_10),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_237),
.B1(n_10),
.B2(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_240),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.C(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_37),
.C(n_5),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_234),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_275),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_236),
.B1(n_233),
.B2(n_235),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_279),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_242),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_280),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_241),
.C(n_232),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_278),
.B(n_261),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_287),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_257),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_261),
.B(n_265),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_293),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_266),
.B(n_263),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_291),
.B(n_270),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_252),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_269),
.A2(n_262),
.B(n_267),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_295),
.B(n_298),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_282),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_288),
.A2(n_281),
.B1(n_252),
.B2(n_276),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_301),
.B1(n_284),
.B2(n_3),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_272),
.B(n_256),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_284),
.B(n_9),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_7),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_7),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_283),
.C(n_287),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_308),
.C(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_297),
.C(n_10),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_307),
.B(n_301),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_309),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

AOI321xp33_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_310),
.A3(n_311),
.B1(n_304),
.B2(n_9),
.C(n_13),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_314),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_13),
.B(n_37),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);


endmodule