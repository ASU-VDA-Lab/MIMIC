module fake_jpeg_26271_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

INVx13_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

AOI22xp5_ASAP7_75t_L g8 ( 
.A1(n_4),
.A2(n_1),
.B1(n_0),
.B2(n_5),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_5),
.B(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx4_ASAP7_75t_SL g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_4),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_16),
.B(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_13),
.Y(n_17)
);

OR2x4_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_11),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_19),
.B1(n_21),
.B2(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_6),
.B(n_10),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_11),
.Y(n_23)
);

FAx1_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_27),
.CI(n_28),
.CON(n_31),
.SN(n_31)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_17),
.C(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_18),
.B1(n_28),
.B2(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_33),
.B(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_31),
.Y(n_36)
);


endmodule