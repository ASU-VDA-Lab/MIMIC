module fake_netlist_6_193_n_1771 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1771);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1771;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_79),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_14),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_48),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_25),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_160),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_139),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_65),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_31),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_66),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_123),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_32),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_109),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_80),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_97),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_104),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_88),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_6),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_43),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_99),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_96),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_22),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_70),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_58),
.Y(n_205)
);

BUFx8_ASAP7_75t_SL g206 ( 
.A(n_17),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_37),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_124),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_74),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_4),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_158),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_0),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_115),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_26),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_85),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_147),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_111),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_20),
.Y(n_222)
);

INVx4_ASAP7_75t_R g223 ( 
.A(n_132),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_35),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_42),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_93),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_51),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_62),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_59),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_24),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_69),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_7),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_113),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_13),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_103),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_7),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_22),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_16),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_64),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_72),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_153),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_43),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_27),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_30),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_8),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_29),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_101),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_116),
.Y(n_251)
);

BUFx2_ASAP7_75t_SL g252 ( 
.A(n_91),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_68),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_73),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_6),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_95),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_129),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_21),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_4),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_86),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_46),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_19),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_81),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_84),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_140),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_16),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_110),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_49),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_10),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_57),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_40),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_3),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_41),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_98),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_27),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_83),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_15),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_151),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_29),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_5),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_2),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_122),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_12),
.Y(n_286)
);

INVxp33_ASAP7_75t_R g287 ( 
.A(n_114),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_23),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_100),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_3),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_155),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_78),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_50),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_44),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_45),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_0),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_15),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_107),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_2),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_148),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_71),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_14),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_76),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_23),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_19),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_108),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_157),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_117),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_41),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_120),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_127),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_37),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_55),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_39),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_30),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_11),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_92),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_128),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_18),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_36),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_144),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_47),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_18),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_44),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_135),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_137),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_165),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_167),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_175),
.B(n_1),
.Y(n_330)
);

BUFx6f_ASAP7_75t_SL g331 ( 
.A(n_271),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_206),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_309),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_183),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_239),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_178),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_183),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_248),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_271),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_239),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_249),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_249),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_249),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_185),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_214),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_249),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_249),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_274),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_304),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_274),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_168),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_193),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_238),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_274),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_207),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_253),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_238),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_217),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_225),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_237),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_264),
.Y(n_363)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_174),
.B(n_1),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_278),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_200),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_221),
.B(n_5),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_202),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_221),
.B(n_8),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_211),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_264),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_172),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_221),
.B(n_9),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_181),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_188),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_189),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_191),
.Y(n_384)
);

BUFx6f_ASAP7_75t_SL g385 ( 
.A(n_271),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_205),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_213),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_222),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_216),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_220),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_224),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_230),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_240),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_241),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_243),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_245),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_247),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_166),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_261),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_232),
.B(n_9),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_258),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_262),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_227),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_232),
.B(n_10),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_228),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_266),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_268),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_285),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_184),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_332),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_328),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_332),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_329),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_333),
.B(n_198),
.Y(n_416)
);

CKINVDCx8_ASAP7_75t_R g417 ( 
.A(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_343),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_345),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_353),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_349),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_353),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_379),
.A2(n_382),
.B(n_381),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_368),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_336),
.B(n_234),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_333),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_368),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_334),
.B(n_296),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_331),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_354),
.B(n_233),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_350),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_337),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g446 ( 
.A(n_331),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_344),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_341),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_370),
.B(n_253),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_342),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_351),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_355),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_403),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_356),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_359),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_363),
.B(n_296),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_374),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_402),
.B(n_233),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_409),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_371),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_409),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_405),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_357),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_331),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_380),
.B(n_251),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_383),
.B(n_251),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_372),
.B(n_319),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_408),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_407),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_339),
.Y(n_477)
);

BUFx8_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_377),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_373),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_360),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_373),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_376),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_451),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_420),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_415),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_435),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_338),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_439),
.B(n_460),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_443),
.B(n_376),
.Y(n_493)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_473),
.B(n_208),
.Y(n_494)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_438),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_428),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_435),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_439),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_473),
.B(n_319),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_460),
.B(n_388),
.Y(n_500)
);

BUFx8_ASAP7_75t_SL g501 ( 
.A(n_449),
.Y(n_501)
);

BUFx10_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_481),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_388),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_473),
.B(n_253),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_398),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_420),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_411),
.B(n_398),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_411),
.B(n_445),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_413),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_411),
.B(n_335),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_412),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_481),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_466),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_445),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

BUFx4f_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

INVx4_ASAP7_75t_SL g521 ( 
.A(n_451),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_479),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_445),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_479),
.B(n_253),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_462),
.B(n_391),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_433),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_447),
.B(n_391),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_480),
.B(n_393),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_466),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_L g532 ( 
.A(n_451),
.B(n_393),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_425),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_451),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_466),
.Y(n_536)
);

CKINVDCx11_ASAP7_75t_R g537 ( 
.A(n_417),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_421),
.B(n_287),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_423),
.A2(n_330),
.B1(n_394),
.B2(n_401),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_456),
.Y(n_540)
);

BUFx4f_ASAP7_75t_L g541 ( 
.A(n_447),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_479),
.B(n_253),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_463),
.B(n_340),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_477),
.B(n_293),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_476),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_433),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_436),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_425),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_463),
.B(n_361),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_476),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_468),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_422),
.B(n_394),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_476),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_476),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_436),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_476),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_425),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_441),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_476),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_424),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_479),
.B(n_236),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_437),
.B(n_396),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_479),
.B(n_386),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_471),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_465),
.B(n_362),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_475),
.B(n_396),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_479),
.B(n_397),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_425),
.Y(n_574)
);

INVx4_ASAP7_75t_SL g575 ( 
.A(n_451),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_451),
.A2(n_404),
.B1(n_400),
.B2(n_184),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_475),
.B(n_397),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_475),
.B(n_401),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_451),
.B(n_387),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_452),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_452),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_422),
.B(n_365),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_437),
.B(n_364),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_475),
.B(n_289),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_426),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_467),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_418),
.Y(n_587)
);

INVx8_ASAP7_75t_L g588 ( 
.A(n_432),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_446),
.B(n_292),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_464),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_452),
.Y(n_592)
);

BUFx8_ASAP7_75t_SL g593 ( 
.A(n_482),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_410),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_418),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_450),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_455),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_419),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_472),
.B(n_352),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_455),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_457),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_452),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_457),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_483),
.A2(n_298),
.B1(n_385),
.B2(n_176),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_L g605 ( 
.A(n_467),
.B(n_164),
.Y(n_605)
);

AND2x6_ASAP7_75t_L g606 ( 
.A(n_419),
.B(n_303),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_440),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_430),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_452),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_452),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_430),
.B(n_308),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_453),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_434),
.B(n_389),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_453),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_448),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_446),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_434),
.B(n_390),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_442),
.B(n_392),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_465),
.B(n_366),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_442),
.B(n_395),
.Y(n_621)
);

BUFx4f_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_440),
.B(n_166),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_444),
.B(n_399),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_444),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_467),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_474),
.B(n_385),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_448),
.B(n_454),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_448),
.B(n_406),
.Y(n_629)
);

NAND2x1p5_ASAP7_75t_L g630 ( 
.A(n_474),
.B(n_310),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_446),
.B(n_311),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_446),
.B(n_367),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_498),
.A2(n_235),
.B1(n_195),
.B2(n_196),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_586),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_501),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_484),
.B(n_313),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_526),
.B(n_417),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_583),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_494),
.B(n_526),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_L g640 ( 
.A(n_554),
.B(n_440),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_492),
.A2(n_326),
.B(n_315),
.C(n_474),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_494),
.B(n_470),
.Y(n_642)
);

O2A1O1Ixp5_ASAP7_75t_L g643 ( 
.A1(n_491),
.A2(n_458),
.B(n_454),
.C(n_448),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_500),
.B(n_470),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_489),
.B(n_199),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_569),
.B(n_454),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_493),
.B(n_231),
.Y(n_647)
);

AO221x1_ASAP7_75t_L g648 ( 
.A1(n_517),
.A2(n_194),
.B1(n_260),
.B2(n_369),
.C(n_223),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_507),
.B(n_478),
.C(n_440),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_491),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_507),
.B(n_246),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_569),
.A2(n_458),
.B(n_454),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_571),
.B(n_458),
.Y(n_653)
);

AND2x2_ASAP7_75t_SL g654 ( 
.A(n_576),
.B(n_194),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_571),
.B(n_263),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_616),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_616),
.Y(n_657)
);

AND3x1_ASAP7_75t_L g658 ( 
.A(n_528),
.B(n_260),
.C(n_321),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_576),
.A2(n_164),
.B1(n_187),
.B2(n_186),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_577),
.B(n_458),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_496),
.A2(n_410),
.B(n_427),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_498),
.A2(n_218),
.B1(n_190),
.B2(n_192),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_577),
.B(n_586),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_488),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_498),
.B(n_410),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_513),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_498),
.A2(n_219),
.B1(n_197),
.B2(n_201),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_498),
.B(n_427),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_513),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_599),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_505),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_578),
.B(n_530),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_509),
.B(n_470),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_566),
.A2(n_187),
.B1(n_186),
.B2(n_182),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_587),
.B(n_427),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_578),
.B(n_267),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_490),
.A2(n_226),
.B(n_265),
.C(n_259),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_503),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_566),
.A2(n_212),
.B1(n_203),
.B2(n_204),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_530),
.B(n_539),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_509),
.B(n_470),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_567),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_496),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_518),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_495),
.B(n_255),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_632),
.B(n_582),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_499),
.A2(n_327),
.B1(n_252),
.B2(n_305),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_582),
.A2(n_536),
.B1(n_531),
.B2(n_587),
.Y(n_688)
);

INVx6_ASAP7_75t_L g689 ( 
.A(n_510),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_531),
.B(n_169),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_625),
.B(n_429),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_516),
.A2(n_210),
.B(n_256),
.C(n_254),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_572),
.B(n_169),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_591),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_572),
.B(n_518),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_495),
.B(n_478),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_596),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_484),
.B(n_327),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_597),
.B(n_429),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_486),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_540),
.Y(n_702)
);

BUFx8_ASAP7_75t_L g703 ( 
.A(n_585),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_499),
.A2(n_327),
.B1(n_305),
.B2(n_312),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_600),
.B(n_429),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_601),
.B(n_453),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_603),
.B(n_453),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_487),
.B(n_180),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_497),
.B(n_180),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_520),
.B(n_478),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_595),
.B(n_209),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_595),
.B(n_229),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_598),
.B(n_242),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_551),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_524),
.B(n_478),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_598),
.B(n_608),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_520),
.B(n_270),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_608),
.B(n_244),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_551),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_541),
.B(n_272),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_541),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_626),
.B(n_257),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_579),
.A2(n_291),
.B(n_269),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_627),
.B(n_275),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_570),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_604),
.B(n_170),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_627),
.B(n_277),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_553),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_629),
.B(n_485),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_544),
.B(n_170),
.Y(n_730)
);

INVx8_ASAP7_75t_L g731 ( 
.A(n_588),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_504),
.A2(n_301),
.B1(n_300),
.B2(n_281),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_565),
.A2(n_320),
.B1(n_316),
.B2(n_324),
.Y(n_733)
);

NOR2x1_ASAP7_75t_L g734 ( 
.A(n_589),
.B(n_250),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_580),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_570),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_511),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_485),
.B(n_171),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_620),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_546),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_620),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_502),
.B(n_171),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_515),
.B(n_173),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_544),
.B(n_623),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_613),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_532),
.A2(n_173),
.B(n_176),
.C(n_177),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_617),
.B(n_177),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_502),
.B(n_589),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_618),
.A2(n_280),
.B1(n_273),
.B2(n_282),
.C(n_283),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_515),
.B(n_179),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_484),
.B(n_179),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_512),
.B(n_302),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_606),
.A2(n_327),
.B1(n_325),
.B2(n_324),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_484),
.B(n_182),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_590),
.B(n_279),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_631),
.A2(n_605),
.B1(n_606),
.B2(n_611),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_508),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_522),
.B(n_306),
.Y(n_758)
);

BUFx5_ASAP7_75t_L g759 ( 
.A(n_606),
.Y(n_759)
);

INVx5_ASAP7_75t_L g760 ( 
.A(n_606),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_619),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_522),
.B(n_306),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_535),
.B(n_307),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_538),
.B(n_325),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_580),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_631),
.B(n_322),
.C(n_307),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_529),
.B(n_534),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_527),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_529),
.B(n_323),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_527),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_628),
.A2(n_322),
.B(n_323),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_535),
.B(n_279),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_584),
.A2(n_295),
.B(n_288),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_545),
.B(n_297),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_621),
.B(n_294),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_534),
.B(n_327),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_624),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_593),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_542),
.B(n_299),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_548),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_535),
.B(n_279),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_535),
.B(n_318),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_SL g783 ( 
.A(n_630),
.B(n_312),
.C(n_316),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_521),
.B(n_318),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_549),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_549),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_514),
.B(n_290),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_521),
.B(n_318),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_555),
.B(n_286),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_558),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_588),
.Y(n_791)
);

INVxp33_ASAP7_75t_L g792 ( 
.A(n_537),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_559),
.Y(n_793)
);

AOI21x1_ASAP7_75t_L g794 ( 
.A1(n_652),
.A2(n_557),
.B(n_560),
.Y(n_794)
);

INVx11_ASAP7_75t_L g795 ( 
.A(n_703),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_752),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_646),
.A2(n_622),
.B(n_615),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_701),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_661),
.A2(n_622),
.B(n_615),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_680),
.A2(n_611),
.B1(n_606),
.B2(n_584),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_663),
.B(n_611),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_650),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_655),
.B(n_745),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_643),
.A2(n_556),
.B(n_547),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_672),
.B(n_568),
.C(n_525),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_653),
.A2(n_592),
.B(n_602),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_698),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_655),
.A2(n_525),
.B(n_543),
.C(n_630),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_757),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_698),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_672),
.B(n_514),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_683),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_702),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_728),
.Y(n_814)
);

OA21x2_ASAP7_75t_L g815 ( 
.A1(n_643),
.A2(n_564),
.B(n_552),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_660),
.A2(n_592),
.B(n_602),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_740),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_635),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_761),
.B(n_611),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_665),
.A2(n_523),
.B(n_561),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_638),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_SL g822 ( 
.A1(n_637),
.A2(n_538),
.B1(n_320),
.B2(n_284),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_639),
.B(n_533),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_651),
.B(n_537),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_716),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_664),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_L g827 ( 
.A(n_759),
.B(n_588),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_668),
.A2(n_523),
.B(n_550),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_760),
.B(n_614),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_651),
.B(n_533),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_689),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_654),
.A2(n_607),
.B1(n_594),
.B2(n_543),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_654),
.A2(n_563),
.B(n_559),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_682),
.B(n_538),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_683),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_729),
.A2(n_561),
.B(n_550),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_757),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_652),
.A2(n_573),
.B(n_562),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_671),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_676),
.A2(n_573),
.B(n_562),
.C(n_563),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_689),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_675),
.A2(n_561),
.B(n_508),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_777),
.B(n_611),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_746),
.A2(n_574),
.B(n_555),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_682),
.B(n_574),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_775),
.B(n_506),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_670),
.B(n_521),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_647),
.B(n_561),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_647),
.B(n_686),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_767),
.A2(n_508),
.B(n_519),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_735),
.A2(n_508),
.B(n_519),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_688),
.A2(n_506),
.B(n_612),
.Y(n_852)
);

OAI21xp33_ASAP7_75t_L g853 ( 
.A1(n_676),
.A2(n_614),
.B(n_610),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_735),
.A2(n_519),
.B(n_550),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_695),
.A2(n_689),
.B1(n_693),
.B2(n_756),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_693),
.A2(n_614),
.B(n_580),
.C(n_610),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_L g857 ( 
.A(n_774),
.B(n_726),
.C(n_685),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_765),
.A2(n_519),
.B(n_550),
.Y(n_858)
);

AOI221x1_ASAP7_75t_L g859 ( 
.A1(n_641),
.A2(n_614),
.B1(n_580),
.B2(n_610),
.C(n_609),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_775),
.B(n_506),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_659),
.A2(n_634),
.B(n_677),
.C(n_692),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_695),
.A2(n_506),
.B1(n_575),
.B2(n_609),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_SL g863 ( 
.A(n_755),
.B(n_506),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_638),
.B(n_609),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_645),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_757),
.Y(n_866)
);

BUFx12f_ASAP7_75t_L g867 ( 
.A(n_703),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_666),
.Y(n_868)
);

O2A1O1Ixp5_ASAP7_75t_L g869 ( 
.A1(n_723),
.A2(n_575),
.B(n_610),
.C(n_609),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_765),
.A2(n_612),
.B(n_581),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_678),
.B(n_694),
.Y(n_871)
);

AND2x6_ASAP7_75t_L g872 ( 
.A(n_734),
.B(n_575),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_717),
.B(n_11),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_760),
.A2(n_612),
.B(n_581),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_697),
.B(n_612),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_760),
.A2(n_581),
.B(n_56),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_753),
.A2(n_581),
.B(n_67),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_731),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_760),
.A2(n_54),
.B(n_152),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_681),
.B(n_690),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_742),
.B(n_12),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_SL g882 ( 
.A1(n_784),
.A2(n_13),
.B(n_21),
.C(n_24),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_690),
.B(n_724),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_742),
.B(n_28),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_726),
.A2(n_28),
.B(n_33),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_727),
.B(n_33),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_706),
.A2(n_82),
.B(n_149),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_748),
.B(n_34),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_748),
.A2(n_75),
.B1(n_146),
.B2(n_145),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_753),
.A2(n_53),
.B(n_141),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_766),
.B(n_52),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_723),
.A2(n_780),
.B(n_786),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_707),
.A2(n_691),
.B(n_700),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_705),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_714),
.B(n_34),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_633),
.A2(n_87),
.B1(n_119),
.B2(n_106),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_720),
.B(n_35),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_708),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_779),
.A2(n_789),
.B(n_699),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_657),
.A2(n_161),
.B(n_105),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_711),
.A2(n_94),
.B(n_89),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_709),
.B(n_36),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_719),
.B(n_38),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_725),
.A2(n_45),
.B(n_39),
.C(n_40),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_736),
.A2(n_38),
.B(n_42),
.C(n_739),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_712),
.A2(n_713),
.B(n_718),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_738),
.A2(n_750),
.B(n_769),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_737),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_741),
.B(n_684),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_766),
.A2(n_687),
.B(n_771),
.C(n_704),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_684),
.B(n_687),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_731),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_L g913 ( 
.A(n_759),
.B(n_791),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_662),
.A2(n_667),
.B1(n_669),
.B2(n_642),
.Y(n_914)
);

NAND3xp33_ASAP7_75t_L g915 ( 
.A(n_704),
.B(n_771),
.C(n_749),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_743),
.A2(n_758),
.B(n_762),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_673),
.A2(n_732),
.B1(n_644),
.B2(n_715),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_731),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_722),
.A2(n_776),
.B(n_790),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_744),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_768),
.A2(n_793),
.B(n_770),
.Y(n_921)
);

NAND3xp33_ASAP7_75t_L g922 ( 
.A(n_658),
.B(n_773),
.C(n_679),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_785),
.A2(n_788),
.B(n_754),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_751),
.A2(n_763),
.B(n_636),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_636),
.A2(n_781),
.B(n_782),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_730),
.B(n_787),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_730),
.B(n_759),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_772),
.A2(n_747),
.B(n_744),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_648),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_773),
.A2(n_783),
.B(n_674),
.C(n_649),
.Y(n_930)
);

BUFx4f_ASAP7_75t_L g931 ( 
.A(n_764),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_783),
.A2(n_710),
.B(n_696),
.C(n_640),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_759),
.A2(n_733),
.B(n_792),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_733),
.A2(n_672),
.B1(n_655),
.B2(n_663),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_759),
.A2(n_646),
.B(n_661),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_759),
.A2(n_680),
.B1(n_639),
.B2(n_672),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_778),
.B(n_569),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_643),
.A2(n_661),
.B(n_654),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_650),
.Y(n_939)
);

INVx6_ASAP7_75t_L g940 ( 
.A(n_703),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_646),
.A2(n_661),
.B(n_660),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_651),
.B(n_670),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_716),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_637),
.B(n_672),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_716),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_651),
.B(n_670),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_637),
.B(n_672),
.Y(n_947)
);

NOR2xp67_ASAP7_75t_L g948 ( 
.A(n_721),
.B(n_617),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_651),
.B(n_670),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_757),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_637),
.B(n_672),
.Y(n_951)
);

AOI22x1_ASAP7_75t_L g952 ( 
.A1(n_650),
.A2(n_683),
.B1(n_657),
.B2(n_656),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_672),
.B(n_637),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_646),
.A2(n_661),
.B(n_660),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_672),
.A2(n_655),
.B(n_680),
.C(n_676),
.Y(n_955)
);

BUFx4f_ASAP7_75t_L g956 ( 
.A(n_731),
.Y(n_956)
);

BUFx4f_ASAP7_75t_L g957 ( 
.A(n_731),
.Y(n_957)
);

OAI21xp33_ASAP7_75t_L g958 ( 
.A1(n_651),
.A2(n_655),
.B(n_647),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_672),
.B(n_637),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_701),
.Y(n_960)
);

OAI321xp33_ASAP7_75t_L g961 ( 
.A1(n_655),
.A2(n_651),
.A3(n_680),
.B1(n_672),
.B2(n_637),
.C(n_676),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_740),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_646),
.A2(n_661),
.B(n_660),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_SL g964 ( 
.A1(n_746),
.A2(n_641),
.B(n_639),
.C(n_677),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_646),
.A2(n_661),
.B(n_660),
.Y(n_965)
);

AO21x1_ASAP7_75t_L g966 ( 
.A1(n_672),
.A2(n_639),
.B(n_655),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_637),
.B(n_672),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_646),
.A2(n_661),
.B(n_660),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_716),
.Y(n_969)
);

INVx11_ASAP7_75t_L g970 ( 
.A(n_703),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_638),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_650),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_757),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_802),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_955),
.A2(n_938),
.B(n_961),
.Y(n_975)
);

AOI21x1_ASAP7_75t_SL g976 ( 
.A1(n_911),
.A2(n_886),
.B(n_860),
.Y(n_976)
);

AO31x2_ASAP7_75t_L g977 ( 
.A1(n_859),
.A2(n_856),
.A3(n_966),
.B(n_855),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_826),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_942),
.B(n_946),
.Y(n_980)
);

BUFx12f_ASAP7_75t_L g981 ( 
.A(n_867),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_812),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_835),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_804),
.A2(n_919),
.B(n_836),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_804),
.A2(n_850),
.B(n_842),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_949),
.B(n_944),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_947),
.B(n_951),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_963),
.A2(n_968),
.B(n_965),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_967),
.B(n_803),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_958),
.A2(n_961),
.B(n_849),
.C(n_888),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_938),
.A2(n_936),
.B(n_877),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_935),
.A2(n_801),
.B(n_893),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_877),
.A2(n_881),
.B(n_884),
.C(n_934),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_880),
.A2(n_953),
.B(n_959),
.C(n_890),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_821),
.Y(n_996)
);

NAND2x1p5_ASAP7_75t_L g997 ( 
.A(n_878),
.B(n_912),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_830),
.B(n_865),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_825),
.B(n_943),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_813),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_885),
.A2(n_910),
.B(n_796),
.C(n_857),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_890),
.A2(n_861),
.B(n_883),
.C(n_915),
.Y(n_1002)
);

BUFx2_ASAP7_75t_R g1003 ( 
.A(n_818),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_833),
.A2(n_915),
.B(n_805),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_899),
.A2(n_869),
.B(n_828),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_833),
.A2(n_805),
.B(n_840),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_821),
.B(n_971),
.Y(n_1007)
);

AOI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_922),
.A2(n_914),
.B(n_873),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_918),
.B(n_831),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_922),
.A2(n_906),
.B(n_800),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_907),
.A2(n_916),
.B(n_806),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_816),
.A2(n_797),
.B(n_820),
.Y(n_1012)
);

BUFx2_ASAP7_75t_SL g1013 ( 
.A(n_798),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_892),
.A2(n_844),
.B(n_923),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_971),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_945),
.A2(n_969),
.B(n_819),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_848),
.B(n_894),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_898),
.B(n_824),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_SL g1019 ( 
.A(n_918),
.B(n_878),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_851),
.A2(n_858),
.B(n_854),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_921),
.A2(n_924),
.B(n_815),
.Y(n_1021)
);

AO31x2_ASAP7_75t_L g1022 ( 
.A1(n_929),
.A2(n_930),
.A3(n_846),
.B(n_832),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_871),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_SL g1024 ( 
.A1(n_928),
.A2(n_843),
.B(n_933),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_815),
.A2(n_829),
.B(n_870),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_808),
.A2(n_852),
.B(n_964),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_845),
.B(n_897),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_926),
.B(n_807),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_898),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_795),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_852),
.A2(n_891),
.B(n_927),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_864),
.B(n_810),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_939),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_913),
.A2(n_827),
.B(n_853),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_810),
.B(n_908),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_811),
.A2(n_917),
.B1(n_834),
.B2(n_823),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_831),
.B(n_841),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_817),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_841),
.B(n_909),
.Y(n_1039)
);

AOI21xp33_ASAP7_75t_L g1040 ( 
.A1(n_895),
.A2(n_903),
.B(n_863),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_829),
.A2(n_874),
.B(n_925),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_972),
.A2(n_875),
.B(n_876),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_932),
.A2(n_862),
.B1(n_889),
.B2(n_905),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_847),
.B(n_839),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_900),
.A2(n_901),
.B(n_887),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_918),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_879),
.A2(n_896),
.B(n_948),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_872),
.A2(n_902),
.B(n_973),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_904),
.A2(n_863),
.B(n_872),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_872),
.A2(n_809),
.B(n_950),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_962),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_809),
.A2(n_973),
.B(n_837),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_809),
.B(n_973),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_920),
.A2(n_931),
.B(n_937),
.C(n_956),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_872),
.A2(n_950),
.B(n_866),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_837),
.A2(n_950),
.B(n_866),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_912),
.B(n_868),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_931),
.B(n_868),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_814),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_920),
.A2(n_957),
.B1(n_956),
.B2(n_822),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_868),
.B(n_960),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_882),
.A2(n_957),
.B(n_970),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_940),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_940),
.A2(n_799),
.B(n_941),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_955),
.A2(n_938),
.B(n_961),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_798),
.B(n_731),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_813),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_898),
.B(n_413),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_798),
.B(n_731),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_955),
.A2(n_938),
.B(n_961),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_918),
.B(n_831),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_799),
.A2(n_935),
.B(n_801),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_813),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_944),
.B(n_947),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_944),
.B(n_947),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_859),
.A2(n_856),
.A3(n_966),
.B(n_855),
.Y(n_1084)
);

AOI21x1_ASAP7_75t_L g1085 ( 
.A1(n_799),
.A2(n_935),
.B(n_801),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_817),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_859),
.A2(n_856),
.A3(n_966),
.B(n_855),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_944),
.B(n_951),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_944),
.A2(n_947),
.B1(n_951),
.B2(n_967),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_L g1093 ( 
.A(n_958),
.B(n_955),
.C(n_947),
.Y(n_1093)
);

AO21x1_ASAP7_75t_L g1094 ( 
.A1(n_944),
.A2(n_947),
.B(n_951),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_878),
.B(n_912),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_944),
.A2(n_947),
.B1(n_951),
.B2(n_967),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_799),
.A2(n_935),
.B(n_801),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_944),
.B(n_947),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_SL g1099 ( 
.A1(n_944),
.A2(n_680),
.B(n_637),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_944),
.B(n_951),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_799),
.A2(n_935),
.B(n_801),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_826),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_809),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_794),
.A2(n_838),
.B(n_952),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_944),
.B(n_947),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_SL g1108 ( 
.A1(n_911),
.A2(n_886),
.B(n_860),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_944),
.A2(n_947),
.B1(n_951),
.B2(n_967),
.Y(n_1109)
);

BUFx2_ASAP7_75t_SL g1110 ( 
.A(n_798),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_821),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_826),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_944),
.B(n_947),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_799),
.A2(n_954),
.B(n_941),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_944),
.B(n_947),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_955),
.A2(n_938),
.B(n_961),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_944),
.B(n_947),
.Y(n_1117)
);

BUFx4f_ASAP7_75t_L g1118 ( 
.A(n_918),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1118),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_978),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1103),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1038),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_988),
.A2(n_1107),
.B1(n_1083),
.B2(n_1117),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1034),
.A2(n_1011),
.B(n_1002),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1010),
.A2(n_1067),
.B(n_979),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_1069),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1010),
.A2(n_1072),
.B(n_1070),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1118),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1092),
.A2(n_1096),
.B1(n_1109),
.B2(n_1115),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_987),
.B(n_980),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_1068),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1057),
.B(n_1058),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1086),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_997),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1112),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1080),
.B(n_1113),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1098),
.B(n_990),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_1061),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1078),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1092),
.A2(n_1096),
.B1(n_1109),
.B2(n_1098),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1068),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1057),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1018),
.B(n_998),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_999),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1093),
.A2(n_1008),
.B1(n_1094),
.B2(n_975),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_974),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1099),
.B(n_1023),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_994),
.A2(n_975),
.B(n_1075),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1017),
.B(n_995),
.Y(n_1150)
);

BUFx12f_ASAP7_75t_L g1151 ( 
.A(n_981),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1027),
.B(n_991),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1015),
.B(n_1111),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1095),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1068),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1015),
.B(n_1111),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1003),
.B(n_1060),
.Y(n_1157)
);

INVx5_ASAP7_75t_L g1158 ( 
.A(n_1073),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1051),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1095),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_996),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1029),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1028),
.B(n_1036),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_992),
.A2(n_1116),
.B1(n_1065),
.B2(n_1075),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1009),
.B(n_1076),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1029),
.B(n_1007),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1001),
.B(n_1039),
.Y(n_1167)
);

INVx3_ASAP7_75t_SL g1168 ( 
.A(n_1030),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1074),
.A2(n_1088),
.B(n_1114),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1059),
.B(n_1071),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1000),
.B(n_1054),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1013),
.B(n_1110),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1065),
.B(n_1116),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1009),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1076),
.B(n_1073),
.Y(n_1175)
);

NAND2x1_ASAP7_75t_L g1176 ( 
.A(n_1046),
.B(n_1024),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_992),
.A2(n_1008),
.B1(n_1043),
.B2(n_1026),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1050),
.Y(n_1178)
);

BUFx4_ASAP7_75t_SL g1179 ( 
.A(n_1073),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1032),
.B(n_1016),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1000),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1037),
.B(n_1060),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1063),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1043),
.A2(n_1026),
.B1(n_1016),
.B2(n_982),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1062),
.B(n_1033),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1040),
.B(n_983),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1055),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1035),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1019),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1035),
.B(n_1044),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1004),
.B(n_1022),
.Y(n_1191)
);

CKINVDCx8_ASAP7_75t_R g1192 ( 
.A(n_1062),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1004),
.B(n_1022),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1053),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1087),
.A2(n_1089),
.B(n_989),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1040),
.A2(n_1031),
.B(n_1064),
.C(n_1049),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1048),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1031),
.A2(n_1049),
.B1(n_1006),
.B2(n_1105),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1052),
.B(n_1097),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1022),
.B(n_1006),
.Y(n_1200)
);

NAND3xp33_ASAP7_75t_L g1201 ( 
.A(n_1012),
.B(n_976),
.C(n_1108),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1077),
.A2(n_1102),
.B1(n_1085),
.B2(n_993),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1056),
.B(n_1047),
.Y(n_1203)
);

OAI321xp33_ASAP7_75t_L g1204 ( 
.A1(n_977),
.A2(n_1090),
.A3(n_1084),
.B1(n_1014),
.B2(n_1045),
.C(n_985),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_986),
.A2(n_1021),
.B1(n_1042),
.B2(n_1106),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1041),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_977),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_977),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1084),
.B(n_1090),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1005),
.A2(n_984),
.B(n_1104),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1020),
.B(n_1025),
.Y(n_1211)
);

AOI222xp33_ASAP7_75t_L g1212 ( 
.A1(n_1066),
.A2(n_1079),
.B1(n_1081),
.B2(n_1082),
.C1(n_1101),
.C2(n_1090),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1084),
.A2(n_1100),
.B1(n_1091),
.B2(n_947),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_987),
.B(n_1091),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1034),
.A2(n_1011),
.B(n_1002),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1118),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_994),
.A2(n_955),
.B(n_1002),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1098),
.B(n_988),
.Y(n_1219)
);

AND2x6_ASAP7_75t_L g1220 ( 
.A(n_1023),
.B(n_936),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1057),
.B(n_1058),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1222)
);

INVxp67_ASAP7_75t_L g1223 ( 
.A(n_1007),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1057),
.B(n_1058),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1091),
.A2(n_947),
.B1(n_951),
.B2(n_944),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1061),
.Y(n_1227)
);

NAND2x2_ASAP7_75t_L g1228 ( 
.A(n_1051),
.B(n_640),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1007),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_1069),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1098),
.B(n_988),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1099),
.A2(n_961),
.B(n_955),
.C(n_958),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1233)
);

OAI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1091),
.A2(n_958),
.B(n_1100),
.Y(n_1234)
);

AND2x2_ASAP7_75t_SL g1235 ( 
.A(n_1091),
.B(n_944),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1091),
.A2(n_947),
.B(n_951),
.C(n_944),
.Y(n_1237)
);

BUFx4f_ASAP7_75t_SL g1238 ( 
.A(n_981),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1068),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1061),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_1099),
.B(n_958),
.C(n_955),
.Y(n_1242)
);

BUFx4f_ASAP7_75t_L g1243 ( 
.A(n_981),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1091),
.A2(n_947),
.B(n_951),
.C(n_944),
.Y(n_1244)
);

OAI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1091),
.A2(n_958),
.B(n_1100),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_978),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_978),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1091),
.B(n_1100),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1118),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_978),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1029),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1091),
.A2(n_1100),
.B1(n_947),
.B2(n_951),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1015),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1061),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1091),
.A2(n_958),
.B1(n_944),
.B2(n_951),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_978),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_1162),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1153),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1156),
.Y(n_1259)
);

INVx6_ASAP7_75t_L g1260 ( 
.A(n_1119),
.Y(n_1260)
);

NAND2x1p5_ASAP7_75t_L g1261 ( 
.A(n_1132),
.B(n_1142),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1120),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1121),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1123),
.A2(n_1224),
.B1(n_1244),
.B2(n_1237),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_1253),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1210),
.A2(n_1215),
.B(n_1125),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1197),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_SL g1268 ( 
.A1(n_1252),
.A2(n_1226),
.B1(n_1235),
.B2(n_1141),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1130),
.B(n_1145),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1200),
.B(n_1191),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1251),
.Y(n_1271)
);

CKINVDCx6p67_ASAP7_75t_R g1272 ( 
.A(n_1168),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1251),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1247),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1255),
.A2(n_1252),
.B1(n_1218),
.B2(n_1233),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1256),
.Y(n_1276)
);

NAND2x1p5_ASAP7_75t_L g1277 ( 
.A(n_1132),
.B(n_1142),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1136),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1246),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1250),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1159),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1170),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1152),
.B(n_1242),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1222),
.A2(n_1240),
.B1(n_1248),
.B2(n_1236),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1129),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1242),
.A2(n_1234),
.B1(n_1245),
.B2(n_1217),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1161),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1194),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1147),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1234),
.A2(n_1245),
.B1(n_1217),
.B2(n_1220),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1220),
.A2(n_1177),
.B1(n_1213),
.B2(n_1148),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1157),
.A2(n_1124),
.B1(n_1213),
.B2(n_1149),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1190),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1140),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1220),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1166),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1220),
.A2(n_1149),
.B1(n_1124),
.B2(n_1164),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1185),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1185),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1150),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1137),
.B(n_1214),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1182),
.A2(n_1163),
.B1(n_1131),
.B2(n_1144),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1122),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1216),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1232),
.A2(n_1167),
.B(n_1186),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1203),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1134),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1184),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1127),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1178),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1169),
.A2(n_1195),
.B(n_1128),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1184),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1180),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1146),
.B(n_1173),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1219),
.A2(n_1231),
.B1(n_1138),
.B2(n_1229),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1216),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1193),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1208),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1178),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1187),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1187),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1230),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1181),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1151),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1211),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1126),
.A2(n_1205),
.B(n_1176),
.Y(n_1326)
);

OAI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1157),
.A2(n_1192),
.B1(n_1223),
.B2(n_1181),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1139),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1174),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1174),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1238),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1201),
.A2(n_1209),
.B(n_1171),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1206),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1198),
.A2(n_1189),
.B1(n_1254),
.B2(n_1241),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1198),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1199),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1207),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1227),
.A2(n_1132),
.B1(n_1158),
.B2(n_1239),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1175),
.Y(n_1339)
);

AOI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1204),
.A2(n_1212),
.B(n_1196),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_1243),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1175),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1142),
.B(n_1158),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1135),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_SL g1345 ( 
.A(n_1243),
.B(n_1230),
.Y(n_1345)
);

CKINVDCx6p67_ASAP7_75t_R g1346 ( 
.A(n_1181),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1165),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1165),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1133),
.B(n_1225),
.Y(n_1349)
);

NAND2x1p5_ASAP7_75t_L g1350 ( 
.A(n_1158),
.B(n_1239),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1207),
.Y(n_1351)
);

OAI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1228),
.A2(n_1239),
.B1(n_1183),
.B2(n_1155),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1155),
.A2(n_1133),
.B1(n_1225),
.B2(n_1221),
.Y(n_1353)
);

CKINVDCx6p67_ASAP7_75t_R g1354 ( 
.A(n_1249),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1221),
.A2(n_1155),
.B1(n_1143),
.B2(n_1172),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1249),
.A2(n_1154),
.B1(n_1160),
.B2(n_1143),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1160),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1179),
.A2(n_1204),
.B1(n_1212),
.B2(n_944),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1120),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1120),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1119),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1188),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1197),
.B(n_1176),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1210),
.A2(n_1202),
.B(n_1085),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1153),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1197),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1197),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1197),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1226),
.A2(n_1091),
.B1(n_1100),
.B2(n_958),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1226),
.A2(n_1099),
.B1(n_1080),
.B2(n_1083),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1120),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1210),
.A2(n_1005),
.B(n_1012),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1175),
.B(n_1132),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1140),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1153),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1364),
.A2(n_1326),
.B(n_1372),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1306),
.B(n_1337),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1283),
.B(n_1314),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1283),
.B(n_1314),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1273),
.Y(n_1380)
);

OAI21xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1297),
.A2(n_1290),
.B(n_1286),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1317),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1318),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1336),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1336),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1270),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1270),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1337),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1266),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1273),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1343),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1335),
.Y(n_1392)
);

BUFx4f_ASAP7_75t_SL g1393 ( 
.A(n_1331),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1291),
.B(n_1305),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1301),
.B(n_1284),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1271),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1308),
.B(n_1312),
.Y(n_1397)
);

INVxp33_ASAP7_75t_L g1398 ( 
.A(n_1282),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1332),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1258),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1259),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1343),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1295),
.B(n_1292),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1260),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1375),
.B(n_1295),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1343),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1269),
.B(n_1299),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1296),
.B(n_1293),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1287),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1351),
.B(n_1325),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1275),
.B(n_1315),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1328),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1299),
.B(n_1333),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1264),
.B(n_1370),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1269),
.B(n_1351),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1340),
.A2(n_1310),
.B(n_1320),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1265),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1362),
.Y(n_1419)
);

AOI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1358),
.A2(n_1338),
.B(n_1334),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1319),
.A2(n_1321),
.B(n_1300),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1333),
.B(n_1313),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1278),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1279),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1280),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1268),
.A2(n_1369),
.B1(n_1302),
.B2(n_1327),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1300),
.B(n_1257),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1311),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1298),
.B(n_1289),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1267),
.B(n_1366),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1320),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1261),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1357),
.A2(n_1371),
.B(n_1360),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1320),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1262),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1263),
.B(n_1359),
.Y(n_1436)
);

BUFx4f_ASAP7_75t_SL g1437 ( 
.A(n_1331),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1274),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1363),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1267),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1261),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1276),
.B(n_1347),
.Y(n_1442)
);

AO21x2_ASAP7_75t_L g1443 ( 
.A1(n_1329),
.A2(n_1330),
.B(n_1342),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1373),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1367),
.B(n_1368),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1395),
.B(n_1339),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1417),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1399),
.B(n_1378),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1421),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1394),
.A2(n_1288),
.B1(n_1345),
.B2(n_1341),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1378),
.B(n_1379),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1379),
.B(n_1368),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1439),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_L g1454 ( 
.A(n_1415),
.B(n_1368),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1422),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1421),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1386),
.B(n_1363),
.Y(n_1457)
);

INVxp67_ASAP7_75t_L g1458 ( 
.A(n_1418),
.Y(n_1458)
);

INVx4_ASAP7_75t_SL g1459 ( 
.A(n_1439),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1393),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1433),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1433),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1433),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1437),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1417),
.Y(n_1465)
);

INVxp67_ASAP7_75t_SL g1466 ( 
.A(n_1392),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1387),
.B(n_1344),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1428),
.B(n_1288),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1394),
.A2(n_1348),
.B1(n_1353),
.B2(n_1349),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1431),
.B(n_1355),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1443),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1440),
.Y(n_1472)
);

AO21x2_ASAP7_75t_L g1473 ( 
.A1(n_1389),
.A2(n_1352),
.B(n_1356),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1443),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1392),
.B(n_1346),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1382),
.B(n_1346),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1416),
.B(n_1277),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1416),
.B(n_1350),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1431),
.B(n_1323),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1412),
.B(n_1361),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1434),
.B(n_1408),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1443),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1450),
.A2(n_1426),
.B1(n_1422),
.B2(n_1404),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1480),
.A2(n_1381),
.B1(n_1404),
.B2(n_1441),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1450),
.B(n_1381),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1455),
.B(n_1380),
.Y(n_1486)
);

NAND4xp25_ASAP7_75t_L g1487 ( 
.A(n_1446),
.B(n_1409),
.C(n_1427),
.D(n_1413),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1455),
.B(n_1390),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1451),
.B(n_1396),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1451),
.B(n_1400),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1480),
.B(n_1398),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1469),
.B(n_1384),
.C(n_1385),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1446),
.B(n_1414),
.Y(n_1493)
);

OAI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1469),
.A2(n_1303),
.B1(n_1409),
.B2(n_1401),
.C(n_1403),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1458),
.B(n_1410),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1458),
.B(n_1382),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1468),
.B(n_1423),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1448),
.B(n_1423),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1454),
.B(n_1384),
.C(n_1385),
.Y(n_1499)
);

OAI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1476),
.A2(n_1307),
.B1(n_1407),
.B2(n_1391),
.C(n_1444),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1448),
.B(n_1424),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1447),
.A2(n_1376),
.B(n_1465),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1452),
.B(n_1425),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1475),
.A2(n_1322),
.B1(n_1406),
.B2(n_1420),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1454),
.B(n_1388),
.C(n_1442),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1477),
.B(n_1445),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1454),
.B(n_1430),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1475),
.B(n_1420),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1476),
.A2(n_1438),
.B1(n_1435),
.B2(n_1436),
.C(n_1383),
.Y(n_1509)
);

AOI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1457),
.A2(n_1438),
.B1(n_1435),
.B2(n_1436),
.C(n_1383),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1473),
.A2(n_1397),
.B1(n_1377),
.B2(n_1411),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1473),
.A2(n_1441),
.B1(n_1432),
.B2(n_1402),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1481),
.B(n_1457),
.Y(n_1513)
);

NAND3xp33_ASAP7_75t_L g1514 ( 
.A(n_1471),
.B(n_1388),
.C(n_1411),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1460),
.A2(n_1322),
.B1(n_1405),
.B2(n_1341),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1481),
.B(n_1440),
.Y(n_1516)
);

OAI21xp33_ASAP7_75t_L g1517 ( 
.A1(n_1457),
.A2(n_1397),
.B(n_1429),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1477),
.B(n_1445),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1479),
.B(n_1388),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1467),
.B(n_1419),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1471),
.B(n_1388),
.C(n_1377),
.Y(n_1521)
);

NOR3xp33_ASAP7_75t_SL g1522 ( 
.A(n_1460),
.B(n_1374),
.C(n_1294),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1513),
.B(n_1459),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1502),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1508),
.Y(n_1525)
);

INVxp67_ASAP7_75t_SL g1526 ( 
.A(n_1502),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1508),
.B(n_1466),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1502),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1486),
.B(n_1488),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1513),
.B(n_1447),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1514),
.B(n_1459),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1506),
.B(n_1465),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1518),
.B(n_1465),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1511),
.B(n_1456),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1493),
.B(n_1466),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1474),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1498),
.B(n_1474),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1497),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_1516),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1521),
.B(n_1459),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1485),
.A2(n_1473),
.B1(n_1478),
.B2(n_1470),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1499),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1501),
.B(n_1482),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1496),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1503),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1489),
.B(n_1461),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1512),
.B(n_1449),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1520),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1507),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1507),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1495),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_1510),
.B(n_1472),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1490),
.B(n_1461),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1547),
.B(n_1519),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1538),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_L g1557 ( 
.A(n_1550),
.B(n_1487),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1523),
.B(n_1459),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1462),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1538),
.Y(n_1560)
);

NAND2x1_ASAP7_75t_L g1561 ( 
.A(n_1531),
.B(n_1449),
.Y(n_1561)
);

OAI21xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1553),
.A2(n_1485),
.B(n_1509),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1523),
.B(n_1459),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1525),
.B(n_1542),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1523),
.B(n_1459),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1537),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1525),
.B(n_1462),
.Y(n_1567)
);

INVx2_ASAP7_75t_SL g1568 ( 
.A(n_1523),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1527),
.B(n_1463),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1523),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1463),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1530),
.B(n_1459),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1530),
.B(n_1519),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1554),
.B(n_1517),
.Y(n_1574)
);

NOR4xp25_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1483),
.C(n_1494),
.D(n_1504),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1524),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1524),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1524),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1532),
.B(n_1533),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1550),
.B(n_1551),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1531),
.B(n_1453),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1528),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1481),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1537),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1528),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1537),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1528),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1543),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1568),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1556),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1556),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1560),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1575),
.B(n_1552),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1563),
.B(n_1550),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1557),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1549),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1577),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1564),
.B(n_1536),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1557),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1580),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1560),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1561),
.Y(n_1604)
);

NAND4xp25_ASAP7_75t_L g1605 ( 
.A(n_1564),
.B(n_1580),
.C(n_1484),
.D(n_1571),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1577),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1562),
.A2(n_1553),
.B1(n_1491),
.B2(n_1492),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1566),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1577),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1574),
.B(n_1529),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1575),
.B(n_1552),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1555),
.B(n_1551),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1566),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1565),
.B(n_1549),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1555),
.B(n_1544),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1565),
.B(n_1549),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1578),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1584),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1562),
.A2(n_1553),
.B1(n_1540),
.B2(n_1531),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1558),
.B(n_1531),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_L g1621 ( 
.A(n_1558),
.B(n_1570),
.Y(n_1621)
);

NOR3xp33_ASAP7_75t_L g1622 ( 
.A(n_1571),
.B(n_1500),
.C(n_1515),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1578),
.Y(n_1623)
);

NAND2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1570),
.B(n_1531),
.Y(n_1624)
);

NAND2x1_ASAP7_75t_L g1625 ( 
.A(n_1558),
.B(n_1568),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1574),
.B(n_1554),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1555),
.B(n_1544),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1584),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1583),
.B(n_1535),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1558),
.B(n_1540),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1586),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1608),
.Y(n_1633)
);

AO21x2_ASAP7_75t_L g1634 ( 
.A1(n_1601),
.A2(n_1526),
.B(n_1578),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.B(n_1624),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1596),
.B(n_1568),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1602),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1595),
.B(n_1586),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1624),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1599),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1597),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1621),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1611),
.B(n_1587),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1613),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1618),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1590),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1591),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1629),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1625),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1599),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1607),
.A2(n_1581),
.B1(n_1540),
.B2(n_1547),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1598),
.B(n_1614),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1632),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1598),
.B(n_1581),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_R g1655 ( 
.A(n_1607),
.B(n_1324),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1606),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1592),
.B(n_1587),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1594),
.B(n_1589),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1590),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1610),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1600),
.B(n_1567),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1614),
.B(n_1581),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1606),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1603),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1609),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1609),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1600),
.B(n_1567),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1612),
.Y(n_1668)
);

OAI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1655),
.A2(n_1619),
.B(n_1605),
.C(n_1622),
.Y(n_1669)
);

OAI21xp33_ASAP7_75t_L g1670 ( 
.A1(n_1651),
.A2(n_1626),
.B(n_1615),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1639),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1641),
.A2(n_1522),
.B(n_1526),
.Y(n_1672)
);

AOI322xp5_ASAP7_75t_L g1673 ( 
.A1(n_1641),
.A2(n_1637),
.A3(n_1643),
.B1(n_1638),
.B2(n_1668),
.C1(n_1660),
.C2(n_1647),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1637),
.B(n_1627),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1635),
.A2(n_1631),
.B1(n_1620),
.B2(n_1616),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1635),
.A2(n_1631),
.B1(n_1620),
.B2(n_1616),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1633),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1633),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1644),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1638),
.A2(n_1547),
.B1(n_1626),
.B2(n_1620),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1644),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1660),
.B(n_1324),
.Y(n_1682)
);

AOI32xp33_ASAP7_75t_L g1683 ( 
.A1(n_1643),
.A2(n_1534),
.A3(n_1581),
.B1(n_1589),
.B2(n_1539),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1668),
.B(n_1628),
.Y(n_1684)
);

OAI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1639),
.A2(n_1649),
.B1(n_1642),
.B2(n_1659),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1661),
.B(n_1667),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1642),
.A2(n_1630),
.B(n_1464),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1649),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1636),
.B(n_1572),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1645),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1649),
.A2(n_1540),
.B1(n_1572),
.B2(n_1579),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1573),
.Y(n_1692)
);

CKINVDCx14_ASAP7_75t_R g1693 ( 
.A(n_1636),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1659),
.A2(n_1569),
.B(n_1559),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1671),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1693),
.B(n_1652),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1673),
.B(n_1647),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1689),
.B(n_1642),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1688),
.B(n_1664),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1677),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1682),
.B(n_1464),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1685),
.B(n_1664),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1678),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1674),
.B(n_1646),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1679),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1686),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1675),
.B(n_1642),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1684),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1687),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1672),
.A2(n_1654),
.B1(n_1662),
.B2(n_1667),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1692),
.B(n_1657),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1669),
.B(n_1646),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1676),
.Y(n_1713)
);

NOR2x1_ASAP7_75t_L g1714 ( 
.A(n_1672),
.B(n_1681),
.Y(n_1714)
);

OAI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1714),
.A2(n_1683),
.B(n_1670),
.C(n_1694),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1696),
.B(n_1690),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1696),
.Y(n_1717)
);

AOI211xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1697),
.A2(n_1712),
.B(n_1702),
.C(n_1706),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1695),
.B(n_1680),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1695),
.B(n_1654),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1713),
.A2(n_1680),
.B1(n_1645),
.B2(n_1648),
.C(n_1653),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1707),
.A2(n_1691),
.B(n_1653),
.C(n_1648),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1709),
.A2(n_1662),
.B1(n_1657),
.B2(n_1658),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1708),
.B(n_1707),
.Y(n_1724)
);

NAND4xp75_ASAP7_75t_L g1725 ( 
.A(n_1704),
.B(n_1666),
.C(n_1665),
.D(n_1663),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1698),
.B(n_1661),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1726),
.Y(n_1727)
);

NOR3xp33_ASAP7_75t_L g1728 ( 
.A(n_1724),
.B(n_1699),
.C(n_1701),
.Y(n_1728)
);

INVxp33_ASAP7_75t_L g1729 ( 
.A(n_1717),
.Y(n_1729)
);

NOR3xp33_ASAP7_75t_L g1730 ( 
.A(n_1715),
.B(n_1703),
.C(n_1700),
.Y(n_1730)
);

NAND4xp75_ASAP7_75t_L g1731 ( 
.A(n_1721),
.B(n_1698),
.C(n_1700),
.D(n_1705),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1716),
.Y(n_1732)
);

NOR2x1_ASAP7_75t_L g1733 ( 
.A(n_1725),
.B(n_1705),
.Y(n_1733)
);

XNOR2xp5_ASAP7_75t_L g1734 ( 
.A(n_1720),
.B(n_1710),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1719),
.Y(n_1735)
);

NOR3xp33_ASAP7_75t_L g1736 ( 
.A(n_1723),
.B(n_1711),
.C(n_1374),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1718),
.B(n_1711),
.Y(n_1737)
);

NAND5xp2_ASAP7_75t_L g1738 ( 
.A(n_1728),
.B(n_1718),
.C(n_1722),
.D(n_1666),
.E(n_1665),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1737),
.A2(n_1658),
.B(n_1663),
.C(n_1656),
.Y(n_1739)
);

AOI211xp5_ASAP7_75t_L g1740 ( 
.A1(n_1730),
.A2(n_1663),
.B(n_1656),
.C(n_1650),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1735),
.A2(n_1656),
.B(n_1650),
.C(n_1640),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1727),
.B(n_1294),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1729),
.A2(n_1650),
.B(n_1640),
.C(n_1593),
.Y(n_1743)
);

NAND5xp2_ASAP7_75t_L g1744 ( 
.A(n_1736),
.B(n_1491),
.C(n_1272),
.D(n_1539),
.E(n_1534),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_L g1745 ( 
.A(n_1738),
.B(n_1732),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1739),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1742),
.A2(n_1734),
.B1(n_1733),
.B2(n_1731),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1743),
.B(n_1640),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1740),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1741),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1744),
.A2(n_1634),
.B1(n_1272),
.B2(n_1623),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_L g1752 ( 
.A(n_1749),
.B(n_1634),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1747),
.B(n_1745),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1750),
.Y(n_1754)
);

AOI311xp33_ASAP7_75t_L g1755 ( 
.A1(n_1746),
.A2(n_1634),
.A3(n_1546),
.B(n_1548),
.C(n_1545),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1751),
.B(n_1281),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1753),
.A2(n_1748),
.B1(n_1634),
.B2(n_1623),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1755),
.B(n_1309),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1754),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1759),
.Y(n_1760)
);

OAI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1757),
.B1(n_1758),
.B2(n_1752),
.C(n_1756),
.Y(n_1761)
);

OAI21xp33_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1281),
.B(n_1593),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1761),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1763),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1762),
.B(n_1593),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1765),
.B(n_1309),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1764),
.A2(n_1617),
.B(n_1604),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1617),
.B(n_1585),
.Y(n_1768)
);

AOI322xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1766),
.A3(n_1604),
.B1(n_1576),
.B2(n_1585),
.C1(n_1588),
.C2(n_1582),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_R g1770 ( 
.A1(n_1769),
.A2(n_1309),
.B1(n_1604),
.B2(n_1576),
.C(n_1354),
.Y(n_1770)
);

AOI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1316),
.B(n_1304),
.C(n_1285),
.Y(n_1771)
);


endmodule