module fake_jpeg_27767_n_73 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_15),
.B1(n_26),
.B2(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_36),
.B1(n_32),
.B2(n_13),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_8),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_14),
.B1(n_24),
.B2(n_23),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_42),
.Y(n_44)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_52),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_49),
.B1(n_3),
.B2(n_4),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_6),
.B1(n_44),
.B2(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_12),
.B1(n_22),
.B2(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

A2O1A1O1Ixp25_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_27),
.B(n_20),
.C(n_19),
.D(n_17),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_1),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.C(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.C(n_62),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_4),
.C(n_5),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_5),
.B(n_6),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_56),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_67),
.C(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_62),
.Y(n_70)
);

OAI21x1_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_58),
.B(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_63),
.B(n_46),
.Y(n_72)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_72),
.Y(n_73)
);


endmodule