module fake_jpeg_10369_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_1),
.B(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_44),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_27),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_21),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_63),
.Y(n_69)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_1),
.B(n_2),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_16),
.B1(n_26),
.B2(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_16),
.B1(n_26),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_18),
.B1(n_32),
.B2(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_18),
.B1(n_33),
.B2(n_28),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_29),
.B1(n_28),
.B2(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_23),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_27),
.B(n_19),
.C(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_87),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_48),
.B1(n_62),
.B2(n_3),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_74),
.Y(n_98)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_77),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_0),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_91),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_80),
.Y(n_117)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_86),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_44),
.B1(n_40),
.B2(n_29),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_90),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_8),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_48),
.B1(n_56),
.B2(n_4),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_89),
.B(n_93),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_44),
.B1(n_37),
.B2(n_27),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_0),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_62),
.B(n_0),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_6),
.B(n_7),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_101),
.B1(n_106),
.B2(n_109),
.Y(n_127)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_94),
.B1(n_71),
.B2(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_90),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_62),
.B1(n_48),
.B2(n_56),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_1),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_115),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_10),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_79),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_121),
.C(n_131),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_125),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_70),
.C(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_77),
.C(n_76),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_135),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_66),
.C(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_80),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_117),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_83),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_101),
.C(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_145),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_101),
.B(n_111),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_156),
.B(n_119),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_134),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_109),
.B1(n_115),
.B2(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_129),
.B(n_127),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_125),
.Y(n_169)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_134),
.B1(n_127),
.B2(n_102),
.C(n_124),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_160),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_180),
.B1(n_181),
.B2(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_116),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_166),
.B1(n_164),
.B2(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_169),
.B1(n_164),
.B2(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_123),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_116),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_140),
.C(n_147),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_161),
.C(n_131),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_156),
.B1(n_141),
.B2(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_151),
.B1(n_140),
.B2(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_185),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_168),
.B(n_163),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_186),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_154),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_107),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_188),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_175),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_193),
.B1(n_104),
.B2(n_96),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_174),
.B1(n_176),
.B2(n_172),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_171),
.B(n_180),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_196),
.A2(n_198),
.B(n_190),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_96),
.B1(n_104),
.B2(n_92),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_190),
.B1(n_195),
.B2(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_195),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_201),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_203),
.Y(n_206)
);


endmodule