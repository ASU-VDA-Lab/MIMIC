module fake_jpeg_25011_n_85 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_27),
.B(n_4),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_51),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_13),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_47),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_44),
.B1(n_55),
.B2(n_42),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_63),
.B1(n_57),
.B2(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_58),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_42),
.B1(n_41),
.B2(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_60),
.B(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_66),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_57),
.B1(n_39),
.B2(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_71),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_35),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_72),
.B(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_29),
.Y(n_77)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g80 ( 
.A1(n_77),
.A2(n_16),
.B(n_17),
.C(n_19),
.D(n_22),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_37),
.B1(n_41),
.B2(n_18),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_79),
.A2(n_80),
.B1(n_26),
.B2(n_54),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_79),
.B(n_23),
.Y(n_81)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_81),
.B(n_82),
.CI(n_32),
.CON(n_83),
.SN(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_43),
.Y(n_85)
);


endmodule