module fake_jpeg_17327_n_25 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_25;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_3),
.Y(n_8)
);

AOI22xp33_ASAP7_75t_SL g9 ( 
.A1(n_4),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_4),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_8),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_16),
.C(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_0),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_9),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_13),
.B(n_10),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_11),
.B1(n_8),
.B2(n_13),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_23),
.C(n_17),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

AOI322xp5_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_15),
.A3(n_20),
.B1(n_14),
.B2(n_10),
.C1(n_16),
.C2(n_11),
.Y(n_25)
);


endmodule