module fake_jpeg_31145_n_512 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_512);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_512;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_84),
.Y(n_106)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_8),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_54),
.B(n_63),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_66),
.Y(n_164)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_8),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_99),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_50),
.B(n_6),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_23),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_156),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_50),
.B1(n_25),
.B2(n_26),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_123),
.A2(n_149),
.B1(n_66),
.B2(n_64),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_37),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_142),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_78),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_65),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_79),
.A2(n_50),
.B1(n_26),
.B2(n_18),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_149),
.B1(n_85),
.B2(n_91),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_51),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

AO22x2_ASAP7_75t_L g149 ( 
.A1(n_93),
.A2(n_101),
.B1(n_98),
.B2(n_96),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_76),
.B(n_51),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_69),
.B(n_37),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_72),
.A2(n_24),
.B(n_39),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_73),
.B(n_20),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_23),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_165),
.A2(n_181),
.B1(n_193),
.B2(n_196),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_182),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_106),
.A2(n_27),
.B(n_33),
.C(n_29),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_168),
.B(n_171),
.Y(n_240)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_33),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_109),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_172),
.B(n_173),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_26),
.B1(n_92),
.B2(n_81),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_177),
.A2(n_190),
.B1(n_203),
.B2(n_205),
.Y(n_221)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_105),
.A2(n_90),
.B1(n_89),
.B2(n_77),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_140),
.B(n_0),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_18),
.C(n_24),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_42),
.B1(n_29),
.B2(n_20),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_75),
.B1(n_70),
.B2(n_55),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_120),
.A2(n_19),
.B1(n_47),
.B2(n_42),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_147),
.Y(n_228)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_131),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_207),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_202),
.B1(n_137),
.B2(n_134),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_149),
.A2(n_61),
.B1(n_27),
.B2(n_47),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_144),
.A2(n_17),
.B1(n_40),
.B2(n_19),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_141),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_204),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_135),
.A2(n_40),
.B1(n_68),
.B2(n_39),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_206),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_142),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_151),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVxp67_ASAP7_75t_R g211 ( 
.A(n_129),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_211),
.B(n_13),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_161),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_213),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_108),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_39),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_214),
.Y(n_219)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_215),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_195),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_187),
.A2(n_112),
.B1(n_122),
.B2(n_132),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_230),
.A2(n_248),
.B1(n_199),
.B2(n_183),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_231),
.A2(n_165),
.B1(n_123),
.B2(n_196),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_228),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_238),
.B(n_251),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_169),
.A2(n_107),
.B1(n_148),
.B2(n_139),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_104),
.C(n_162),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_209),
.C(n_188),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_174),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_167),
.B(n_68),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_255),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_174),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_271),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_257),
.Y(n_294)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_259),
.A2(n_277),
.B1(n_289),
.B2(n_170),
.Y(n_293)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_262),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_182),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_209),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_269),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_167),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_270),
.B(n_273),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_211),
.C(n_188),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_236),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_274),
.Y(n_305)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_176),
.C(n_198),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_288),
.Y(n_292)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_276),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_231),
.A2(n_134),
.B1(n_119),
.B2(n_138),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_168),
.B(n_204),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_220),
.B(n_237),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_219),
.B(n_179),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_282),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_180),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_234),
.A2(n_221),
.B1(n_254),
.B2(n_238),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_224),
.B(n_218),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_283),
.A2(n_222),
.B1(n_242),
.B2(n_236),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_234),
.A2(n_226),
.B1(n_247),
.B2(n_178),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_287),
.B1(n_237),
.B2(n_220),
.Y(n_295)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_285),
.B(n_286),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_229),
.B(n_189),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_233),
.A2(n_175),
.B1(n_185),
.B2(n_197),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_233),
.A2(n_164),
.B1(n_138),
.B2(n_145),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_246),
.Y(n_290)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_290),
.A2(n_24),
.B(n_250),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_293),
.A2(n_301),
.B1(n_257),
.B2(n_265),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_295),
.A2(n_319),
.B1(n_263),
.B2(n_273),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_296),
.B(n_280),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_281),
.A2(n_164),
.B1(n_160),
.B2(n_191),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_298),
.A2(n_300),
.B1(n_310),
.B2(n_313),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_245),
.B1(n_192),
.B2(n_184),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_272),
.A2(n_222),
.B1(n_183),
.B2(n_242),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_303),
.A2(n_289),
.B1(n_258),
.B2(n_276),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_267),
.A2(n_220),
.B(n_237),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_304),
.A2(n_307),
.B(n_321),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_241),
.B(n_206),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_269),
.A2(n_235),
.B1(n_241),
.B2(n_194),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_259),
.A2(n_235),
.B1(n_217),
.B2(n_239),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_215),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_318),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_227),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_277),
.A2(n_110),
.B1(n_239),
.B2(n_227),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_274),
.A2(n_186),
.B(n_225),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_322),
.Y(n_366)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_323),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_299),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_324),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_325),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_282),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_326),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_279),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_327),
.B(n_328),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_309),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_264),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_329),
.B(n_336),
.Y(n_358)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_330),
.Y(n_355)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_274),
.B(n_280),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_335),
.A2(n_337),
.B(n_338),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_310),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_260),
.B(n_261),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_275),
.Y(n_339)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_340),
.A2(n_341),
.B1(n_301),
.B2(n_296),
.Y(n_359)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_308),
.Y(n_342)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_343),
.A2(n_348),
.B1(n_313),
.B2(n_298),
.Y(n_361)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_344),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_306),
.B(n_271),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_345),
.B(n_346),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_270),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_256),
.B1(n_285),
.B2(n_287),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_352),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_305),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_350),
.Y(n_378)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_292),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_369),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_359),
.A2(n_352),
.B1(n_325),
.B2(n_328),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_315),
.C(n_292),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_363),
.C(n_364),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_361),
.A2(n_380),
.B1(n_381),
.B2(n_347),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_307),
.B1(n_291),
.B2(n_295),
.Y(n_362)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_315),
.C(n_314),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_304),
.C(n_305),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_305),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_331),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_305),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_300),
.C(n_319),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_370),
.B(n_347),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_294),
.C(n_229),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_322),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_348),
.A2(n_294),
.B1(n_317),
.B2(n_312),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_317),
.B1(n_312),
.B2(n_257),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_377),
.B(n_327),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_384),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_402),
.Y(n_431)
);

A2O1A1Ixp33_ASAP7_75t_SL g386 ( 
.A1(n_356),
.A2(n_349),
.B(n_338),
.C(n_343),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_386),
.A2(n_411),
.B(n_244),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_381),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_387),
.B(n_390),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_383),
.B(n_326),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_398),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_391),
.A2(n_404),
.B1(n_389),
.B2(n_406),
.Y(n_430)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_393),
.A2(n_400),
.B1(n_380),
.B2(n_370),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_401),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_342),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_396),
.Y(n_428)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_397),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_375),
.B(n_346),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_324),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_399),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_368),
.A2(n_323),
.B1(n_340),
.B2(n_349),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_356),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_336),
.Y(n_402)
);

A2O1A1O1Ixp25_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_329),
.B(n_349),
.C(n_330),
.D(n_333),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_SL g414 ( 
.A1(n_403),
.A2(n_409),
.B(n_410),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_361),
.A2(n_341),
.B1(n_340),
.B2(n_351),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_344),
.Y(n_406)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_407),
.B(n_408),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_379),
.A2(n_317),
.B(n_322),
.Y(n_408)
);

OAI32xp33_ASAP7_75t_L g410 ( 
.A1(n_378),
.A2(n_225),
.A3(n_250),
.B1(n_244),
.B2(n_110),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_379),
.A2(n_364),
.B(n_368),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_433),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_387),
.A2(n_371),
.B1(n_353),
.B2(n_374),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_419),
.A2(n_420),
.B1(n_425),
.B2(n_432),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_393),
.A2(n_374),
.B1(n_355),
.B2(n_365),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_360),
.C(n_354),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_422),
.C(n_429),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_373),
.C(n_369),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_400),
.A2(n_365),
.B1(n_382),
.B2(n_366),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_405),
.C(n_409),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_430),
.A2(n_28),
.B1(n_22),
.B2(n_39),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_408),
.A2(n_382),
.B1(n_367),
.B2(n_217),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_426),
.Y(n_436)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_428),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_437),
.B(n_438),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_416),
.B(n_390),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_405),
.C(n_385),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_441),
.C(n_447),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_406),
.C(n_391),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_403),
.B1(n_404),
.B2(n_386),
.Y(n_444)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_423),
.B(n_252),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_446),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_423),
.B(n_410),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_386),
.C(n_104),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_448),
.A2(n_424),
.B1(n_415),
.B2(n_412),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_386),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_451),
.C(n_424),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_450),
.A2(n_432),
.B1(n_420),
.B2(n_425),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_118),
.C(n_39),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_452),
.A2(n_457),
.B1(n_459),
.B2(n_466),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_414),
.B1(n_413),
.B2(n_427),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_427),
.B1(n_430),
.B2(n_415),
.Y(n_459)
);

XOR2x1_ASAP7_75t_SL g460 ( 
.A(n_449),
.B(n_433),
.Y(n_460)
);

MAJx2_ASAP7_75t_L g470 ( 
.A(n_460),
.B(n_9),
.C(n_15),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_9),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_32),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_447),
.A2(n_412),
.B1(n_10),
.B2(n_4),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_6),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_28),
.C(n_22),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_468),
.C(n_32),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_450),
.B1(n_441),
.B2(n_451),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_22),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_467),
.A2(n_435),
.B(n_439),
.Y(n_469)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_32),
.C(n_28),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_472),
.B(n_477),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_474),
.Y(n_485)
);

BUFx24_ASAP7_75t_SL g474 ( 
.A(n_454),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_460),
.A2(n_9),
.B(n_15),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_475),
.A2(n_480),
.B(n_5),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_478),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_32),
.C(n_6),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_481),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_453),
.A2(n_6),
.B(n_12),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_32),
.C(n_4),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_482),
.B(n_465),
.C(n_458),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_483),
.B(n_1),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_SL g487 ( 
.A1(n_475),
.A2(n_452),
.B(n_459),
.C(n_457),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_487),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_466),
.B1(n_463),
.B2(n_464),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_490),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_462),
.B1(n_5),
.B2(n_10),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_10),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_476),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_495),
.A2(n_499),
.B(n_500),
.Y(n_502)
);

AOI21xp33_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_487),
.B(n_2),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_484),
.A2(n_470),
.B(n_10),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_498),
.A2(n_487),
.B(n_483),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_12),
.Y(n_499)
);

A2O1A1O1Ixp25_ASAP7_75t_L g501 ( 
.A1(n_497),
.A2(n_486),
.B(n_489),
.C(n_487),
.D(n_493),
.Y(n_501)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_503),
.A2(n_504),
.B(n_494),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_502),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_507),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_506),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_495),
.B(n_1),
.Y(n_510)
);

NAND3xp33_ASAP7_75t_L g511 ( 
.A(n_510),
.B(n_1),
.C(n_2),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_511),
.A2(n_2),
.B(n_505),
.Y(n_512)
);


endmodule