module real_aes_2960_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_0), .B(n_136), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_1), .A2(n_144), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_2), .B(n_777), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_3), .A2(n_105), .B1(n_773), .B2(n_780), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_4), .B(n_136), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_5), .B(n_163), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_6), .B(n_163), .Y(n_485) );
INVx1_ASAP7_75t_L g132 ( .A(n_7), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_8), .B(n_163), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g777 ( .A(n_9), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g762 ( .A1(n_10), .A2(n_14), .B1(n_763), .B2(n_764), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_10), .Y(n_763) );
NAND2xp33_ASAP7_75t_L g526 ( .A(n_11), .B(n_161), .Y(n_526) );
AND2x2_ASAP7_75t_L g166 ( .A(n_12), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g177 ( .A(n_13), .B(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_14), .Y(n_764) );
INVx2_ASAP7_75t_L g123 ( .A(n_15), .Y(n_123) );
AOI221x1_ASAP7_75t_L g470 ( .A1(n_16), .A2(n_29), .B1(n_136), .B2(n_144), .C(n_471), .Y(n_470) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_17), .A2(n_22), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_17), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_18), .B(n_163), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_19), .Y(n_110) );
NOR3xp33_ASAP7_75t_L g775 ( .A(n_19), .B(n_776), .C(n_778), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_20), .B(n_136), .Y(n_522) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_21), .A2(n_178), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_22), .B(n_121), .Y(n_474) );
INVxp67_ASAP7_75t_L g768 ( .A(n_22), .Y(n_768) );
AOI22xp5_ASAP7_75t_SL g732 ( .A1(n_23), .A2(n_733), .B1(n_734), .B2(n_740), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_23), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_24), .B(n_163), .Y(n_459) );
AO21x1_ASAP7_75t_L g480 ( .A1(n_25), .A2(n_136), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_26), .B(n_136), .Y(n_219) );
INVx1_ASAP7_75t_L g744 ( .A(n_27), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_28), .A2(n_92), .B1(n_127), .B2(n_136), .Y(n_126) );
NAND2x1_ASAP7_75t_L g501 ( .A(n_30), .B(n_163), .Y(n_501) );
NAND2x1_ASAP7_75t_L g533 ( .A(n_31), .B(n_161), .Y(n_533) );
OR2x2_ASAP7_75t_L g124 ( .A(n_32), .B(n_89), .Y(n_124) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_32), .A2(n_89), .B(n_123), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_33), .B(n_161), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_34), .B(n_163), .Y(n_525) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_35), .A2(n_167), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_36), .B(n_161), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_37), .A2(n_144), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_38), .B(n_163), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_39), .A2(n_144), .B(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g134 ( .A(n_40), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g142 ( .A(n_40), .B(n_132), .Y(n_142) );
INVx1_ASAP7_75t_L g148 ( .A(n_40), .Y(n_148) );
OR2x6_ASAP7_75t_L g742 ( .A(n_41), .B(n_743), .Y(n_742) );
INVxp67_ASAP7_75t_L g778 ( .A(n_41), .Y(n_778) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_42), .B(n_136), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_43), .B(n_136), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_44), .B(n_163), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_45), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_46), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_47), .B(n_161), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_48), .B(n_136), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_49), .A2(n_144), .B(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_50), .A2(n_735), .B1(n_736), .B2(n_739), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_50), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_51), .A2(n_144), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_52), .B(n_161), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_53), .B(n_161), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_54), .B(n_136), .Y(n_200) );
INVx1_ASAP7_75t_L g130 ( .A(n_55), .Y(n_130) );
INVx1_ASAP7_75t_L g139 ( .A(n_55), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_56), .B(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g209 ( .A(n_57), .B(n_121), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_58), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_59), .B(n_163), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_60), .B(n_161), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_61), .A2(n_144), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_62), .B(n_136), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_63), .B(n_136), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_64), .A2(n_144), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g225 ( .A(n_65), .B(n_122), .Y(n_225) );
AO21x1_ASAP7_75t_L g482 ( .A1(n_66), .A2(n_144), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_67), .B(n_136), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_68), .B(n_161), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_69), .B(n_136), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_70), .B(n_161), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_71), .A2(n_96), .B1(n_144), .B2(n_146), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_72), .B(n_163), .Y(n_222) );
AND2x2_ASAP7_75t_L g495 ( .A(n_73), .B(n_122), .Y(n_495) );
INVx1_ASAP7_75t_L g135 ( .A(n_74), .Y(n_135) );
INVx1_ASAP7_75t_L g141 ( .A(n_74), .Y(n_141) );
AND2x2_ASAP7_75t_L g536 ( .A(n_75), .B(n_167), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_76), .B(n_161), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_77), .A2(n_144), .B(n_213), .Y(n_212) );
AOI22xp5_ASAP7_75t_SL g736 ( .A1(n_78), .A2(n_83), .B1(n_737), .B2(n_738), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_78), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_79), .A2(n_144), .B(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_80), .A2(n_144), .B(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g235 ( .A(n_81), .B(n_122), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_82), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g737 ( .A(n_83), .Y(n_737) );
INVx1_ASAP7_75t_L g745 ( .A(n_84), .Y(n_745) );
AND2x2_ASAP7_75t_L g447 ( .A(n_85), .B(n_167), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_86), .B(n_136), .Y(n_461) );
AND2x2_ASAP7_75t_L g190 ( .A(n_87), .B(n_178), .Y(n_190) );
AND2x2_ASAP7_75t_L g481 ( .A(n_88), .B(n_205), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_90), .B(n_161), .Y(n_460) );
AND2x2_ASAP7_75t_L g504 ( .A(n_91), .B(n_167), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_93), .B(n_163), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_94), .A2(n_144), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_95), .B(n_161), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_97), .A2(n_144), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_98), .B(n_163), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_99), .B(n_163), .Y(n_452) );
BUFx2_ASAP7_75t_L g224 ( .A(n_100), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_101), .Y(n_749) );
BUFx2_ASAP7_75t_L g754 ( .A(n_102), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_103), .A2(n_144), .B(n_524), .Y(n_523) );
AO221x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_750), .B1(n_755), .B2(n_758), .C(n_770), .Y(n_105) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_741), .B1(n_746), .B2(n_749), .Y(n_106) );
XOR2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_732), .Y(n_107) );
OAI22xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_110), .B1(n_111), .B2(n_440), .Y(n_108) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g748 ( .A(n_110), .B(n_742), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_110), .B(n_741), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_111), .A2(n_761), .B1(n_762), .B2(n_765), .Y(n_760) );
INVx3_ASAP7_75t_L g761 ( .A(n_111), .Y(n_761) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_365), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_301), .C(n_348), .Y(n_112) );
NAND4xp25_ASAP7_75t_SL g113 ( .A(n_114), .B(n_236), .C(n_254), .D(n_280), .Y(n_113) );
OAI21xp33_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_194), .B(n_195), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_116), .B(n_179), .Y(n_115) );
INVx1_ASAP7_75t_L g416 ( .A(n_116), .Y(n_416) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_151), .Y(n_116) );
INVx2_ASAP7_75t_L g240 ( .A(n_117), .Y(n_240) );
AND2x2_ASAP7_75t_L g260 ( .A(n_117), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g362 ( .A(n_117), .B(n_181), .Y(n_362) );
AND2x2_ASAP7_75t_L g422 ( .A(n_117), .B(n_241), .Y(n_422) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_118), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g306 ( .A(n_119), .B(n_154), .Y(n_306) );
BUFx3_ASAP7_75t_L g316 ( .A(n_119), .Y(n_316) );
AND2x2_ASAP7_75t_L g379 ( .A(n_119), .B(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_125), .Y(n_119) );
AND2x4_ASAP7_75t_L g193 ( .A(n_120), .B(n_125), .Y(n_193) );
AO21x2_ASAP7_75t_L g125 ( .A1(n_121), .A2(n_126), .B(n_143), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_121), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_121), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_121), .A2(n_449), .B(n_450), .Y(n_448) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_121), .A2(n_470), .B(n_474), .Y(n_469) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_121), .A2(n_470), .B(n_474), .Y(n_540) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_SL g122 ( .A(n_123), .B(n_124), .Y(n_122) );
AND2x4_ASAP7_75t_L g205 ( .A(n_123), .B(n_124), .Y(n_205) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_133), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g145 ( .A(n_130), .B(n_132), .Y(n_145) );
AND2x4_ASAP7_75t_L g163 ( .A(n_130), .B(n_140), .Y(n_163) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x6_ASAP7_75t_L g144 ( .A(n_134), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g150 ( .A(n_135), .Y(n_150) );
AND2x6_ASAP7_75t_L g161 ( .A(n_135), .B(n_138), .Y(n_161) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_142), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx5_ASAP7_75t_L g164 ( .A(n_142), .Y(n_164) );
AND2x4_ASAP7_75t_L g146 ( .A(n_145), .B(n_147), .Y(n_146) );
NOR2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g425 ( .A(n_152), .Y(n_425) );
AND2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_168), .Y(n_152) );
AND2x2_ASAP7_75t_L g192 ( .A(n_153), .B(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g380 ( .A(n_153), .Y(n_380) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g194 ( .A(n_154), .B(n_183), .Y(n_194) );
AND2x2_ASAP7_75t_L g257 ( .A(n_154), .B(n_168), .Y(n_257) );
INVx2_ASAP7_75t_L g262 ( .A(n_154), .Y(n_262) );
AND2x2_ASAP7_75t_L g264 ( .A(n_154), .B(n_169), .Y(n_264) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_166), .Y(n_154) );
INVx4_ASAP7_75t_L g167 ( .A(n_155), .Y(n_167) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx4f_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_165), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_164), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_161), .B(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_164), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_164), .A2(n_188), .B(n_189), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_164), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_164), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_164), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_164), .A2(n_452), .B(n_453), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_164), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_164), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_164), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_164), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_164), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_164), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_164), .A2(n_533), .B(n_534), .Y(n_532) );
INVx3_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
INVx1_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
INVx2_ASAP7_75t_L g246 ( .A(n_168), .Y(n_246) );
AND2x4_ASAP7_75t_SL g277 ( .A(n_168), .B(n_183), .Y(n_277) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_168), .Y(n_309) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_169), .Y(n_191) );
AOI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_177), .Y(n_169) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_170), .A2(n_530), .B(n_536), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_176), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_178), .A2(n_219), .B(n_220), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_192), .Y(n_179) );
AND2x2_ASAP7_75t_L g343 ( .A(n_180), .B(n_288), .Y(n_343) );
INVx2_ASAP7_75t_SL g431 ( .A(n_180), .Y(n_431) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_191), .Y(n_181) );
NAND2x1p5_ASAP7_75t_L g244 ( .A(n_182), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g351 ( .A(n_182), .B(n_264), .Y(n_351) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx2_ASAP7_75t_L g239 ( .A(n_183), .Y(n_239) );
AND2x4_ASAP7_75t_L g241 ( .A(n_183), .B(n_242), .Y(n_241) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_183), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g334 ( .A(n_183), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_183), .B(n_292), .Y(n_353) );
AND2x2_ASAP7_75t_L g384 ( .A(n_183), .B(n_293), .Y(n_384) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_190), .Y(n_183) );
AND2x2_ASAP7_75t_L g323 ( .A(n_192), .B(n_277), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_192), .B(n_334), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_192), .A2(n_434), .B1(n_436), .B2(n_437), .Y(n_433) );
AND2x2_ASAP7_75t_L g436 ( .A(n_192), .B(n_243), .Y(n_436) );
INVx3_ASAP7_75t_L g289 ( .A(n_193), .Y(n_289) );
AND2x2_ASAP7_75t_L g292 ( .A(n_193), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g308 ( .A(n_194), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g317 ( .A(n_194), .Y(n_317) );
AND2x4_ASAP7_75t_SL g195 ( .A(n_196), .B(n_206), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_196), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g368 ( .A(n_196), .B(n_369), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g420 ( .A(n_196), .B(n_330), .C(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g438 ( .A(n_196), .B(n_332), .Y(n_438) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g253 ( .A(n_198), .B(n_217), .Y(n_253) );
INVx1_ASAP7_75t_L g270 ( .A(n_198), .Y(n_270) );
INVx2_ASAP7_75t_L g283 ( .A(n_198), .Y(n_283) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_198), .Y(n_298) );
AND2x2_ASAP7_75t_L g312 ( .A(n_198), .B(n_285), .Y(n_312) );
AND2x2_ASAP7_75t_L g391 ( .A(n_198), .B(n_208), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_205), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_205), .A2(n_211), .B(n_212), .Y(n_210) );
INVx1_ASAP7_75t_SL g455 ( .A(n_205), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_205), .B(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_205), .A2(n_522), .B(n_523), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g254 ( .A1(n_206), .A2(n_255), .B1(n_258), .B2(n_265), .C(n_271), .Y(n_254) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_206), .A2(n_384), .B1(n_385), .B2(n_386), .C(n_387), .Y(n_383) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
INVx2_ASAP7_75t_L g325 ( .A(n_207), .Y(n_325) );
AND2x2_ASAP7_75t_L g385 ( .A(n_207), .B(n_269), .Y(n_385) );
AND2x2_ASAP7_75t_L g395 ( .A(n_207), .B(n_281), .Y(n_395) );
OR2x2_ASAP7_75t_L g435 ( .A(n_207), .B(n_319), .Y(n_435) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_SL g252 ( .A(n_208), .B(n_253), .Y(n_252) );
NAND2x1_ASAP7_75t_L g268 ( .A(n_208), .B(n_217), .Y(n_268) );
INVx4_ASAP7_75t_L g297 ( .A(n_208), .Y(n_297) );
OR2x2_ASAP7_75t_L g339 ( .A(n_208), .B(n_226), .Y(n_339) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
AND2x2_ASAP7_75t_L g390 ( .A(n_216), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_226), .Y(n_216) );
INVx2_ASAP7_75t_SL g278 ( .A(n_217), .Y(n_278) );
NOR2x1_ASAP7_75t_SL g284 ( .A(n_217), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g299 ( .A(n_217), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g330 ( .A(n_217), .B(n_297), .Y(n_330) );
AND2x2_ASAP7_75t_L g337 ( .A(n_217), .B(n_283), .Y(n_337) );
BUFx2_ASAP7_75t_L g371 ( .A(n_217), .Y(n_371) );
AND2x2_ASAP7_75t_L g382 ( .A(n_217), .B(n_297), .Y(n_382) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_225), .Y(n_217) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_226), .Y(n_250) );
AND2x2_ASAP7_75t_L g269 ( .A(n_226), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g300 ( .A(n_226), .Y(n_300) );
AND2x2_ASAP7_75t_L g326 ( .A(n_226), .B(n_282), .Y(n_326) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_227) );
AO21x1_ASAP7_75t_SL g285 ( .A1(n_228), .A2(n_229), .B(n_235), .Y(n_285) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_228), .A2(n_489), .B(n_495), .Y(n_488) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_228), .A2(n_498), .B(n_504), .Y(n_497) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_228), .A2(n_498), .B(n_504), .Y(n_510) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_228), .A2(n_489), .B(n_495), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_234), .Y(n_229) );
OAI31xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_241), .A3(n_243), .B(n_247), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g345 ( .A(n_239), .Y(n_345) );
NOR2xp67_ASAP7_75t_L g255 ( .A(n_240), .B(n_256), .Y(n_255) );
AOI322xp5_ASAP7_75t_L g335 ( .A1(n_240), .A2(n_329), .A3(n_336), .B1(n_340), .B2(n_341), .C1(n_343), .C2(n_344), .Y(n_335) );
AND2x2_ASAP7_75t_L g407 ( .A(n_240), .B(n_384), .Y(n_407) );
AOI221xp5_ASAP7_75t_SL g320 ( .A1(n_241), .A2(n_321), .B1(n_323), .B2(n_324), .C(n_327), .Y(n_320) );
INVx2_ASAP7_75t_L g340 ( .A(n_241), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_243), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_243), .B(n_336), .Y(n_439) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g314 ( .A(n_244), .B(n_289), .Y(n_314) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g293 ( .A(n_246), .B(n_262), .Y(n_293) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g364 ( .A(n_250), .Y(n_364) );
O2A1O1Ixp5_ASAP7_75t_L g355 ( .A1(n_251), .A2(n_356), .B(n_358), .C(n_360), .Y(n_355) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_252), .A2(n_388), .B1(n_389), .B2(n_392), .Y(n_387) );
OR2x2_ASAP7_75t_L g342 ( .A(n_253), .B(n_339), .Y(n_342) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_259), .B(n_263), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_264), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g318 ( .A(n_268), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_268), .B(n_269), .Y(n_361) );
OR2x2_ASAP7_75t_L g363 ( .A(n_268), .B(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_268), .B(n_412), .Y(n_411) );
BUFx2_ASAP7_75t_L g279 ( .A(n_270), .Y(n_279) );
NOR4xp25_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .C(n_278), .D(n_279), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g399 ( .A(n_273), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g427 ( .A(n_273), .B(n_276), .Y(n_427) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g357 ( .A(n_275), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_276), .B(n_305), .Y(n_392) );
AOI321xp33_ASAP7_75t_L g394 ( .A1(n_276), .A2(n_395), .A3(n_396), .B1(n_397), .B2(n_399), .C(n_402), .Y(n_394) );
INVx2_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_277), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_277), .B(n_316), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_278), .B(n_300), .Y(n_405) );
OR2x2_ASAP7_75t_L g432 ( .A(n_279), .B(n_316), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_286), .B(n_290), .Y(n_280) );
AND2x2_ASAP7_75t_L g321 ( .A(n_281), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g347 ( .A(n_283), .B(n_285), .Y(n_347) );
INVx2_ASAP7_75t_L g332 ( .A(n_284), .Y(n_332) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_287), .B(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g388 ( .A(n_288), .B(n_340), .Y(n_388) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g346 ( .A(n_289), .B(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_289), .B(n_425), .Y(n_424) );
NOR2xp67_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g375 ( .A(n_293), .Y(n_375) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_297), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
BUFx2_ASAP7_75t_L g404 ( .A(n_297), .Y(n_404) );
INVxp67_ASAP7_75t_L g412 ( .A(n_300), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_320), .C(n_335), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_310), .B(n_313), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g333 ( .A(n_306), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g386 ( .A(n_307), .Y(n_386) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g401 ( .A(n_309), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_310), .A2(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g319 ( .A(n_312), .Y(n_319) );
AND2x2_ASAP7_75t_L g381 ( .A(n_312), .B(n_382), .Y(n_381) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_318), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_314), .A2(n_361), .B1(n_362), .B2(n_363), .Y(n_360) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g350 ( .A(n_316), .Y(n_350) );
OR2x2_ASAP7_75t_L g398 ( .A(n_319), .B(n_330), .Y(n_398) );
NOR4xp25_ASAP7_75t_L g430 ( .A(n_322), .B(n_371), .C(n_431), .D(n_432), .Y(n_430) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
OR2x2_ASAP7_75t_L g331 ( .A(n_325), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_325), .B(n_347), .Y(n_429) );
AOI21xp33_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_331), .B(n_333), .Y(n_327) );
INVx2_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g418 ( .A(n_330), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g426 ( .A(n_332), .Y(n_426) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVxp67_ASAP7_75t_L g354 ( .A(n_337), .Y(n_354) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g370 ( .A(n_339), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AND2x2_ASAP7_75t_L g373 ( .A(n_345), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g419 ( .A(n_347), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B(n_354), .C(n_355), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g409 ( .A(n_351), .Y(n_409) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g413 ( .A(n_356), .Y(n_413) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR3xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_393), .C(n_414), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_372), .B(n_376), .C(n_383), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_379), .B(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g415 ( .A1(n_379), .A2(n_416), .B(n_417), .C(n_420), .Y(n_415) );
BUFx2_ASAP7_75t_L g396 ( .A(n_380), .Y(n_396) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_406), .Y(n_393) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_403), .A2(n_409), .B1(n_410), .B2(n_413), .Y(n_408) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_415), .B(n_423), .C(n_433), .D(n_439), .Y(n_414) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_427), .B2(n_428), .C(n_430), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_619), .Y(n_440) );
AO211x2_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_464), .B(n_514), .C(n_587), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
AND3x2_ASAP7_75t_L g668 ( .A(n_444), .B(n_549), .C(n_565), .Y(n_668) );
AND2x4_ASAP7_75t_L g671 ( .A(n_444), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_445), .B(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g580 ( .A(n_445), .Y(n_580) );
AND2x2_ASAP7_75t_SL g665 ( .A(n_445), .B(n_574), .Y(n_665) );
AND2x2_ASAP7_75t_L g708 ( .A(n_445), .B(n_529), .Y(n_708) );
INVx5_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g557 ( .A(n_446), .Y(n_557) );
AND2x2_ASAP7_75t_L g576 ( .A(n_446), .B(n_520), .Y(n_576) );
AND2x2_ASAP7_75t_L g594 ( .A(n_446), .B(n_529), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_446), .B(n_528), .Y(n_654) );
NOR2x1_ASAP7_75t_SL g681 ( .A(n_446), .B(n_454), .Y(n_681) );
OR2x6_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_454), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B(n_462), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_455), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_455), .A2(n_456), .B(n_462), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
AO21x1_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_496), .B(n_505), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_466), .A2(n_563), .B1(n_567), .B2(n_568), .Y(n_562) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
AND2x2_ASAP7_75t_L g623 ( .A(n_467), .B(n_511), .Y(n_623) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g556 ( .A(n_468), .B(n_539), .Y(n_556) );
AND2x2_ASAP7_75t_L g628 ( .A(n_468), .B(n_513), .Y(n_628) );
AND2x2_ASAP7_75t_L g647 ( .A(n_468), .B(n_613), .Y(n_647) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g506 ( .A(n_469), .Y(n_506) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_469), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_475), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g607 ( .A(n_476), .B(n_508), .Y(n_607) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_488), .Y(n_476) );
AND2x2_ASAP7_75t_L g511 ( .A(n_477), .B(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g544 ( .A(n_477), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_477), .B(n_540), .Y(n_604) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g697 ( .A(n_478), .Y(n_697) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g539 ( .A(n_479), .Y(n_539) );
OAI21x1_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_482), .B(n_486), .Y(n_479) );
INVx1_ASAP7_75t_L g487 ( .A(n_481), .Y(n_487) );
INVx2_ASAP7_75t_L g545 ( .A(n_488), .Y(n_545) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_488), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_490), .B(n_494), .Y(n_489) );
INVx2_ASAP7_75t_L g541 ( .A(n_496), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_496), .B(n_673), .Y(n_699) );
AND2x2_ASAP7_75t_L g718 ( .A(n_496), .B(n_708), .Y(n_718) );
BUFx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_SL g586 ( .A(n_497), .B(n_545), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_506), .B(n_507), .Y(n_505) );
AND2x2_ASAP7_75t_L g585 ( .A(n_506), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_506), .B(n_555), .Y(n_590) );
INVx1_ASAP7_75t_SL g717 ( .A(n_506), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_507), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g543 ( .A(n_508), .Y(n_543) );
AND2x2_ASAP7_75t_L g729 ( .A(n_508), .B(n_730), .Y(n_729) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g605 ( .A(n_509), .B(n_512), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_509), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g659 ( .A(n_509), .B(n_513), .Y(n_659) );
AND2x2_ASAP7_75t_L g690 ( .A(n_509), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g555 ( .A(n_510), .B(n_513), .Y(n_555) );
INVxp67_ASAP7_75t_L g572 ( .A(n_510), .Y(n_572) );
BUFx3_ASAP7_75t_L g613 ( .A(n_510), .Y(n_613) );
AND2x2_ASAP7_75t_L g633 ( .A(n_511), .B(n_634), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g646 ( .A(n_511), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_512), .B(n_539), .Y(n_602) );
AND2x2_ASAP7_75t_L g691 ( .A(n_512), .B(n_540), .Y(n_691) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g618 ( .A(n_513), .B(n_540), .Y(n_618) );
OR3x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_562), .C(n_577), .Y(n_514) );
OAI321xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_527), .A3(n_537), .B1(n_542), .B2(n_546), .C(n_554), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_519), .Y(n_593) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_519), .Y(n_611) );
OR2x2_ASAP7_75t_L g615 ( .A(n_519), .B(n_527), .Y(n_615) );
BUFx3_ASAP7_75t_L g549 ( .A(n_520), .Y(n_549) );
AND2x2_ASAP7_75t_L g566 ( .A(n_520), .B(n_552), .Y(n_566) );
INVx1_ASAP7_75t_L g583 ( .A(n_520), .Y(n_583) );
INVx2_ASAP7_75t_L g599 ( .A(n_520), .Y(n_599) );
OR2x2_ASAP7_75t_L g638 ( .A(n_520), .B(n_528), .Y(n_638) );
INVx2_ASAP7_75t_L g626 ( .A(n_527), .Y(n_626) );
AND2x2_ASAP7_75t_L g550 ( .A(n_528), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g565 ( .A(n_528), .Y(n_565) );
AND2x4_ASAP7_75t_L g574 ( .A(n_528), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_528), .B(n_551), .Y(n_597) );
AND2x2_ASAP7_75t_L g704 ( .A(n_528), .B(n_599), .Y(n_704) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_529), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
INVx1_ASAP7_75t_L g591 ( .A(n_537), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_538), .B(n_541), .Y(n_537) );
AND2x2_ASAP7_75t_L g678 ( .A(n_538), .B(n_605), .Y(n_678) );
INVx1_ASAP7_75t_SL g695 ( .A(n_538), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_538), .B(n_671), .Y(n_724) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OR2x2_ASAP7_75t_L g567 ( .A(n_539), .B(n_540), .Y(n_567) );
AND2x2_ASAP7_75t_L g660 ( .A(n_541), .B(n_556), .Y(n_660) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_545), .B(n_556), .Y(n_683) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_547), .A2(n_696), .B1(n_701), .B2(n_703), .Y(n_700) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g625 ( .A(n_548), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g720 ( .A(n_548), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g676 ( .A(n_549), .B(n_594), .Y(n_676) );
AND2x4_ASAP7_75t_L g630 ( .A(n_550), .B(n_576), .Y(n_630) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_552), .Y(n_728) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g561 ( .A(n_553), .Y(n_561) );
INVx1_ASAP7_75t_L g575 ( .A(n_553), .Y(n_575) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_557), .D(n_558), .Y(n_554) );
AND2x2_ASAP7_75t_L g712 ( .A(n_555), .B(n_697), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_555), .B(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_556), .B(n_632), .Y(n_631) );
OAI322xp33_ASAP7_75t_L g639 ( .A1(n_556), .A2(n_640), .A3(n_644), .B1(n_646), .B2(n_648), .C1(n_650), .C2(n_655), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_556), .B(n_605), .Y(n_655) );
INVx1_ASAP7_75t_L g723 ( .A(n_556), .Y(n_723) );
INVx2_ASAP7_75t_L g569 ( .A(n_557), .Y(n_569) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_560), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_561), .B(n_580), .Y(n_637) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_564), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g610 ( .A(n_565), .Y(n_610) );
AND2x2_ASAP7_75t_L g682 ( .A(n_565), .B(n_593), .Y(n_682) );
AOI31xp33_ASAP7_75t_L g568 ( .A1(n_566), .A2(n_569), .A3(n_570), .B(n_573), .Y(n_568) );
AND2x2_ASAP7_75t_L g579 ( .A(n_566), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g707 ( .A(n_566), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_SL g714 ( .A(n_566), .B(n_594), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_566), .Y(n_715) );
INVx1_ASAP7_75t_SL g673 ( .A(n_567), .Y(n_673) );
NAND3xp33_ASAP7_75t_SL g701 ( .A(n_567), .B(n_695), .C(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g601 ( .A(n_572), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
AND2x2_ASAP7_75t_L g582 ( .A(n_574), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g643 ( .A(n_574), .Y(n_643) );
AOI322xp5_ASAP7_75t_L g725 ( .A1(n_574), .A2(n_604), .A3(n_607), .B1(n_726), .B2(n_727), .C1(n_729), .C2(n_731), .Y(n_725) );
AND2x2_ASAP7_75t_L g731 ( .A(n_574), .B(n_580), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_584), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_580), .B(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g726 ( .A(n_580), .B(n_613), .Y(n_726) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g652 ( .A(n_583), .Y(n_652) );
AND2x2_ASAP7_75t_L g680 ( .A(n_583), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g727 ( .A(n_583), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g632 ( .A(n_586), .Y(n_632) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
O2A1O1Ixp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B(n_592), .C(n_595), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g649 ( .A(n_594), .B(n_599), .Y(n_649) );
OAI211xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_600), .B(n_606), .C(n_608), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_596), .A2(n_622), .B1(n_624), .B2(n_627), .C(n_629), .Y(n_621) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g641 ( .A(n_598), .Y(n_641) );
OR2x2_ASAP7_75t_L g661 ( .A(n_598), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g706 ( .A(n_601), .Y(n_706) );
INVx1_ASAP7_75t_L g730 ( .A(n_602), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g612 ( .A(n_604), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_604), .B(n_674), .Y(n_686) );
INVx1_ASAP7_75t_L g666 ( .A(n_605), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B1(n_614), .B2(n_616), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_SL g674 ( .A(n_613), .Y(n_674) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND4xp75_ASAP7_75t_L g619 ( .A(n_620), .B(n_656), .C(n_684), .D(n_709), .Y(n_619) );
NOR2xp67_ASAP7_75t_L g620 ( .A(n_621), .B(n_639), .Y(n_620) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_628), .B(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_633), .B2(n_635), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_632), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx2_ASAP7_75t_L g672 ( .A(n_638), .Y(n_672) );
OR2x2_ASAP7_75t_L g687 ( .A(n_638), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g702 ( .A(n_647), .Y(n_702) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_649), .A2(n_694), .B(n_696), .Y(n_693) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_669), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B1(n_664), .B2(n_666), .C(n_667), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g705 ( .A1(n_659), .A2(n_706), .B(n_707), .Y(n_705) );
INVx3_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
OAI322xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_673), .A3(n_674), .B1(n_675), .B2(n_677), .C1(n_679), .C2(n_683), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g692 ( .A(n_680), .Y(n_692) );
INVx1_ASAP7_75t_L g688 ( .A(n_681), .Y(n_688) );
AND2x2_ASAP7_75t_L g703 ( .A(n_681), .B(n_704), .Y(n_703) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_685), .B(n_698), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_689), .B2(n_692), .C(n_693), .Y(n_685) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_692), .A2(n_699), .B(n_700), .C(n_705), .Y(n_698) );
INVx2_ASAP7_75t_SL g721 ( .A(n_708), .Y(n_721) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_710), .B(n_719), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .B1(n_715), .B2(n_716), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
OAI211xp5_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_722), .B(n_724), .C(n_725), .Y(n_719) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx12_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
CKINVDCx5p33_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_744), .B(n_745), .Y(n_779) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR2x1_ASAP7_75t_R g755 ( .A(n_754), .B(n_756), .Y(n_755) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g772 ( .A(n_757), .Y(n_772) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_759), .A2(n_760), .B1(n_766), .B2(n_767), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g765 ( .A(n_762), .Y(n_765) );
INVxp33_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_773), .Y(n_780) );
CKINVDCx6p67_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g774 ( .A(n_775), .B(n_779), .Y(n_774) );
endmodule