module real_jpeg_25657_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_34),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_1),
.A2(n_43),
.B1(n_58),
.B2(n_60),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_1),
.A2(n_22),
.B1(n_28),
.B2(n_43),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_1),
.A2(n_43),
.B1(n_56),
.B2(n_131),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_2),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_2),
.A2(n_58),
.B1(n_60),
.B2(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_2),
.A2(n_34),
.B1(n_37),
.B2(n_106),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_2),
.A2(n_22),
.B1(n_28),
.B2(n_106),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_4),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_4),
.A2(n_29),
.B1(n_56),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_29),
.B1(n_34),
.B2(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_29),
.B1(n_58),
.B2(n_60),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_54),
.B(n_107),
.C(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_4),
.B(n_57),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_60),
.B(n_78),
.C(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_22),
.C(n_36),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_4),
.B(n_76),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_4),
.B(n_11),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_4),
.B(n_38),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_7),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_40),
.B1(n_58),
.B2(n_60),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_7),
.A2(n_22),
.B1(n_28),
.B2(n_40),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_11),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_135),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_133),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_108),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_15),
.B(n_108),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_85),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_65),
.B2(n_66),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_20),
.A2(n_30),
.B1(n_45),
.B2(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_20),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_20),
.A2(n_45),
.B1(n_191),
.B2(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B(n_27),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_21),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_21),
.B(n_27),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_21),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_22),
.B(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_26),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_29),
.A2(n_53),
.B(n_60),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_29),
.A2(n_37),
.B(n_79),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_30),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_39),
.B(n_41),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_31),
.A2(n_69),
.B(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_32),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_32),
.B(n_70),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_32),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_34),
.A2(n_37),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_34),
.B(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_38),
.B(n_196),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_39),
.A2(n_71),
.B(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_41),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_41),
.B(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_61),
.B(n_62),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_49),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_49),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_49),
.B(n_63),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_57),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_57),
.B(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_57),
.B(n_130),
.Y(n_161)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_60),
.B1(n_78),
.B2(n_79),
.Y(n_82)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_74),
.B(n_84),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_68),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_73),
.B(n_206),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_80),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_76),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_83),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_77),
.A2(n_81),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_77),
.B(n_126),
.Y(n_159)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_80),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_81),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_94),
.C(n_100),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_87),
.B(n_93),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_88),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_91),
.A2(n_118),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_91),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_100),
.B1(n_101),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_95),
.B(n_157),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_97),
.B(n_150),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_114),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_109),
.B(n_112),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_114),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_125),
.C(n_127),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_115),
.A2(n_116),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_123),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_120),
.B(n_219),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_124),
.B(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_125),
.A2(n_127),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_125),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_127),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_273),
.B(n_277),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_184),
.B(n_259),
.C(n_272),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_172),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_138),
.B(n_172),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_154),
.B2(n_171),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_152),
.B2(n_153),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_141),
.B(n_153),
.C(n_171),
.Y(n_260)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_148),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_144),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_151),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_156),
.B(n_163),
.C(n_164),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.C(n_179),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_173),
.A2(n_174),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_179),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.C(n_182),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_182),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_258),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_200),
.B(n_257),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_187),
.B(n_197),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_193),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_190),
.B(n_193),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_191),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_252),
.B(n_256),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_243),
.B(n_251),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_223),
.B(n_242),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_230),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_217),
.B2(n_222),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_213),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_216),
.C(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_231),
.B(n_241),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_225),
.B(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_237),
.B(n_240),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_248),
.C(n_249),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_271),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_269),
.B2(n_270),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_270),
.C(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);


endmodule