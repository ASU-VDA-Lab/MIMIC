module fake_jpeg_297_n_704 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_704);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_704;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_60),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_61),
.Y(n_187)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_64),
.B(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_69),
.Y(n_171)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_76),
.Y(n_183)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_80),
.A2(n_57),
.B1(n_55),
.B2(n_31),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_81),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_82),
.Y(n_203)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_83),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_84),
.Y(n_227)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_19),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_104),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_91),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_93),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_95),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_101),
.Y(n_221)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_21),
.B(n_19),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_43),
.B(n_18),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_18),
.Y(n_182)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_54),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_59),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_44),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_115),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_22),
.Y(n_120)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_22),
.Y(n_121)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_24),
.Y(n_125)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_28),
.Y(n_126)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_24),
.Y(n_127)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_25),
.Y(n_128)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_25),
.Y(n_129)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_25),
.Y(n_130)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_25),
.Y(n_131)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_132),
.A2(n_59),
.B(n_27),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_79),
.B1(n_92),
.B2(n_93),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_136),
.A2(n_138),
.B1(n_152),
.B2(n_204),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_83),
.A2(n_26),
.B1(n_21),
.B2(n_50),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_71),
.B(n_26),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_139),
.B(n_182),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_145),
.A2(n_157),
.B1(n_158),
.B2(n_173),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_50),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_147),
.B(n_167),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_58),
.B1(n_39),
.B2(n_49),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_20),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_154),
.A2(n_197),
.B(n_95),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_57),
.B1(n_55),
.B2(n_31),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_61),
.A2(n_58),
.B1(n_39),
.B2(n_49),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_73),
.B(n_58),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_72),
.A2(n_49),
.B1(n_39),
.B2(n_55),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_105),
.B(n_28),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_176),
.B(n_192),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_185),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_105),
.B(n_28),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_76),
.B(n_20),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_196),
.B(n_10),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_82),
.A2(n_20),
.B1(n_57),
.B2(n_31),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_199),
.A2(n_223),
.B1(n_9),
.B2(n_10),
.Y(n_292)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_80),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_121),
.Y(n_209)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_62),
.A2(n_40),
.B1(n_33),
.B2(n_67),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_210),
.A2(n_214),
.B1(n_219),
.B2(n_0),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_130),
.A2(n_94),
.B1(n_91),
.B2(n_84),
.Y(n_214)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_108),
.B(n_33),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_16),
.C(n_15),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_120),
.B(n_40),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_225),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_96),
.A2(n_59),
.B1(n_37),
.B2(n_42),
.Y(n_219)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_129),
.A2(n_36),
.B1(n_42),
.B2(n_41),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_114),
.B(n_32),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_116),
.A2(n_36),
.B1(n_42),
.B2(n_41),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_229),
.A2(n_36),
.B(n_35),
.Y(n_245)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_119),
.Y(n_230)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_230),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_232),
.B(n_304),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_37),
.B1(n_32),
.B2(n_35),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_235),
.A2(n_255),
.B1(n_277),
.B2(n_282),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_134),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_236),
.B(n_307),
.Y(n_319)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_148),
.Y(n_237)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_237),
.Y(n_336)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_37),
.B1(n_32),
.B2(n_35),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_241),
.A2(n_245),
.B1(n_259),
.B2(n_287),
.Y(n_322)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_242),
.Y(n_366)
);

BUFx8_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

INVx11_ASAP7_75t_L g346 ( 
.A(n_243),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_246),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_247),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_154),
.A2(n_27),
.B1(n_132),
.B2(n_52),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_248),
.A2(n_257),
.B1(n_263),
.B2(n_264),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_249),
.B(n_261),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_250),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_159),
.B(n_27),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_251),
.B(n_276),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_144),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_252),
.Y(n_330)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_253),
.Y(n_368)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_136),
.A2(n_75),
.B1(n_99),
.B2(n_52),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_184),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_185),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_259)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_162),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_227),
.Y(n_262)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_180),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_264)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_181),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_265),
.Y(n_339)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_177),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_266),
.B(n_269),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_180),
.A2(n_13),
.B1(n_11),
.B2(n_2),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_270),
.A2(n_274),
.B1(n_288),
.B2(n_290),
.Y(n_341)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_156),
.Y(n_271)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_271),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_231),
.Y(n_272)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_146),
.B(n_0),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_273),
.B(n_175),
.C(n_164),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_207),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_206),
.Y(n_275)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_275),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_150),
.B(n_0),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_157),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_143),
.A2(n_1),
.B(n_5),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_279),
.A2(n_302),
.B(n_289),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_179),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_160),
.B(n_5),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_283),
.B(n_285),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_223),
.B(n_6),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_213),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_286)
);

OA22x2_ASAP7_75t_L g379 ( 
.A1(n_286),
.A2(n_292),
.B1(n_260),
.B2(n_253),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_191),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_207),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_141),
.B(n_9),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g372 ( 
.A(n_289),
.B(n_252),
.Y(n_372)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_181),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_156),
.Y(n_291)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_291),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_140),
.Y(n_293)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_155),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_296),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_295),
.B(n_305),
.Y(n_343)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_161),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_186),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_297),
.B(n_298),
.Y(n_373)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_165),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_174),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_299),
.B(n_301),
.Y(n_375)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_212),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_137),
.A2(n_10),
.B(n_142),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_153),
.A2(n_171),
.B1(n_221),
.B2(n_135),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_303),
.A2(n_306),
.B1(n_309),
.B2(n_311),
.Y(n_360)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_170),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_153),
.B(n_171),
.Y(n_305)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_181),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_140),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

INVx11_ASAP7_75t_L g309 ( 
.A(n_144),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_172),
.B(n_195),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_211),
.Y(n_340)
);

INVx11_ASAP7_75t_L g311 ( 
.A(n_178),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_215),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_186),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_208),
.B(n_194),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_314),
.B(n_178),
.Y(n_348)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_215),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_315),
.B(n_316),
.Y(n_344)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_202),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_300),
.A2(n_198),
.B(n_149),
.C(n_169),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_321),
.B(n_332),
.Y(n_391)
);

NOR2x1_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_193),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_325),
.A2(n_355),
.B(n_237),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_281),
.A2(n_226),
.B1(n_211),
.B2(n_166),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_331),
.A2(n_246),
.B1(n_256),
.B2(n_272),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_251),
.A2(n_208),
.B(n_183),
.C(n_163),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_234),
.A2(n_183),
.B1(n_163),
.B2(n_228),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_333),
.A2(n_374),
.B(n_249),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_340),
.B(n_352),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_258),
.B(n_133),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_353),
.C(n_243),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_358),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g352 ( 
.A(n_280),
.B(n_168),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_239),
.B(n_238),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_302),
.A2(n_228),
.B(n_189),
.C(n_206),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_354),
.B(n_315),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_281),
.B(n_151),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_297),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_277),
.A2(n_205),
.B1(n_226),
.B2(n_189),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_359),
.A2(n_311),
.B1(n_316),
.B2(n_268),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_241),
.A2(n_205),
.B1(n_175),
.B2(n_166),
.Y(n_361)
);

OAI21xp33_ASAP7_75t_SL g386 ( 
.A1(n_361),
.A2(n_365),
.B(n_379),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_276),
.B(n_164),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_364),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_363),
.B(n_372),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_283),
.B(n_273),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_255),
.A2(n_220),
.B1(n_291),
.B2(n_271),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_273),
.B(n_220),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_310),
.B(n_289),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_243),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_330),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_279),
.B(n_245),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_284),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_355),
.A2(n_292),
.B1(n_308),
.B2(n_293),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_380),
.A2(n_383),
.B1(n_390),
.B2(n_403),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_385),
.C(n_401),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_355),
.A2(n_262),
.B1(n_235),
.B2(n_240),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_375),
.Y(n_384)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_318),
.B(n_244),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_375),
.Y(n_387)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_387),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_334),
.A2(n_247),
.B1(n_267),
.B2(n_250),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

INVx3_ASAP7_75t_SL g393 ( 
.A(n_349),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_337),
.A2(n_309),
.B1(n_242),
.B2(n_290),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_394),
.A2(n_411),
.B1(n_417),
.B2(n_420),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_357),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_402),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_378),
.A2(n_254),
.B(n_278),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_396),
.A2(n_415),
.B(n_341),
.Y(n_460)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_398),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_406),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_294),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_320),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_334),
.A2(n_304),
.B1(n_301),
.B2(n_299),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_298),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_419),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_410),
.B1(n_421),
.B2(n_422),
.Y(n_438)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_409),
.B(n_412),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_331),
.A2(n_233),
.B1(n_307),
.B2(n_268),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_414),
.Y(n_452)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_354),
.A2(n_374),
.B(n_332),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_328),
.B(n_296),
.C(n_278),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_401),
.C(n_372),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_337),
.A2(n_233),
.B1(n_284),
.B2(n_312),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_418),
.B(n_348),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_318),
.B(n_275),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_328),
.A2(n_265),
.B1(n_306),
.B2(n_362),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_333),
.A2(n_322),
.B1(n_370),
.B2(n_363),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_322),
.A2(n_364),
.B1(n_328),
.B2(n_317),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_373),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_429),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_371),
.B(n_340),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_425),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_326),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_325),
.A2(n_379),
.B1(n_327),
.B2(n_319),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_426),
.A2(n_376),
.B1(n_342),
.B2(n_336),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_326),
.B(n_343),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_428),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_373),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_344),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_425),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_433),
.B(n_457),
.Y(n_488)
);

AO22x1_ASAP7_75t_SL g437 ( 
.A1(n_380),
.A2(n_325),
.B1(n_379),
.B2(n_352),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_437),
.B(n_441),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_395),
.B(n_372),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_451),
.C(n_455),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_385),
.B(n_372),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_447),
.B(n_448),
.Y(n_479)
);

AO22x2_ASAP7_75t_L g450 ( 
.A1(n_383),
.A2(n_379),
.B1(n_321),
.B2(n_345),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_450),
.B(n_458),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_323),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_422),
.B1(n_400),
.B2(n_406),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_454),
.A2(n_456),
.B1(n_459),
.B2(n_461),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_407),
.B(n_376),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_386),
.A2(n_327),
.B1(n_329),
.B2(n_366),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_398),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_366),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_415),
.A2(n_329),
.B1(n_351),
.B2(n_338),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_460),
.A2(n_396),
.B(n_418),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_424),
.B(n_342),
.Y(n_462)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_462),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_391),
.A2(n_360),
.B(n_377),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_463),
.A2(n_392),
.B(n_391),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_381),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_464),
.B(n_470),
.Y(n_508)
);

FAx1_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_330),
.CI(n_339),
.CON(n_466),
.SN(n_466)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_466),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_336),
.Y(n_467)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_467),
.A2(n_420),
.B(n_381),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_407),
.B(n_369),
.C(n_339),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_411),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_419),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_458),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_472),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_467),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_511),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_475),
.A2(n_478),
.B(n_496),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_451),
.B(n_382),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_476),
.B(n_437),
.Y(n_546)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_430),
.Y(n_480)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_480),
.Y(n_516)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_481),
.Y(n_521)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_482),
.Y(n_538)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_486),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_453),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_510),
.Y(n_528)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_440),
.Y(n_489)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_489),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_432),
.B(n_388),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_500),
.C(n_505),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_438),
.A2(n_399),
.B1(n_417),
.B2(n_384),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_493),
.A2(n_499),
.B1(n_501),
.B2(n_506),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_494),
.B(n_442),
.Y(n_529)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_495),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_445),
.A2(n_466),
.B(n_465),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_445),
.A2(n_397),
.B(n_387),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_497),
.A2(n_503),
.B(n_504),
.Y(n_515)
);

OAI32xp33_ASAP7_75t_L g498 ( 
.A1(n_435),
.A2(n_466),
.A3(n_445),
.B1(n_439),
.B2(n_462),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_498),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_438),
.A2(n_390),
.B1(n_388),
.B2(n_405),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_404),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_434),
.A2(n_405),
.B1(n_428),
.B2(n_408),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_471),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_502),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_445),
.A2(n_427),
.B(n_416),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_460),
.A2(n_389),
.B(n_403),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_434),
.A2(n_389),
.B1(n_393),
.B2(n_413),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_466),
.A2(n_369),
.B(n_412),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_507),
.A2(n_496),
.B(n_491),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_470),
.A2(n_393),
.B1(n_413),
.B2(n_412),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_509),
.A2(n_449),
.B1(n_469),
.B2(n_444),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_453),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_444),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_451),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_512),
.B(n_518),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_473),
.B(n_443),
.C(n_468),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_517),
.B(n_525),
.C(n_526),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_455),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_508),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_519),
.B(n_495),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_508),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_520),
.B(n_532),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_488),
.A2(n_464),
.B1(n_433),
.B2(n_457),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_522),
.A2(n_533),
.B(n_536),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_497),
.B(n_455),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_492),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_435),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_500),
.B(n_441),
.C(n_447),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_L g563 ( 
.A1(n_529),
.A2(n_479),
.B(n_502),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_488),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_509),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_534),
.B(n_537),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_535),
.A2(n_539),
.B1(n_543),
.B2(n_545),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_485),
.A2(n_442),
.B1(n_461),
.B2(n_439),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_472),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_485),
.A2(n_454),
.B1(n_449),
.B2(n_463),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_504),
.A2(n_456),
.B1(n_437),
.B2(n_448),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_475),
.A2(n_459),
.B(n_431),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_544),
.A2(n_507),
.B(n_478),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_491),
.A2(n_437),
.B1(n_450),
.B2(n_431),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_546),
.B(n_479),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_503),
.B(n_450),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_550),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_452),
.C(n_446),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_524),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_551),
.B(n_555),
.Y(n_599)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_552),
.Y(n_603)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_541),
.Y(n_553)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_541),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g600 ( 
.A(n_556),
.B(n_565),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_527),
.A2(n_480),
.B1(n_481),
.B2(n_474),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_558),
.A2(n_559),
.B1(n_563),
.B2(n_578),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_527),
.A2(n_513),
.B1(n_539),
.B2(n_549),
.Y(n_559)
);

XNOR2x1_ASAP7_75t_L g589 ( 
.A(n_560),
.B(n_582),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_516),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_561),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_531),
.A2(n_498),
.B(n_492),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_566),
.A2(n_567),
.B(n_570),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_531),
.A2(n_477),
.B(n_484),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_530),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_568),
.B(n_576),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_482),
.Y(n_569)
);

CKINVDCx14_ASAP7_75t_R g611 ( 
.A(n_569),
.Y(n_611)
);

AO32x1_ASAP7_75t_L g570 ( 
.A1(n_515),
.A2(n_477),
.A3(n_493),
.B1(n_450),
.B2(n_501),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_515),
.A2(n_484),
.B(n_499),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_533),
.A2(n_544),
.B(n_543),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_572),
.A2(n_547),
.B(n_542),
.Y(n_605)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_516),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_579),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_525),
.B(n_350),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_528),
.B(n_483),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_514),
.B(n_519),
.Y(n_580)
);

AOI21xp33_ASAP7_75t_SL g596 ( 
.A1(n_580),
.A2(n_489),
.B(n_511),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_514),
.B(n_486),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_518),
.Y(n_586)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_521),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_583),
.A2(n_584),
.B1(n_548),
.B2(n_547),
.Y(n_592)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_538),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_586),
.B(n_596),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_517),
.C(n_526),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_587),
.B(n_590),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_562),
.B(n_512),
.C(n_523),
.Y(n_590)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_592),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_581),
.B(n_557),
.C(n_573),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_593),
.B(n_594),
.C(n_607),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_557),
.B(n_546),
.C(n_522),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_558),
.A2(n_513),
.B1(n_536),
.B2(n_545),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_595),
.A2(n_567),
.B1(n_560),
.B2(n_572),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_554),
.A2(n_535),
.B1(n_506),
.B2(n_542),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_601),
.A2(n_570),
.B1(n_583),
.B2(n_576),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_SL g602 ( 
.A(n_556),
.B(n_548),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_602),
.B(n_604),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_SL g604 ( 
.A(n_573),
.B(n_566),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_605),
.B(n_610),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_574),
.B(n_540),
.C(n_538),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_540),
.C(n_452),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_608),
.B(n_577),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_571),
.B(n_446),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_598),
.A2(n_552),
.B1(n_551),
.B2(n_568),
.Y(n_612)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_612),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_609),
.B(n_577),
.Y(n_614)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_614),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_615),
.B(n_616),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_611),
.B(n_579),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_618),
.A2(n_619),
.B1(n_624),
.B2(n_627),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_598),
.A2(n_559),
.B1(n_570),
.B2(n_575),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_591),
.A2(n_564),
.B(n_582),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_620),
.A2(n_591),
.B(n_589),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_606),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_621),
.B(n_631),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_595),
.B(n_555),
.Y(n_622)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_622),
.Y(n_645)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_609),
.Y(n_625)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_625),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_601),
.A2(n_553),
.B1(n_561),
.B2(n_584),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_606),
.Y(n_628)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_628),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_603),
.A2(n_561),
.B1(n_450),
.B2(n_414),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_629),
.A2(n_630),
.B1(n_633),
.B2(n_597),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_588),
.A2(n_450),
.B1(n_402),
.B2(n_338),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_592),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_605),
.A2(n_409),
.B1(n_350),
.B2(n_335),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_620),
.B(n_586),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g660 ( 
.A(n_636),
.B(n_639),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_626),
.B(n_587),
.C(n_593),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_637),
.B(n_642),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_619),
.B(n_604),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_641),
.B(n_638),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_626),
.B(n_607),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_SL g643 ( 
.A(n_617),
.B(n_594),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_SL g656 ( 
.A(n_643),
.B(n_617),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_646),
.A2(n_649),
.B1(n_653),
.B2(n_625),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_614),
.B(n_597),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_613),
.B(n_608),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_651),
.B(n_621),
.Y(n_662)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_613),
.B(n_590),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_652),
.B(n_632),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_628),
.Y(n_653)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_655),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g679 ( 
.A(n_656),
.B(n_658),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_637),
.B(n_634),
.C(n_631),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_657),
.B(n_659),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_SL g658 ( 
.A(n_639),
.B(n_632),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_644),
.B(n_585),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_661),
.B(n_662),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_663),
.A2(n_665),
.B(n_667),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_645),
.A2(n_627),
.B1(n_624),
.B2(n_623),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_664),
.B(n_668),
.C(n_610),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_SL g665 ( 
.A1(n_635),
.A2(n_623),
.B1(n_599),
.B2(n_633),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_651),
.B(n_599),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_666),
.B(n_648),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_650),
.A2(n_618),
.B1(n_589),
.B2(n_630),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_636),
.B(n_646),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_638),
.B(n_652),
.C(n_643),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_669),
.B(n_640),
.C(n_647),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_671),
.B(n_677),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_654),
.A2(n_647),
.B(n_649),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_673),
.A2(n_680),
.B(n_668),
.Y(n_685)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_674),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_657),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_678),
.B(n_658),
.Y(n_686)
);

OAI221xp5_ASAP7_75t_L g680 ( 
.A1(n_656),
.A2(n_641),
.B1(n_629),
.B2(n_602),
.C(n_600),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g681 ( 
.A(n_655),
.B(n_600),
.C(n_351),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g689 ( 
.A(n_681),
.B(n_356),
.C(n_367),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_676),
.B(n_669),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_682),
.B(n_683),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_676),
.B(n_660),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_685),
.A2(n_675),
.B(n_672),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_686),
.B(n_687),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_SL g687 ( 
.A1(n_670),
.A2(n_409),
.B1(n_349),
.B2(n_356),
.Y(n_687)
);

AOI31xp33_ASAP7_75t_L g694 ( 
.A1(n_689),
.A2(n_681),
.A3(n_679),
.B(n_678),
.Y(n_694)
);

AOI21x1_ASAP7_75t_L g697 ( 
.A1(n_690),
.A2(n_694),
.B(n_346),
.Y(n_697)
);

OAI21xp33_ASAP7_75t_L g692 ( 
.A1(n_684),
.A2(n_688),
.B(n_671),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_692),
.A2(n_679),
.B(n_689),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_695),
.A2(n_696),
.B(n_697),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_SL g696 ( 
.A1(n_691),
.A2(n_687),
.B(n_324),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_696),
.B(n_693),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_699),
.Y(n_700)
);

MAJIxp5_ASAP7_75t_L g701 ( 
.A(n_700),
.B(n_698),
.C(n_356),
.Y(n_701)
);

MAJIxp5_ASAP7_75t_L g702 ( 
.A(n_701),
.B(n_367),
.C(n_346),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_702),
.B(n_367),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_SL g704 ( 
.A1(n_703),
.A2(n_324),
.B(n_335),
.Y(n_704)
);


endmodule