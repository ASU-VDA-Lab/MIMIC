module fake_jpeg_22230_n_303 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_46),
.B(n_26),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_30),
.B1(n_31),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_47),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_25),
.B(n_23),
.C(n_18),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_40),
.B(n_8),
.C(n_9),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_54),
.Y(n_82)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_24),
.C(n_34),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_18),
.C(n_20),
.Y(n_92)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_59),
.B1(n_29),
.B2(n_18),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_17),
.B1(n_31),
.B2(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_32),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_75),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_25),
.B(n_36),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_92),
.C(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_19),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_79),
.B1(n_97),
.B2(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_81),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_21),
.B1(n_28),
.B2(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_26),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_96),
.B1(n_100),
.B2(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_98),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_45),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_54),
.B(n_29),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_20),
.B1(n_42),
.B2(n_40),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_20),
.B1(n_42),
.B2(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_61),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_12),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_106),
.A2(n_129),
.B1(n_69),
.B2(n_103),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_109),
.B1(n_126),
.B2(n_76),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_92),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_67),
.B1(n_50),
.B2(n_51),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_124),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_78),
.A2(n_57),
.A3(n_8),
.B1(n_10),
.B2(n_16),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_1),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_130),
.A2(n_98),
.B(n_85),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_142),
.C(n_69),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_154),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_135),
.A2(n_162),
.B(n_1),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_73),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_143),
.B(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_124),
.B1(n_123),
.B2(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_146),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_86),
.B(n_89),
.C(n_91),
.D(n_84),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_153),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_83),
.B(n_74),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_151),
.B1(n_15),
.B2(n_13),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_106),
.A2(n_111),
.B1(n_104),
.B2(n_119),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_94),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_159),
.B(n_160),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_80),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_113),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_74),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_156),
.B(n_158),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_87),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g160 ( 
.A1(n_107),
.A2(n_129),
.B1(n_127),
.B2(n_105),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_93),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_130),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_115),
.B(n_128),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_172),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_170),
.A2(n_174),
.B(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_69),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_176),
.B1(n_187),
.B2(n_192),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_70),
.C(n_121),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_177),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_93),
.B1(n_95),
.B2(n_99),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_178),
.B(n_181),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_121),
.Y(n_179)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_116),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_189),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_93),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_57),
.C(n_90),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_90),
.Y(n_186)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_1),
.Y(n_188)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_191),
.B1(n_141),
.B2(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_149),
.B1(n_146),
.B2(n_163),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_191),
.A2(n_149),
.B1(n_160),
.B2(n_162),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_201),
.B1(n_192),
.B2(n_181),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_206),
.B1(n_215),
.B2(n_5),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_137),
.B(n_148),
.C(n_142),
.D(n_143),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_174),
.C(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_153),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_166),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_186),
.A2(n_147),
.B1(n_137),
.B2(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_167),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_136),
.B(n_151),
.Y(n_206)
);

XOR2x2_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_143),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_R g239 ( 
.A(n_207),
.B(n_4),
.Y(n_239)
);

OAI322xp33_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_159),
.A3(n_155),
.B1(n_150),
.B2(n_7),
.C1(n_4),
.C2(n_6),
.Y(n_208)
);

OAI322xp33_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_188),
.A3(n_164),
.B1(n_193),
.B2(n_173),
.C1(n_183),
.C2(n_185),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_4),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_218),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_4),
.B(n_5),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_167),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_166),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_220),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_169),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_177),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_229),
.A2(n_235),
.B1(n_211),
.B2(n_206),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_189),
.B1(n_178),
.B2(n_164),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_196),
.B1(n_201),
.B2(n_214),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_208),
.C(n_198),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_175),
.C(n_176),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_237),
.C(n_203),
.Y(n_245)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_238),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_187),
.B1(n_190),
.B2(n_6),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_10),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_240),
.B1(n_209),
.B2(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_233),
.C(n_221),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_231),
.B1(n_210),
.B2(n_225),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_253),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_252),
.B(n_219),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_265),
.C(n_249),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_251),
.A2(n_238),
.B1(n_223),
.B2(n_224),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_199),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_243),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_227),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_222),
.B(n_225),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_242),
.B(n_218),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_210),
.C(n_217),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_243),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_246),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_205),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_270),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_277),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_267),
.A2(n_248),
.B1(n_249),
.B2(n_247),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_281),
.B1(n_260),
.B2(n_264),
.Y(n_282)
);

OAI221xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_242),
.B1(n_217),
.B2(n_253),
.C(n_229),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_275),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_265),
.B(n_237),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_195),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_278),
.B(n_280),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_195),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_279),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_274),
.B(n_263),
.C(n_244),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_289),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_241),
.C(n_10),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_271),
.A2(n_203),
.B1(n_258),
.B2(n_204),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_279),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_292),
.C(n_284),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_294),
.B(n_295),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_283),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_284),
.B(n_286),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_297),
.Y(n_300)
);

OAI321xp33_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_284),
.A3(n_241),
.B1(n_11),
.B2(n_7),
.C(n_6),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_299),
.B1(n_11),
.B2(n_5),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_300),
.C(n_296),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_5),
.Y(n_303)
);


endmodule