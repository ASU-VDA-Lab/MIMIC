module fake_jpeg_14454_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_7),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_13),
.A2(n_0),
.B1(n_5),
.B2(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_30),
.A2(n_37),
.B1(n_43),
.B2(n_51),
.Y(n_78)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_38),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_18),
.A2(n_8),
.B1(n_10),
.B2(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_5),
.C(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_5),
.B1(n_14),
.B2(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_21),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_25),
.B1(n_24),
.B2(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_15),
.B1(n_21),
.B2(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_32),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_23),
.A2(n_13),
.B1(n_16),
.B2(n_25),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_72),
.Y(n_80)
);

OR2x4_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_17),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_43),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_51),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_77),
.Y(n_87)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_63),
.B1(n_89),
.B2(n_94),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_92),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_35),
.B(n_64),
.C(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_93),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_78),
.B1(n_69),
.B2(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_90),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_62),
.B1(n_58),
.B2(n_61),
.Y(n_90)
);

OR2x6_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_95),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_56),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_58),
.B1(n_68),
.B2(n_59),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_73),
.B1(n_71),
.B2(n_57),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_80),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_108),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_91),
.B1(n_88),
.B2(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_85),
.C(n_96),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_115),
.B1(n_97),
.B2(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_111),
.B(n_98),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_81),
.B1(n_91),
.B2(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_106),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_86),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_116),
.C(n_99),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_91),
.B1(n_93),
.B2(n_79),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_91),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_121),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_120),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_117),
.C(n_101),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_118),
.B1(n_106),
.B2(n_104),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_112),
.C(n_114),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_124),
.C(n_116),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_112),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_127),
.B(n_128),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_132),
.B(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_131),
.B(n_130),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_125),
.Y(n_137)
);


endmodule