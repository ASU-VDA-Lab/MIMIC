module fake_jpeg_19652_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_35),
.B(n_43),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_56),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_57),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_43),
.CON(n_56),
.SN(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_39),
.B1(n_37),
.B2(n_49),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_63),
.B1(n_62),
.B2(n_67),
.Y(n_78)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_71),
.B1(n_64),
.B2(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_39),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_51),
.B1(n_50),
.B2(n_38),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_47),
.B1(n_44),
.B2(n_40),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_20),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_78),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_1),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_93),
.A2(n_77),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_87),
.B(n_83),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_98),
.B1(n_90),
.B2(n_92),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_25),
.B1(n_7),
.B2(n_9),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_89),
.B1(n_92),
.B2(n_94),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_102),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_101),
.C(n_100),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_96),
.B(n_99),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_6),
.B(n_12),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_34),
.B(n_15),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_14),
.C(n_16),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_30),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_24),
.Y(n_111)
);


endmodule