module real_jpeg_25251_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_249;
wire n_176;
wire n_292;
wire n_215;
wire n_221;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_295;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_0),
.B(n_36),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_0),
.B(n_31),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_0),
.B(n_133),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_2),
.B(n_36),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_2),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_3),
.B(n_43),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_3),
.B(n_25),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_45),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_36),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_3),
.B(n_31),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_7),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_7),
.B(n_31),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_7),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_7),
.B(n_36),
.Y(n_236)
);

INVx8_ASAP7_75t_SL g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_10),
.B(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_10),
.B(n_25),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_10),
.B(n_36),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_10),
.B(n_17),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_10),
.B(n_31),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_10),
.B(n_45),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_10),
.B(n_43),
.Y(n_241)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_12),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_12),
.B(n_43),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_25),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_12),
.B(n_36),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_12),
.B(n_31),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_12),
.B(n_45),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_43),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_14),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_14),
.B(n_31),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_15),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_15),
.B(n_45),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_15),
.B(n_36),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_43),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_15),
.B(n_25),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_15),
.B(n_51),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_16),
.B(n_51),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_16),
.B(n_31),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_16),
.B(n_36),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_16),
.B(n_45),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_16),
.B(n_43),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_16),
.B(n_25),
.Y(n_246)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_17),
.Y(n_134)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_17),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_154),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_31),
.Y(n_182)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_38),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_56),
.C(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_35),
.B(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_69),
.SN(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_47),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_70),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_63),
.C(n_69),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_61),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_64),
.C(n_65),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_63),
.B(n_69),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_66),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_69),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_84),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_82),
.C(n_83),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_73),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.C(n_79),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_79),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_83),
.B1(n_91),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_107),
.C(n_111),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_103),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_95),
.B(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_97),
.B(n_103),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.C(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_100),
.B(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.C(n_119),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.C(n_116),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_127),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_297)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_127),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_140),
.C(n_142),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_128),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_136),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_129),
.B(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_131),
.A2(n_132),
.B(n_135),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_131),
.B(n_136),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.C(n_139),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_137),
.B(n_138),
.CI(n_139),
.CON(n_256),
.SN(n_256)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_140),
.B(n_142),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_150),
.C(n_152),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_143),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_144),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_182),
.Y(n_181)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_148),
.B(n_149),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_295),
.C(n_296),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_285),
.C(n_286),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_270),
.C(n_271),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_249),
.C(n_250),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_229),
.C(n_230),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_209),
.C(n_210),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_187),
.C(n_188),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_174),
.C(n_179),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_170),
.B2(n_171),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_172),
.C(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.C(n_183),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_200),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_193),
.C(n_200),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_199),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_208),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_207),
.C(n_208),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_213),
.C(n_218),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_216),
.C(n_217),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_221),
.C(n_222),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_228),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_244),
.C(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_238),
.C(n_239),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_237),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_239),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.CI(n_242),
.CON(n_239),
.SN(n_239)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.CI(n_247),
.CON(n_244),
.SN(n_244)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_254),
.C(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_258),
.C(n_261),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_256),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_266),
.C(n_268),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_266),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_280),
.B2(n_284),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_281),
.C(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_276),
.C(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_293),
.B2(n_294),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_291),
.C(n_293),
.Y(n_295)
);


endmodule