module fake_ibex_297_n_188 (n_7, n_20, n_40, n_17, n_25, n_36, n_41, n_18, n_3, n_22, n_28, n_32, n_39, n_4, n_33, n_5, n_11, n_30, n_6, n_29, n_13, n_2, n_8, n_26, n_35, n_14, n_0, n_9, n_34, n_12, n_38, n_15, n_37, n_24, n_31, n_10, n_23, n_21, n_27, n_19, n_16, n_1, n_188);

input n_7;
input n_20;
input n_40;
input n_17;
input n_25;
input n_36;
input n_41;
input n_18;
input n_3;
input n_22;
input n_28;
input n_32;
input n_39;
input n_4;
input n_33;
input n_5;
input n_11;
input n_30;
input n_6;
input n_29;
input n_13;
input n_2;
input n_8;
input n_26;
input n_35;
input n_14;
input n_0;
input n_9;
input n_34;
input n_12;
input n_38;
input n_15;
input n_37;
input n_24;
input n_31;
input n_10;
input n_23;
input n_21;
input n_27;
input n_19;
input n_16;
input n_1;

output n_188;

wire n_151;
wire n_147;
wire n_85;
wire n_167;
wire n_128;
wire n_84;
wire n_64;
wire n_73;
wire n_152;
wire n_171;
wire n_145;
wire n_65;
wire n_103;
wire n_95;
wire n_139;
wire n_55;
wire n_130;
wire n_63;
wire n_98;
wire n_129;
wire n_161;
wire n_143;
wire n_106;
wire n_177;
wire n_148;
wire n_76;
wire n_118;
wire n_183;
wire n_67;
wire n_164;
wire n_124;
wire n_110;
wire n_47;
wire n_169;
wire n_108;
wire n_82;
wire n_165;
wire n_78;
wire n_60;
wire n_86;
wire n_70;
wire n_87;
wire n_69;
wire n_75;
wire n_109;
wire n_127;
wire n_121;
wire n_175;
wire n_137;
wire n_48;
wire n_57;
wire n_59;
wire n_125;
wire n_178;
wire n_62;
wire n_71;
wire n_153;
wire n_173;
wire n_120;
wire n_93;
wire n_168;
wire n_155;
wire n_162;
wire n_180;
wire n_122;
wire n_116;
wire n_61;
wire n_94;
wire n_134;
wire n_42;
wire n_77;
wire n_112;
wire n_150;
wire n_88;
wire n_133;
wire n_44;
wire n_142;
wire n_51;
wire n_46;
wire n_80;
wire n_172;
wire n_49;
wire n_66;
wire n_74;
wire n_90;
wire n_176;
wire n_58;
wire n_43;
wire n_140;
wire n_136;
wire n_119;
wire n_100;
wire n_179;
wire n_72;
wire n_166;
wire n_163;
wire n_114;
wire n_97;
wire n_102;
wire n_181;
wire n_131;
wire n_123;
wire n_52;
wire n_99;
wire n_135;
wire n_105;
wire n_156;
wire n_126;
wire n_187;
wire n_154;
wire n_182;
wire n_111;
wire n_104;
wire n_141;
wire n_89;
wire n_83;
wire n_53;
wire n_107;
wire n_115;
wire n_149;
wire n_54;
wire n_186;
wire n_50;
wire n_92;
wire n_144;
wire n_170;
wire n_101;
wire n_113;
wire n_138;
wire n_96;
wire n_185;
wire n_68;
wire n_117;
wire n_79;
wire n_81;
wire n_159;
wire n_158;
wire n_132;
wire n_174;
wire n_157;
wire n_160;
wire n_184;
wire n_56;
wire n_146;
wire n_91;
wire n_45;

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

INVxp67_ASAP7_75t_SL g75 ( 
.A(n_22),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_6),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g79 ( 
.A(n_25),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_1),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_10),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_3),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_11),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_5),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_5),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_6),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_44),
.A2(n_34),
.B1(n_41),
.B2(n_64),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_44),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_78),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_76),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

OAI221xp5_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_79),
.B1(n_80),
.B2(n_51),
.C(n_66),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

OR2x6_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_57),
.B(n_62),
.Y(n_110)
);

OR2x6_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_53),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_74),
.B1(n_59),
.B2(n_43),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_43),
.B(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_43),
.B(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_55),
.B(n_43),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_55),
.B(n_43),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_107),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_114),
.Y(n_121)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_81),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_100),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_112),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_84),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_96),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_91),
.B(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_89),
.B(n_117),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_117),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_94),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_88),
.B(n_90),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_86),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_99),
.B(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_83),
.B(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_83),
.B(n_106),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_83),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_83),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_83),
.B(n_137),
.Y(n_144)
);

CKINVDCx11_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_123),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_133),
.B(n_130),
.C(n_121),
.Y(n_154)
);

OAI21x1_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_141),
.B(n_140),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_132),
.B1(n_139),
.B2(n_142),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_147),
.Y(n_160)
);

OR2x6_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_157),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_R g167 ( 
.A(n_145),
.B(n_153),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_152),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_153),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_151),
.B1(n_149),
.B2(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_150),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_170),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_170),
.B1(n_174),
.B2(n_160),
.Y(n_179)
);

INVxp33_ASAP7_75t_SL g180 ( 
.A(n_179),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_175),
.C(n_178),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_181),
.B(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_173),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_161),
.B(n_166),
.Y(n_185)
);

AOI31xp33_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_184),
.A3(n_163),
.B(n_172),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_176),
.B1(n_171),
.B2(n_172),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_155),
.B1(n_176),
.B2(n_171),
.C(n_177),
.Y(n_188)
);


endmodule