module fake_netlist_6_1615_n_2427 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2427);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2427;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_873;
wire n_461;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_437;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_1070;
wire n_458;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_1207;
wire n_811;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_2416;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2301;
wire n_2209;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_2420;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_SL g238 ( 
.A(n_225),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_120),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_19),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_135),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_176),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_185),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_180),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_86),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_110),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_102),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_129),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_96),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_165),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_60),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_24),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_5),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_119),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_89),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_127),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_143),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_83),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_19),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_26),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_34),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_201),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_74),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_109),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_213),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_134),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_77),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_79),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_27),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_221),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_85),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_30),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_218),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_10),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_35),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_48),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_100),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_138),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_22),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_70),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_72),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_162),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_99),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_121),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_13),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_228),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_24),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_48),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_195),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_51),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_155),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_12),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_91),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_184),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_36),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_1),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_0),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_118),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_12),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_115),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_202),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_94),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_183),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_146),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_196),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_56),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_44),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_14),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_60),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_223),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_45),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_206),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_30),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_71),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_29),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_36),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_74),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_82),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_43),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_156),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_124),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_207),
.Y(n_332)
);

BUFx8_ASAP7_75t_SL g333 ( 
.A(n_29),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_41),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_126),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_39),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_11),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_178),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_107),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_101),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_50),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_77),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_232),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_137),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_76),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_37),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_113),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_80),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_214),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_44),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_43),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_147),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_104),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_25),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_10),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_84),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_160),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_69),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_18),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_2),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_45),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_105),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_16),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_205),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_32),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_173),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_72),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_192),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_106),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_37),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_80),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_90),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_32),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_174),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_210),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_79),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_204),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_108),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_161),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_53),
.Y(n_380)
);

BUFx5_ASAP7_75t_L g381 ( 
.A(n_87),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_190),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_70),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_38),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_139),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_34),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_144),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_211),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_53),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_217),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_97),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_193),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_111),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_212),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_20),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_148),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_237),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_154),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_158),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_46),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_58),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_131),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_65),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_13),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_235),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_125),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_92),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_179),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_230),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_76),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_68),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_26),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_73),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_136),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_0),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_31),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_73),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_181),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_20),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_22),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_166),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_88),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_114),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_149),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_159),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_224),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_38),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_23),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_199),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_27),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_54),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_175),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_123),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_64),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_1),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_197),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_46),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_61),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_61),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_152),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_132),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_140),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_35),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_28),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_6),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_33),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_15),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_47),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_7),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_216),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_75),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_68),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_57),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_186),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_62),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_103),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_31),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_169),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_21),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_116),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_56),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_3),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_57),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_6),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_18),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_130),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_348),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_348),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_263),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_302),
.Y(n_470)
);

BUFx5_ASAP7_75t_L g471 ( 
.A(n_270),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_348),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_333),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_348),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_348),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_256),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_288),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_459),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_320),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_462),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_254),
.Y(n_486)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_256),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_292),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_374),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_405),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_392),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_293),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_414),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_462),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_296),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_299),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_267),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_267),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_329),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_329),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_364),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_334),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_334),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_441),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_345),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_345),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_355),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_355),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_332),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_360),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_274),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_360),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_377),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_449),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_282),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_449),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_282),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_301),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_304),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_456),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_245),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_243),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_245),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_265),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_308),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_310),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_308),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_352),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_269),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_280),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_298),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_321),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_326),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_336),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_337),
.Y(n_537)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_284),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_346),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_257),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_312),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_313),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_351),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_365),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_370),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_380),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_383),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_389),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_314),
.Y(n_549)
);

INVxp33_ASAP7_75t_SL g550 ( 
.A(n_258),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_410),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_352),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_315),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_322),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_258),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_282),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_274),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_415),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_417),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_272),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_331),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_338),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_444),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_447),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_343),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_344),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_347),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_353),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_451),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_452),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_335),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_282),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_268),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_268),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_356),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_273),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_273),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_303),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_303),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_362),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_368),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_274),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_339),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_369),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_339),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_366),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_366),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_382),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_382),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_375),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_418),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_335),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_335),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_469),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_475),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_523),
.B(n_238),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_477),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_475),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_488),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_496),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_553),
.B(n_238),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_553),
.B(n_255),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_517),
.B(n_261),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_496),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_467),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_484),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_527),
.B(n_255),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_467),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_R g612 ( 
.A(n_487),
.B(n_239),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_553),
.B(n_425),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_472),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_517),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_519),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_494),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_474),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_474),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_478),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_478),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_513),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_479),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_519),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_479),
.B(n_425),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_529),
.B(n_239),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_530),
.B(n_241),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_480),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_481),
.B(n_398),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_525),
.B(n_398),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_481),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_557),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_503),
.B(n_261),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_482),
.B(n_241),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_557),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_483),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_483),
.B(n_271),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_485),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_485),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_489),
.B(n_242),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_489),
.Y(n_645)
);

NOR2xp67_ASAP7_75t_L g646 ( 
.A(n_574),
.B(n_277),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_491),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_491),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_476),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_574),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_575),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_525),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_575),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_576),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_576),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_578),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_578),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_490),
.A2(n_285),
.B1(n_359),
.B2(n_240),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_579),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_579),
.B(n_242),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_580),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_580),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_581),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_581),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_585),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_585),
.B(n_244),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_587),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_587),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_573),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_588),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_588),
.B(n_281),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_589),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_589),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_590),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_590),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_591),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_591),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_516),
.B(n_294),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_532),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_471),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_471),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_SL g682 ( 
.A1(n_493),
.A2(n_376),
.B1(n_400),
.B2(n_371),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_497),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_532),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_499),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_516),
.B(n_311),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_499),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_471),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_518),
.B(n_340),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_498),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_520),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_500),
.A2(n_372),
.B(n_357),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_533),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_518),
.B(n_244),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_611),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_598),
.B(n_521),
.Y(n_696)
);

AOI22x1_ASAP7_75t_L g697 ( 
.A1(n_689),
.A2(n_486),
.B1(n_495),
.B2(n_492),
.Y(n_697)
);

NOR2x1p5_ASAP7_75t_L g698 ( 
.A(n_599),
.B(n_473),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_598),
.B(n_528),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_611),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_606),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_613),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_596),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_652),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_637),
.B(n_538),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_678),
.B(n_387),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_613),
.Y(n_707)
);

NAND3xp33_ASAP7_75t_L g708 ( 
.A(n_689),
.B(n_562),
.C(n_506),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_616),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_652),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_637),
.A2(n_511),
.B1(n_515),
.B2(n_540),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_694),
.B(n_388),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_606),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_637),
.B(n_541),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_606),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_628),
.B(n_554),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_615),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_615),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_615),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_622),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_628),
.A2(n_290),
.B1(n_305),
.B2(n_276),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_630),
.A2(n_542),
.B1(n_549),
.B2(n_550),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_598),
.B(n_555),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_620),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_622),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_620),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_623),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_652),
.Y(n_729)
);

AND2x6_ASAP7_75t_L g730 ( 
.A(n_609),
.B(n_261),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_620),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_621),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_617),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_630),
.A2(n_563),
.B1(n_567),
.B2(n_564),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_621),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_621),
.Y(n_736)
);

AOI22x1_ASAP7_75t_L g737 ( 
.A1(n_689),
.A2(n_556),
.B1(n_470),
.B2(n_266),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_623),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_617),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_650),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_617),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_625),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_625),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_629),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_629),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_601),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_624),
.Y(n_747)
);

INVx8_ASAP7_75t_L g748 ( 
.A(n_605),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_631),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_650),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_629),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_619),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_626),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_683),
.B(n_568),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_636),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_609),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_649),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_658),
.B(n_682),
.C(n_584),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_636),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_631),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_650),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_609),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_641),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_650),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_634),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_690),
.B(n_569),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_650),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_617),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_649),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_691),
.B(n_522),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_669),
.B(n_570),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_650),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_L g773 ( 
.A(n_694),
.B(n_573),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_634),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_647),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_640),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_669),
.B(n_577),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_608),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_626),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_647),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_640),
.Y(n_782)
);

AO21x2_ASAP7_75t_L g783 ( 
.A1(n_692),
.A2(n_391),
.B(n_390),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_648),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_669),
.B(n_582),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_681),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_633),
.B(n_500),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_624),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_669),
.B(n_583),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_641),
.Y(n_790)
);

AND3x2_ASAP7_75t_L g791 ( 
.A(n_633),
.B(n_318),
.C(n_558),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_638),
.B(n_586),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_638),
.B(n_592),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_681),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_669),
.B(n_593),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_626),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_603),
.B(n_526),
.C(n_524),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_669),
.B(n_471),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_618),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_640),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_669),
.B(n_594),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_642),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_612),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_626),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_633),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_642),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_R g807 ( 
.A(n_678),
.B(n_246),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_648),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_618),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_618),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_626),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_626),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_644),
.B(n_471),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_626),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_658),
.B(n_342),
.C(n_341),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_618),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_635),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_597),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_644),
.B(n_594),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_660),
.B(n_595),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_678),
.B(n_394),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_660),
.B(n_261),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_627),
.B(n_471),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_627),
.Y(n_824)
);

INVx5_ASAP7_75t_L g825 ( 
.A(n_605),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_635),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_635),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_635),
.Y(n_828)
);

BUFx6f_ASAP7_75t_SL g829 ( 
.A(n_678),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_681),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_639),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_686),
.B(n_501),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_642),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_627),
.B(n_471),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_639),
.Y(n_835)
);

BUFx10_ASAP7_75t_L g836 ( 
.A(n_686),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_682),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_645),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_645),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_627),
.B(n_471),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_639),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_646),
.A2(n_407),
.B(n_399),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_641),
.B(n_471),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_641),
.B(n_595),
.Y(n_844)
);

AOI21x1_ASAP7_75t_L g845 ( 
.A1(n_646),
.A2(n_424),
.B(n_423),
.Y(n_845)
);

NOR2x1p5_ASAP7_75t_L g846 ( 
.A(n_666),
.B(n_259),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_639),
.Y(n_847)
);

INVx5_ASAP7_75t_L g848 ( 
.A(n_605),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_666),
.B(n_385),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_597),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_686),
.B(n_385),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_671),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_632),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_686),
.B(n_349),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_671),
.B(n_426),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_645),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_632),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_632),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_696),
.B(n_361),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_699),
.B(n_431),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_717),
.B(n_603),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_756),
.B(n_604),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_756),
.B(n_604),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_786),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_786),
.B(n_261),
.Y(n_865)
);

OR2x6_ASAP7_75t_L g866 ( 
.A(n_747),
.B(n_531),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_762),
.B(n_693),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_762),
.B(n_693),
.Y(n_868)
);

XNOR2xp5_ASAP7_75t_L g869 ( 
.A(n_703),
.B(n_434),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_853),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_792),
.B(n_614),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_786),
.A2(n_681),
.B(n_680),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_713),
.A2(n_671),
.B1(n_632),
.B2(n_692),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_824),
.B(n_614),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_724),
.B(n_397),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_695),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_786),
.B(n_262),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_853),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_763),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_824),
.A2(n_432),
.B1(n_450),
.B2(n_429),
.Y(n_880)
);

NAND3x1_ASAP7_75t_L g881 ( 
.A(n_758),
.B(n_537),
.C(n_536),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_857),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_829),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_695),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_805),
.Y(n_885)
);

AO22x2_ASAP7_75t_L g886 ( 
.A1(n_815),
.A2(n_460),
.B1(n_466),
.B2(n_454),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_794),
.B(n_262),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_711),
.B(n_671),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_L g889 ( 
.A(n_730),
.B(n_803),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_700),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_819),
.B(n_665),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_700),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_805),
.B(n_715),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_854),
.B(n_665),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_857),
.B(n_665),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_787),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_858),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_858),
.B(n_665),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_852),
.B(n_668),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_787),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_747),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_832),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_852),
.B(n_668),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_788),
.B(n_679),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_734),
.B(n_246),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_852),
.B(n_668),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_757),
.B(n_679),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_711),
.B(n_668),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_729),
.B(n_680),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_702),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_794),
.B(n_262),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_816),
.Y(n_912)
);

AND2x6_ASAP7_75t_L g913 ( 
.A(n_763),
.B(n_262),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_832),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_729),
.B(n_680),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_794),
.B(n_262),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_794),
.B(n_287),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_813),
.B(n_688),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_702),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_830),
.B(n_287),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_763),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_707),
.B(n_709),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_707),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_788),
.B(n_684),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_790),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_709),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_769),
.B(n_684),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_790),
.Y(n_928)
);

NOR2xp67_ASAP7_75t_L g929 ( 
.A(n_746),
.B(n_654),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_710),
.B(n_688),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_713),
.A2(n_692),
.B1(n_605),
.B2(n_381),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_697),
.B(n_286),
.C(n_283),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_830),
.B(n_287),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_710),
.B(n_688),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_790),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_721),
.B(n_685),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_721),
.B(n_685),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_713),
.A2(n_605),
.B1(n_381),
.B2(n_282),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_726),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_726),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_728),
.Y(n_941)
);

INVx8_ASAP7_75t_L g942 ( 
.A(n_829),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_728),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_836),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_738),
.B(n_685),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_830),
.B(n_287),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_830),
.B(n_287),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_773),
.B(n_539),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_773),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_738),
.B(n_685),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_836),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_712),
.B(n_543),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_742),
.B(n_685),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_742),
.B(n_685),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_743),
.B(n_661),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_743),
.B(n_661),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_846),
.B(n_465),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_L g958 ( 
.A(n_730),
.B(n_282),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_836),
.B(n_330),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_749),
.B(n_661),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_749),
.B(n_661),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_760),
.B(n_661),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_708),
.B(n_544),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_713),
.A2(n_605),
.B1(n_381),
.B2(n_282),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_760),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_765),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_708),
.B(n_545),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_705),
.B(n_247),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_765),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_836),
.B(n_330),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_723),
.B(n_533),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_774),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_774),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_820),
.B(n_704),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_775),
.B(n_661),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_846),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_775),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_752),
.B(n_534),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_781),
.B(n_674),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_781),
.B(n_674),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_784),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_722),
.B(n_535),
.C(n_534),
.Y(n_982)
);

AND2x2_ASAP7_75t_SL g983 ( 
.A(n_793),
.B(n_330),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_713),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_784),
.B(n_674),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_849),
.B(n_247),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_823),
.B(n_330),
.Y(n_987)
);

AO22x1_ASAP7_75t_L g988 ( 
.A1(n_844),
.A2(n_266),
.B1(n_275),
.B2(n_259),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_754),
.B(n_248),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_834),
.B(n_330),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_808),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_808),
.B(n_706),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_706),
.B(n_674),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_706),
.B(n_674),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_840),
.B(n_396),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_706),
.B(n_674),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_821),
.B(n_687),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_701),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_816),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_821),
.B(n_687),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_821),
.B(n_687),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_701),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_843),
.B(n_396),
.Y(n_1003)
);

INVxp33_ASAP7_75t_SL g1004 ( 
.A(n_770),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_714),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_821),
.B(n_855),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_816),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_855),
.B(n_687),
.Y(n_1008)
);

AND2x6_ASAP7_75t_SL g1009 ( 
.A(n_837),
.B(n_535),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_766),
.B(n_546),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_714),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_807),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_737),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_797),
.A2(n_547),
.B(n_548),
.C(n_546),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_851),
.B(n_248),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_855),
.B(n_791),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_716),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_855),
.B(n_816),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_827),
.Y(n_1019)
);

INVxp67_ASAP7_75t_SL g1020 ( 
.A(n_827),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_827),
.B(n_396),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_730),
.B(n_687),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_829),
.B(n_249),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_697),
.Y(n_1024)
);

BUFx8_ASAP7_75t_L g1025 ( 
.A(n_730),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_827),
.B(n_249),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_748),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_835),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_835),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_835),
.B(n_825),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_730),
.B(n_687),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_835),
.B(n_250),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_730),
.A2(n_422),
.B1(n_433),
.B2(n_421),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_896),
.B(n_698),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_870),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_871),
.B(n_730),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_876),
.Y(n_1037)
);

BUFx2_ASAP7_75t_SL g1038 ( 
.A(n_929),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_878),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_885),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_902),
.B(n_698),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_861),
.B(n_740),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_951),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_885),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_SL g1045 ( 
.A1(n_1004),
.A2(n_779),
.B1(n_350),
.B2(n_384),
.Y(n_1045)
);

INVxp67_ASAP7_75t_SL g1046 ( 
.A(n_879),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_876),
.Y(n_1047)
);

INVx5_ASAP7_75t_L g1048 ( 
.A(n_951),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_907),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_951),
.B(n_825),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1012),
.B(n_797),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_893),
.A2(n_778),
.B1(n_785),
.B2(n_771),
.Y(n_1052)
);

BUFx10_ASAP7_75t_L g1053 ( 
.A(n_1023),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_893),
.B(n_740),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_862),
.B(n_740),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_882),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_884),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_951),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_863),
.B(n_740),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_879),
.Y(n_1060)
);

AO21x1_ASAP7_75t_L g1061 ( 
.A1(n_905),
.A2(n_822),
.B(n_801),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_983),
.A2(n_737),
.B1(n_783),
.B2(n_282),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_884),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_883),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_869),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_983),
.A2(n_783),
.B1(n_381),
.B2(n_396),
.Y(n_1066)
);

AND3x2_ASAP7_75t_SL g1067 ( 
.A(n_886),
.B(n_350),
.C(n_275),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_890),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_890),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_901),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_875),
.B(n_867),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_914),
.B(n_547),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_1009),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_900),
.B(n_548),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_897),
.Y(n_1075)
);

AND3x2_ASAP7_75t_SL g1076 ( 
.A(n_886),
.B(n_386),
.C(n_384),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_978),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_957),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_875),
.A2(n_655),
.B(n_656),
.C(n_654),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_883),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_868),
.B(n_750),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_864),
.B(n_825),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_892),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_892),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_859),
.B(n_750),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_866),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_866),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_864),
.B(n_825),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_904),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_910),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_992),
.A2(n_750),
.B1(n_764),
.B2(n_761),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_910),
.Y(n_1092)
);

NOR2x1p5_ASAP7_75t_L g1093 ( 
.A(n_952),
.B(n_386),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_924),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_874),
.A2(n_748),
.B(n_789),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1024),
.B(n_859),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_919),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_888),
.B(n_825),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_948),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_860),
.B(n_750),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_883),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_866),
.Y(n_1102)
);

AND2x6_ASAP7_75t_SL g1103 ( 
.A(n_905),
.B(n_551),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_860),
.B(n_761),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_939),
.B(n_943),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_919),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_949),
.B(n_551),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_927),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_923),
.Y(n_1109)
);

CKINVDCx14_ASAP7_75t_R g1110 ( 
.A(n_1016),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_888),
.B(n_1006),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_SL g1112 ( 
.A(n_984),
.B(n_783),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_918),
.A2(n_810),
.B(n_809),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_888),
.B(n_825),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_926),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_L g1116 ( 
.A1(n_891),
.A2(n_845),
.B(n_842),
.C(n_718),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_965),
.B(n_969),
.Y(n_1117)
);

AO22x1_ASAP7_75t_L g1118 ( 
.A1(n_989),
.A2(n_401),
.B1(n_403),
.B2(n_395),
.Y(n_1118)
);

INVx3_ASAP7_75t_SL g1119 ( 
.A(n_942),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_926),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_940),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1010),
.B(n_552),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_940),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_942),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1027),
.B(n_848),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_1027),
.B(n_848),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_974),
.A2(n_795),
.B1(n_764),
.B2(n_767),
.Y(n_1127)
);

AO21x1_ASAP7_75t_L g1128 ( 
.A1(n_968),
.A2(n_845),
.B(n_842),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_941),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_971),
.B(n_552),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_SL g1131 ( 
.A(n_942),
.B(n_385),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_974),
.A2(n_764),
.B1(n_767),
.B2(n_761),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_941),
.B(n_848),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1014),
.A2(n_810),
.B(n_817),
.C(n_809),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_972),
.B(n_761),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_944),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_966),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_930),
.A2(n_826),
.B(n_817),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_966),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_991),
.B(n_921),
.Y(n_1140)
);

BUFx8_ASAP7_75t_L g1141 ( 
.A(n_976),
.Y(n_1141)
);

NAND2x1p5_ASAP7_75t_L g1142 ( 
.A(n_944),
.B(n_848),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_881),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_973),
.B(n_764),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_989),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_991),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_977),
.B(n_767),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_886),
.A2(n_381),
.B1(n_396),
.B2(n_718),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_963),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_981),
.B(n_767),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_988),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_922),
.B(n_772),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_999),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1007),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1019),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_967),
.B(n_559),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_925),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1028),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_894),
.B(n_772),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_928),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1029),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1013),
.B(n_772),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_982),
.A2(n_381),
.B1(n_720),
.B2(n_719),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_998),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_968),
.B(n_772),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1018),
.B(n_848),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_935),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1018),
.A2(n_804),
.B1(n_811),
.B2(n_780),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_912),
.B(n_826),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1002),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_986),
.B(n_559),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1016),
.B(n_560),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_913),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_986),
.B(n_780),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1015),
.B(n_560),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_932),
.A2(n_804),
.B1(n_811),
.B2(n_780),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_899),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1015),
.B(n_561),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1020),
.B(n_828),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1023),
.B(n_561),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1005),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1011),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_903),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1011),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1014),
.A2(n_831),
.B(n_841),
.C(n_828),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1026),
.B(n_831),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1017),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1017),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_913),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1026),
.B(n_841),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_906),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_895),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_898),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1032),
.B(n_847),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_936),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_937),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_945),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_950),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1032),
.B(n_847),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_953),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_934),
.B(n_780),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_880),
.B(n_251),
.C(n_250),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_938),
.A2(n_381),
.B1(n_720),
.B2(n_719),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_889),
.A2(n_811),
.B1(n_812),
.B2(n_804),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_954),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_955),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_956),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_909),
.B(n_915),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1030),
.B(n_565),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_960),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_961),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_993),
.A2(n_811),
.B1(n_812),
.B2(n_804),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_908),
.B(n_873),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_SL g1214 ( 
.A1(n_964),
.A2(n_401),
.B1(n_403),
.B2(n_395),
.Y(n_1214)
);

INVxp33_ASAP7_75t_L g1215 ( 
.A(n_1003),
.Y(n_1215)
);

BUFx4f_ASAP7_75t_L g1216 ( 
.A(n_913),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_962),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_975),
.B(n_812),
.Y(n_1218)
);

OR2x2_ASAP7_75t_SL g1219 ( 
.A(n_994),
.B(n_565),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_931),
.A2(n_812),
.B1(n_814),
.B2(n_748),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_979),
.B(n_814),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_980),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_985),
.Y(n_1223)
);

INVx5_ASAP7_75t_L g1224 ( 
.A(n_913),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1071),
.B(n_1025),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_1058),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1149),
.B(n_865),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1170),
.Y(n_1228)
);

INVx3_ASAP7_75t_SL g1229 ( 
.A(n_1080),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1083),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1096),
.B(n_865),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1156),
.B(n_877),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1145),
.A2(n_996),
.B1(n_970),
.B2(n_959),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1040),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1175),
.B(n_877),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1208),
.A2(n_872),
.B(n_997),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1077),
.B(n_887),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1070),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1122),
.B(n_887),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1094),
.B(n_911),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1213),
.A2(n_1001),
.B(n_1000),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1089),
.B(n_1025),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1040),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1090),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1058),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1042),
.A2(n_1008),
.B(n_970),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1066),
.A2(n_959),
.B(n_916),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1051),
.A2(n_1033),
.B1(n_916),
.B2(n_917),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1094),
.B(n_911),
.Y(n_1249)
);

OR2x6_ASAP7_75t_L g1250 ( 
.A(n_1064),
.B(n_748),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1108),
.B(n_917),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1064),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1049),
.B(n_566),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1186),
.A2(n_933),
.B(n_920),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1064),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1170),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1190),
.A2(n_933),
.B(n_920),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1079),
.A2(n_1117),
.B(n_1105),
.C(n_1104),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1194),
.A2(n_947),
.B(n_946),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1044),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1099),
.B(n_946),
.Y(n_1261)
);

BUFx12f_ASAP7_75t_L g1262 ( 
.A(n_1064),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1099),
.B(n_947),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1199),
.A2(n_1003),
.B(n_990),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1051),
.B(n_1030),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1101),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1097),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1036),
.A2(n_1095),
.B(n_1165),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1106),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1079),
.A2(n_987),
.B(n_995),
.C(n_990),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1095),
.A2(n_995),
.B(n_987),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1180),
.B(n_566),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1177),
.B(n_913),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1044),
.B(n_1171),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1178),
.A2(n_1021),
.B(n_958),
.C(n_727),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1119),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1165),
.A2(n_1031),
.B(n_1022),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1065),
.B(n_814),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1113),
.A2(n_1021),
.B(n_727),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1058),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1177),
.B(n_814),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1093),
.A2(n_440),
.B1(n_442),
.B2(n_436),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1058),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1085),
.A2(n_731),
.B(n_732),
.C(n_725),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1086),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1085),
.A2(n_850),
.B(n_739),
.C(n_741),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1037),
.Y(n_1287)
);

AO32x1_ASAP7_75t_L g1288 ( 
.A1(n_1091),
.A2(n_572),
.A3(n_571),
.B1(n_502),
.B2(n_504),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1130),
.B(n_251),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1172),
.B(n_571),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1100),
.A2(n_850),
.B(n_739),
.C(n_741),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1100),
.A2(n_850),
.B(n_739),
.C(n_741),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1119),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1087),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1046),
.A2(n_748),
.B1(n_796),
.B2(n_753),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1115),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1121),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1041),
.A2(n_253),
.B1(n_260),
.B2(n_252),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1111),
.A2(n_796),
.B(n_753),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1111),
.A2(n_796),
.B(n_753),
.Y(n_1300)
);

NAND2xp33_ASAP7_75t_SL g1301 ( 
.A(n_1101),
.B(n_1078),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1172),
.A2(n_412),
.B(n_411),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1143),
.B(n_1045),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1183),
.B(n_850),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1053),
.B(n_1038),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1102),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1183),
.B(n_1025),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1035),
.B(n_655),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1107),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1039),
.B(n_656),
.Y(n_1310)
);

CKINVDCx16_ASAP7_75t_R g1311 ( 
.A(n_1124),
.Y(n_1311)
);

INVx11_ASAP7_75t_L g1312 ( 
.A(n_1141),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1123),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1174),
.A2(n_1138),
.B(n_1046),
.Y(n_1314)
);

BUFx4f_ASAP7_75t_L g1315 ( 
.A(n_1101),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1174),
.A2(n_796),
.B1(n_753),
.B2(n_253),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1101),
.Y(n_1317)
);

AOI21x1_ASAP7_75t_SL g1318 ( 
.A1(n_1162),
.A2(n_798),
.B(n_381),
.Y(n_1318)
);

OAI21xp33_ASAP7_75t_L g1319 ( 
.A1(n_1131),
.A2(n_412),
.B(n_411),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1054),
.A2(n_1112),
.B(n_1075),
.C(n_1056),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1047),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1041),
.B(n_572),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1201),
.A2(n_796),
.B(n_753),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1054),
.B(n_657),
.Y(n_1324)
);

AOI33xp33_ASAP7_75t_L g1325 ( 
.A1(n_1074),
.A2(n_501),
.A3(n_514),
.B1(n_512),
.B2(n_510),
.B3(n_509),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_SL g1326 ( 
.A(n_1073),
.B(n_252),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1057),
.Y(n_1327)
);

OR2x6_ASAP7_75t_SL g1328 ( 
.A(n_1151),
.B(n_413),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1201),
.A2(n_818),
.B(n_768),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1063),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1140),
.A2(n_759),
.B(n_839),
.C(n_838),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1107),
.B(n_502),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1152),
.A2(n_818),
.B(n_768),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1159),
.A2(n_818),
.B(n_768),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1140),
.A2(n_1202),
.B(n_1137),
.C(n_1146),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1060),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1068),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1202),
.A2(n_260),
.B1(n_409),
.B2(n_458),
.Y(n_1338)
);

INVx4_ASAP7_75t_L g1339 ( 
.A(n_1043),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1069),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1034),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1084),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1139),
.A2(n_755),
.B(n_839),
.C(n_838),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1072),
.B(n_504),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1092),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1128),
.A2(n_731),
.B(n_725),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1192),
.B(n_1193),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1053),
.B(n_289),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1109),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1081),
.A2(n_818),
.B(n_799),
.Y(n_1350)
);

NOR2x1_ASAP7_75t_L g1351 ( 
.A(n_1034),
.B(n_733),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1195),
.A2(n_755),
.B(n_833),
.C(n_806),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1043),
.B(n_264),
.Y(n_1353)
);

NOR3xp33_ASAP7_75t_SL g1354 ( 
.A(n_1214),
.B(n_448),
.C(n_413),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1110),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1052),
.A2(n_264),
.B1(n_278),
.B2(n_279),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1197),
.B(n_657),
.Y(n_1357)
);

AO21x1_ASAP7_75t_L g1358 ( 
.A1(n_1112),
.A2(n_735),
.B(n_732),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1060),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1072),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1118),
.B(n_295),
.C(n_291),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1198),
.B(n_670),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_SL g1363 ( 
.A(n_1062),
.B(n_453),
.C(n_448),
.Y(n_1363)
);

AND3x4_ASAP7_75t_L g1364 ( 
.A(n_1074),
.B(n_455),
.C(n_453),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1120),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1129),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1103),
.B(n_297),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1218),
.A2(n_799),
.B(n_733),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1209),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1043),
.B(n_278),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1066),
.A2(n_279),
.B1(n_378),
.B2(n_379),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1110),
.B(n_300),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1164),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1200),
.B(n_670),
.Y(n_1374)
);

INVxp67_ASAP7_75t_SL g1375 ( 
.A(n_1060),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_SL g1376 ( 
.A(n_1043),
.B(n_378),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1141),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1209),
.B(n_505),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1055),
.A2(n_818),
.B(n_799),
.Y(n_1379)
);

NOR3xp33_ASAP7_75t_SL g1380 ( 
.A(n_1067),
.B(n_457),
.C(n_455),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1219),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_R g1382 ( 
.A(n_1157),
.B(n_379),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1167),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1205),
.B(n_672),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1215),
.A2(n_733),
.B(n_673),
.C(n_677),
.Y(n_1385)
);

INVx5_ASAP7_75t_L g1386 ( 
.A(n_1048),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1048),
.A2(n_393),
.B1(n_402),
.B2(n_406),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1215),
.B(n_306),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1060),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1181),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1207),
.B(n_672),
.Y(n_1391)
);

O2A1O1Ixp5_ASAP7_75t_L g1392 ( 
.A1(n_1358),
.A2(n_1061),
.B(n_1116),
.C(n_1050),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1238),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1268),
.A2(n_1218),
.A3(n_1220),
.B(n_1211),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1315),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1312),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1373),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1265),
.A2(n_1062),
.B1(n_1148),
.B2(n_1048),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1347),
.B(n_1210),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1367),
.A2(n_1153),
.B(n_1155),
.C(n_1154),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1379),
.A2(n_1334),
.B(n_1333),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1315),
.Y(n_1402)
);

AO21x1_ASAP7_75t_L g1403 ( 
.A1(n_1258),
.A2(n_1185),
.B(n_1134),
.Y(n_1403)
);

AOI221x1_ASAP7_75t_L g1404 ( 
.A1(n_1363),
.A2(n_1067),
.B1(n_1076),
.B2(n_1217),
.C(n_1221),
.Y(n_1404)
);

CKINVDCx6p67_ASAP7_75t_R g1405 ( 
.A(n_1229),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1272),
.B(n_1206),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1324),
.B(n_1222),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1255),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1248),
.A2(n_1148),
.B1(n_1048),
.B2(n_1216),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1234),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1346),
.A2(n_1059),
.B(n_1135),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1390),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1235),
.B(n_1223),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1379),
.A2(n_1116),
.B(n_1134),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1334),
.A2(n_1185),
.B(n_1147),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_SL g1416 ( 
.A1(n_1307),
.A2(n_1150),
.B(n_1144),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1247),
.A2(n_1127),
.B(n_1191),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1333),
.A2(n_1204),
.B(n_1176),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1314),
.A2(n_1136),
.B(n_1169),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1314),
.A2(n_1136),
.B(n_1179),
.Y(n_1420)
);

OAI22x1_ASAP7_75t_L g1421 ( 
.A1(n_1381),
.A2(n_1076),
.B1(n_1160),
.B2(n_1157),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1268),
.A2(n_1184),
.A3(n_1188),
.B(n_1187),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1350),
.A2(n_1212),
.B(n_1132),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1357),
.B(n_1196),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1350),
.A2(n_1182),
.B(n_1160),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1318),
.A2(n_1142),
.B(n_1158),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1290),
.B(n_1161),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1341),
.B(n_1136),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1243),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1318),
.A2(n_1142),
.B(n_1126),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_1305),
.B(n_1136),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1299),
.A2(n_1300),
.B(n_1329),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1274),
.A2(n_1216),
.B1(n_1189),
.B2(n_1173),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1299),
.A2(n_1300),
.B(n_1329),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1254),
.A2(n_1163),
.B(n_1168),
.Y(n_1435)
);

AND2x2_ASAP7_75t_SL g1436 ( 
.A(n_1303),
.B(n_1173),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1285),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1254),
.A2(n_1163),
.B(n_1203),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1362),
.B(n_1098),
.Y(n_1439)
);

AOI221x1_ASAP7_75t_L g1440 ( 
.A1(n_1363),
.A2(n_1189),
.B1(n_673),
.B2(n_677),
.C(n_507),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1258),
.A2(n_1098),
.B(n_1114),
.C(n_1203),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1320),
.A2(n_1133),
.B(n_1050),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1278),
.B(n_1133),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1309),
.B(n_1114),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1241),
.A2(n_1126),
.B(n_1125),
.Y(n_1445)
);

AO21x1_ASAP7_75t_L g1446 ( 
.A1(n_1233),
.A2(n_1166),
.B(n_1082),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1241),
.A2(n_1125),
.B(n_1082),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1332),
.B(n_505),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1230),
.Y(n_1449)
);

AO31x2_ASAP7_75t_L g1450 ( 
.A1(n_1271),
.A2(n_759),
.A3(n_735),
.B(n_736),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1253),
.B(n_507),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1244),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1236),
.A2(n_1088),
.B(n_1224),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1374),
.B(n_1166),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1252),
.B(n_1224),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1267),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1384),
.B(n_1088),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1236),
.A2(n_1224),
.B(n_848),
.Y(n_1458)
);

AOI221x1_ASAP7_75t_L g1459 ( 
.A1(n_1271),
.A2(n_509),
.B1(n_514),
.B2(n_512),
.C(n_510),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1239),
.A2(n_1224),
.B1(n_457),
.B2(n_461),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1261),
.A2(n_458),
.B(n_393),
.C(n_402),
.Y(n_1461)
);

OAI21xp33_ASAP7_75t_L g1462 ( 
.A1(n_1338),
.A2(n_463),
.B(n_461),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1344),
.B(n_508),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1386),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1323),
.A2(n_856),
.B(n_744),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1269),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1391),
.B(n_1232),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1257),
.A2(n_856),
.B(n_744),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1386),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1294),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1369),
.B(n_1322),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1360),
.B(n_508),
.Y(n_1472)
);

BUFx8_ASAP7_75t_L g1473 ( 
.A(n_1377),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1257),
.A2(n_856),
.B(n_745),
.Y(n_1474)
);

AOI221x1_ASAP7_75t_L g1475 ( 
.A1(n_1259),
.A2(n_833),
.B1(n_806),
.B2(n_802),
.C(n_800),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1260),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1259),
.A2(n_745),
.B(n_736),
.Y(n_1477)
);

BUFx10_ASAP7_75t_L g1478 ( 
.A(n_1372),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1323),
.A2(n_776),
.B(n_751),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1386),
.B(n_751),
.Y(n_1480)
);

BUFx3_ASAP7_75t_L g1481 ( 
.A(n_1262),
.Y(n_1481)
);

AOI21xp33_ASAP7_75t_L g1482 ( 
.A1(n_1231),
.A2(n_464),
.B(n_463),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1246),
.A2(n_1277),
.B(n_1331),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1322),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1240),
.B(n_776),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_SL g1486 ( 
.A(n_1386),
.B(n_464),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1388),
.B(n_406),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1246),
.A2(n_802),
.B(n_782),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1249),
.B(n_777),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1277),
.A2(n_782),
.B(n_777),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1255),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_SL g1492 ( 
.A1(n_1335),
.A2(n_667),
.B(n_662),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1383),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1289),
.B(n_408),
.Y(n_1494)
);

O2A1O1Ixp5_ASAP7_75t_L g1495 ( 
.A1(n_1225),
.A2(n_800),
.B(n_663),
.C(n_676),
.Y(n_1495)
);

AO31x2_ASAP7_75t_L g1496 ( 
.A1(n_1286),
.A2(n_663),
.A3(n_676),
.B(n_675),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1264),
.A2(n_716),
.B(n_653),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1331),
.A2(n_1343),
.B(n_1352),
.Y(n_1498)
);

AOI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1264),
.A2(n_664),
.B(n_676),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_SL g1500 ( 
.A1(n_1335),
.A2(n_653),
.B(n_675),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1263),
.A2(n_408),
.B(n_409),
.C(n_307),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1355),
.B(n_309),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1270),
.A2(n_663),
.B(n_675),
.Y(n_1503)
);

O2A1O1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1319),
.A2(n_667),
.B(n_664),
.C(n_662),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1291),
.A2(n_653),
.B(n_667),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1348),
.B(n_316),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1255),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1237),
.A2(n_430),
.B(n_319),
.C(n_323),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1378),
.B(n_662),
.Y(n_1509)
);

NOR2xp67_ASAP7_75t_L g1510 ( 
.A(n_1276),
.B(n_93),
.Y(n_1510)
);

AO32x2_ASAP7_75t_L g1511 ( 
.A1(n_1371),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1295),
.A2(n_664),
.B(n_659),
.Y(n_1512)
);

AO31x2_ASAP7_75t_L g1513 ( 
.A1(n_1292),
.A2(n_651),
.A3(n_659),
.B(n_605),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1339),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_SL g1515 ( 
.A1(n_1227),
.A2(n_164),
.B(n_236),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1266),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1251),
.B(n_317),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1270),
.A2(n_602),
.B(n_605),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1296),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1284),
.A2(n_602),
.B(n_605),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1368),
.A2(n_437),
.B(n_325),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1297),
.B(n_687),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_L g1523 ( 
.A(n_1356),
.B(n_428),
.C(n_327),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1284),
.A2(n_602),
.B(n_324),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1313),
.B(n_651),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1287),
.B(n_651),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1322),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1250),
.A2(n_659),
.B(n_651),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1275),
.A2(n_1376),
.B(n_1316),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1343),
.A2(n_602),
.B(n_600),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1352),
.A2(n_600),
.B(n_597),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1306),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1345),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1275),
.A2(n_1279),
.B(n_1288),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1301),
.A2(n_438),
.B1(n_354),
.B2(n_358),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1382),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1321),
.B(n_651),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1304),
.A2(n_1281),
.B(n_1351),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1273),
.A2(n_600),
.B(n_597),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1308),
.B(n_328),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1359),
.A2(n_600),
.B(n_597),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1266),
.B(n_597),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1359),
.A2(n_600),
.B(n_659),
.Y(n_1543)
);

INVx6_ASAP7_75t_L g1544 ( 
.A(n_1311),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1354),
.B(n_363),
.Y(n_1545)
);

NOR2xp67_ASAP7_75t_L g1546 ( 
.A(n_1293),
.B(n_95),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1380),
.B(n_367),
.Y(n_1547)
);

AO31x2_ASAP7_75t_L g1548 ( 
.A1(n_1385),
.A2(n_659),
.A3(n_651),
.B(n_8),
.Y(n_1548)
);

O2A1O1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1242),
.A2(n_373),
.B(n_416),
.C(n_419),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1327),
.B(n_659),
.Y(n_1550)
);

A2O1A1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1302),
.A2(n_446),
.B(n_427),
.C(n_439),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1279),
.A2(n_659),
.B(n_600),
.Y(n_1552)
);

OAI22x1_ASAP7_75t_L g1553 ( 
.A1(n_1364),
.A2(n_420),
.B1(n_443),
.B2(n_445),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1250),
.A2(n_643),
.B(n_610),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1266),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1298),
.B(n_4),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1282),
.B(n_7),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1330),
.B(n_607),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1317),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1310),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1337),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1325),
.A2(n_643),
.B(n_610),
.C(n_607),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1250),
.B(n_607),
.Y(n_1563)
);

INVx3_ASAP7_75t_SL g1564 ( 
.A(n_1317),
.Y(n_1564)
);

AOI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1353),
.A2(n_643),
.B(n_610),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1340),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1342),
.A2(n_117),
.B(n_234),
.Y(n_1567)
);

NOR4xp25_ASAP7_75t_L g1568 ( 
.A(n_1361),
.B(n_1387),
.C(n_1370),
.D(n_1366),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1288),
.A2(n_643),
.B(n_610),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1317),
.B(n_607),
.Y(n_1570)
);

BUFx4_ASAP7_75t_SL g1571 ( 
.A(n_1328),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1349),
.A2(n_112),
.B(n_226),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1456),
.Y(n_1573)
);

OA21x2_ASAP7_75t_L g1574 ( 
.A1(n_1534),
.A2(n_1365),
.B(n_1288),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1539),
.A2(n_1245),
.B(n_1226),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1534),
.A2(n_1375),
.B(n_1228),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1487),
.A2(n_1256),
.B1(n_1326),
.B2(n_1336),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1467),
.B(n_1226),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1432),
.A2(n_1245),
.B(n_1280),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1459),
.A2(n_643),
.B(n_610),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1410),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1467),
.B(n_1280),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1405),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1486),
.A2(n_1406),
.B1(n_1523),
.B2(n_1535),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1419),
.B(n_1389),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1422),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1422),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1434),
.A2(n_1283),
.B(n_1336),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1401),
.A2(n_1283),
.B(n_1336),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1436),
.A2(n_1389),
.B1(n_643),
.B2(n_610),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1490),
.A2(n_1389),
.B(n_607),
.Y(n_1591)
);

AOI21xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1421),
.A2(n_9),
.B(n_14),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1429),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1529),
.A2(n_15),
.B(n_17),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1479),
.A2(n_607),
.B(n_98),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1399),
.B(n_17),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1399),
.B(n_21),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1443),
.A2(n_23),
.B1(n_25),
.B2(n_33),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1422),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1499),
.A2(n_133),
.B(n_220),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1412),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1419),
.A2(n_128),
.B(n_219),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1420),
.A2(n_122),
.B(n_215),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1544),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1488),
.A2(n_222),
.B(n_200),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1464),
.Y(n_1606)
);

AO31x2_ASAP7_75t_L g1607 ( 
.A1(n_1403),
.A2(n_39),
.A3(n_40),
.B(n_41),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1449),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1445),
.A2(n_198),
.B(n_194),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1465),
.A2(n_191),
.B(n_188),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1477),
.A2(n_187),
.B(n_182),
.Y(n_1611)
);

BUFx12f_ASAP7_75t_L g1612 ( 
.A(n_1396),
.Y(n_1612)
);

NAND2x1p5_ASAP7_75t_L g1613 ( 
.A(n_1464),
.B(n_177),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1544),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1452),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1466),
.Y(n_1616)
);

CKINVDCx20_ASAP7_75t_R g1617 ( 
.A(n_1473),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1519),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1533),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1557),
.A2(n_40),
.B1(n_42),
.B2(n_47),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_SL g1621 ( 
.A1(n_1515),
.A2(n_42),
.B(n_49),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1398),
.A2(n_1438),
.B(n_1435),
.C(n_1409),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1477),
.A2(n_172),
.B(n_171),
.Y(n_1623)
);

AO31x2_ASAP7_75t_L g1624 ( 
.A1(n_1446),
.A2(n_1440),
.A3(n_1420),
.B(n_1475),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1447),
.A2(n_170),
.B(n_168),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_SL g1626 ( 
.A1(n_1400),
.A2(n_49),
.B(n_50),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1497),
.A2(n_167),
.B(n_163),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1556),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1476),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1450),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1450),
.Y(n_1631)
);

NOR2xp67_ASAP7_75t_L g1632 ( 
.A(n_1470),
.B(n_157),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1523),
.A2(n_52),
.B1(n_55),
.B2(n_58),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1497),
.A2(n_153),
.B(n_151),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1451),
.B(n_55),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1398),
.B(n_59),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1483),
.A2(n_150),
.B(n_145),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1473),
.Y(n_1638)
);

CKINVDCx11_ASAP7_75t_R g1639 ( 
.A(n_1478),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_1536),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1453),
.A2(n_142),
.B(n_141),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1450),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1482),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.C(n_64),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1566),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1393),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1409),
.A2(n_63),
.B(n_65),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1492),
.Y(n_1647)
);

O2A1O1Ixp5_ASAP7_75t_L g1648 ( 
.A1(n_1417),
.A2(n_66),
.B(n_67),
.C(n_69),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1417),
.A2(n_66),
.B(n_67),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1552),
.A2(n_71),
.B(n_75),
.Y(n_1650)
);

NAND2x1p5_ASAP7_75t_L g1651 ( 
.A(n_1469),
.B(n_82),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1531),
.A2(n_78),
.B(n_81),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1415),
.A2(n_78),
.B(n_81),
.Y(n_1653)
);

OAI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1486),
.A2(n_1424),
.B1(n_1404),
.B2(n_1484),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1425),
.A2(n_1414),
.B(n_1530),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1500),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1418),
.A2(n_1426),
.B(n_1474),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1468),
.A2(n_1474),
.B(n_1430),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1480),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1413),
.B(n_1439),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1427),
.B(n_1424),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1397),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1468),
.A2(n_1423),
.B(n_1569),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1503),
.A2(n_1435),
.B(n_1569),
.Y(n_1664)
);

A2O1A1Ixp33_ASAP7_75t_L g1665 ( 
.A1(n_1438),
.A2(n_1482),
.B(n_1441),
.C(n_1407),
.Y(n_1665)
);

CKINVDCx6p67_ASAP7_75t_R g1666 ( 
.A(n_1564),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1428),
.B(n_1471),
.Y(n_1667)
);

OAI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1568),
.A2(n_1501),
.B(n_1461),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1462),
.A2(n_1506),
.B1(n_1545),
.B2(n_1547),
.Y(n_1669)
);

BUFx8_ASAP7_75t_L g1670 ( 
.A(n_1395),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1448),
.B(n_1463),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_SL g1672 ( 
.A(n_1433),
.B(n_1454),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1493),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1517),
.A2(n_1471),
.B1(n_1527),
.B2(n_1560),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1413),
.B(n_1407),
.Y(n_1675)
);

O2A1O1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1560),
.A2(n_1508),
.B(n_1551),
.C(n_1494),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1561),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1472),
.B(n_1540),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1444),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1532),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1505),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1568),
.A2(n_1460),
.B(n_1439),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1543),
.A2(n_1541),
.B(n_1498),
.Y(n_1683)
);

OA21x2_ASAP7_75t_L g1684 ( 
.A1(n_1392),
.A2(n_1503),
.B(n_1518),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1411),
.A2(n_1416),
.B(n_1458),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1509),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1512),
.A2(n_1572),
.B(n_1567),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1437),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1395),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1511),
.B(n_1509),
.Y(n_1690)
);

INVx6_ASAP7_75t_L g1691 ( 
.A(n_1395),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1505),
.Y(n_1692)
);

NAND2x1p5_ASAP7_75t_L g1693 ( 
.A(n_1514),
.B(n_1402),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1518),
.A2(n_1562),
.B(n_1538),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1520),
.A2(n_1524),
.B(n_1489),
.Y(n_1695)
);

NOR2xp67_ASAP7_75t_SL g1696 ( 
.A(n_1402),
.B(n_1481),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1526),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1565),
.A2(n_1554),
.B(n_1495),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1478),
.B(n_1454),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1522),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1522),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1460),
.A2(n_1553),
.B1(n_1502),
.B2(n_1521),
.Y(n_1702)
);

OAI21x1_ASAP7_75t_L g1703 ( 
.A1(n_1563),
.A2(n_1520),
.B(n_1525),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1549),
.B(n_1521),
.C(n_1546),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1402),
.Y(n_1705)
);

AO21x2_ASAP7_75t_L g1706 ( 
.A1(n_1524),
.A2(n_1489),
.B(n_1485),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_SL g1707 ( 
.A(n_1528),
.B(n_1514),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1555),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1526),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1457),
.A2(n_1485),
.B(n_1431),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1442),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1525),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1457),
.A2(n_1433),
.B(n_1504),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1558),
.Y(n_1714)
);

AND2x6_ASAP7_75t_L g1715 ( 
.A(n_1428),
.B(n_1455),
.Y(n_1715)
);

OAI21x1_ASAP7_75t_L g1716 ( 
.A1(n_1442),
.A2(n_1537),
.B(n_1550),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1537),
.A2(n_1550),
.B(n_1558),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1548),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1408),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1548),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1510),
.B(n_1559),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1480),
.A2(n_1455),
.B1(n_1516),
.B2(n_1570),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1516),
.A2(n_1570),
.B1(n_1408),
.B2(n_1491),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1542),
.A2(n_1496),
.B(n_1513),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1496),
.Y(n_1725)
);

OAI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1408),
.A2(n_1491),
.B1(n_1507),
.B2(n_1571),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1511),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1496),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1542),
.A2(n_1513),
.B(n_1394),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1491),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1507),
.A2(n_1511),
.B1(n_1394),
.B2(n_1513),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1507),
.A2(n_1247),
.B(n_1398),
.C(n_1145),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1406),
.B(n_1145),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1422),
.Y(n_1734)
);

AO21x2_ASAP7_75t_L g1735 ( 
.A1(n_1534),
.A2(n_1420),
.B(n_1419),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1410),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1395),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1422),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1432),
.Y(n_1739)
);

OAI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1432),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1456),
.Y(n_1741)
);

OA21x2_ASAP7_75t_L g1742 ( 
.A1(n_1534),
.A2(n_1459),
.B(n_1483),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1456),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1534),
.A2(n_1459),
.B(n_1483),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1456),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1436),
.A2(n_1145),
.B1(n_1004),
.B2(n_803),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1487),
.A2(n_1145),
.B1(n_905),
.B2(n_1557),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1432),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1467),
.B(n_1413),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1456),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1436),
.A2(n_1145),
.B1(n_1004),
.B2(n_803),
.Y(n_1751)
);

OA21x2_ASAP7_75t_L g1752 ( 
.A1(n_1534),
.A2(n_1459),
.B(n_1483),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1410),
.Y(n_1753)
);

OA21x2_ASAP7_75t_L g1754 ( 
.A1(n_1534),
.A2(n_1459),
.B(n_1483),
.Y(n_1754)
);

NAND2x1_ASAP7_75t_L g1755 ( 
.A(n_1464),
.B(n_1469),
.Y(n_1755)
);

BUFx8_ASAP7_75t_L g1756 ( 
.A(n_1395),
.Y(n_1756)
);

AND2x2_ASAP7_75t_SL g1757 ( 
.A(n_1436),
.B(n_983),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1406),
.B(n_1145),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1544),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1464),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1422),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1422),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1432),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1534),
.A2(n_1459),
.B(n_1483),
.Y(n_1764)
);

OAI21x1_ASAP7_75t_L g1765 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1432),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1432),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1422),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1539),
.A2(n_1434),
.B(n_1432),
.Y(n_1768)
);

AO21x2_ASAP7_75t_L g1769 ( 
.A1(n_1534),
.A2(n_1420),
.B(n_1419),
.Y(n_1769)
);

AO31x2_ASAP7_75t_L g1770 ( 
.A1(n_1534),
.A2(n_1358),
.A3(n_1403),
.B(n_1459),
.Y(n_1770)
);

AO21x2_ASAP7_75t_L g1771 ( 
.A1(n_1534),
.A2(n_1420),
.B(n_1419),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1487),
.A2(n_1145),
.B1(n_1131),
.B2(n_770),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1622),
.A2(n_1757),
.B(n_1636),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1667),
.B(n_1661),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1601),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1601),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1622),
.A2(n_1757),
.B(n_1636),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1673),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1594),
.A2(n_1676),
.B(n_1732),
.Y(n_1779)
);

AOI21x1_ASAP7_75t_SL g1780 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1690),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1667),
.B(n_1679),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1660),
.B(n_1749),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1667),
.B(n_1582),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1747),
.A2(n_1620),
.B1(n_1628),
.B2(n_1633),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1639),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1582),
.B(n_1671),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1732),
.A2(n_1643),
.B1(n_1772),
.B2(n_1665),
.Y(n_1787)
);

O2A1O1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1665),
.A2(n_1592),
.B(n_1668),
.C(n_1598),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1660),
.B(n_1699),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1678),
.B(n_1674),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1749),
.A2(n_1646),
.B1(n_1702),
.B2(n_1733),
.Y(n_1791)
);

CKINVDCx12_ASAP7_75t_R g1792 ( 
.A(n_1578),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1593),
.B(n_1758),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1581),
.B(n_1753),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_SL g1795 ( 
.A1(n_1746),
.A2(n_1751),
.B(n_1590),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1593),
.B(n_1581),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1578),
.B(n_1690),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1753),
.B(n_1736),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1635),
.B(n_1573),
.Y(n_1799)
);

OA21x2_ASAP7_75t_L g1800 ( 
.A1(n_1663),
.A2(n_1685),
.B(n_1657),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1669),
.A2(n_1616),
.B1(n_1608),
.B2(n_1615),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1640),
.B(n_1645),
.Y(n_1802)
);

INVx5_ASAP7_75t_L g1803 ( 
.A(n_1585),
.Y(n_1803)
);

O2A1O1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1584),
.A2(n_1648),
.B(n_1654),
.C(n_1626),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1741),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1629),
.B(n_1680),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1664),
.A2(n_1684),
.B(n_1710),
.Y(n_1807)
);

AOI21x1_ASAP7_75t_SL g1808 ( 
.A1(n_1721),
.A2(n_1688),
.B(n_1649),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1743),
.B(n_1745),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1750),
.B(n_1662),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_L g1811 ( 
.A(n_1614),
.B(n_1759),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1708),
.B(n_1614),
.Y(n_1812)
);

O2A1O1Ixp5_ASAP7_75t_L g1813 ( 
.A1(n_1682),
.A2(n_1603),
.B(n_1713),
.C(n_1704),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1613),
.A2(n_1649),
.B(n_1722),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1686),
.B(n_1677),
.Y(n_1815)
);

NOR2xp67_ASAP7_75t_L g1816 ( 
.A(n_1759),
.B(n_1583),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1618),
.A2(n_1577),
.B1(n_1619),
.B2(n_1727),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1664),
.A2(n_1684),
.B(n_1585),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1726),
.A2(n_1644),
.B1(n_1651),
.B2(n_1701),
.Y(n_1819)
);

BUFx8_ASAP7_75t_L g1820 ( 
.A(n_1612),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1718),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1708),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1585),
.A2(n_1706),
.B(n_1695),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1613),
.A2(n_1649),
.B(n_1651),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1719),
.B(n_1604),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1585),
.A2(n_1706),
.B(n_1695),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1700),
.A2(n_1712),
.B1(n_1640),
.B2(n_1666),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1693),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1714),
.B(n_1697),
.Y(n_1829)
);

BUFx12f_ASAP7_75t_L g1830 ( 
.A(n_1638),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1693),
.Y(n_1831)
);

OA21x2_ASAP7_75t_L g1832 ( 
.A1(n_1663),
.A2(n_1685),
.B(n_1657),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1604),
.B(n_1706),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1697),
.B(n_1709),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1715),
.B(n_1606),
.Y(n_1835)
);

O2A1O1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1621),
.A2(n_1647),
.B(n_1656),
.C(n_1602),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1730),
.B(n_1689),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1720),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1730),
.B(n_1689),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_R g1840 ( 
.A(n_1583),
.B(n_1638),
.Y(n_1840)
);

O2A1O1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1647),
.A2(n_1656),
.B(n_1602),
.C(n_1731),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1709),
.B(n_1672),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1666),
.A2(n_1632),
.B1(n_1695),
.B2(n_1691),
.Y(n_1843)
);

NOR2xp67_ASAP7_75t_L g1844 ( 
.A(n_1612),
.B(n_1606),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1691),
.Y(n_1845)
);

OA21x2_ASAP7_75t_L g1846 ( 
.A1(n_1658),
.A2(n_1740),
.B(n_1739),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1711),
.B(n_1586),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1711),
.B(n_1586),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1705),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1639),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1705),
.B(n_1737),
.Y(n_1851)
);

AOI21x1_ASAP7_75t_SL g1852 ( 
.A1(n_1607),
.A2(n_1602),
.B(n_1707),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1715),
.B(n_1606),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1691),
.A2(n_1617),
.B1(n_1737),
.B2(n_1580),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1587),
.B(n_1599),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1691),
.A2(n_1617),
.B1(n_1737),
.B2(n_1580),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1715),
.B(n_1760),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1715),
.B(n_1607),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1641),
.A2(n_1611),
.B(n_1623),
.C(n_1650),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1587),
.B(n_1599),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1580),
.A2(n_1738),
.B1(n_1767),
.B2(n_1734),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1723),
.Y(n_1862)
);

O2A1O1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1760),
.A2(n_1755),
.B(n_1767),
.C(n_1734),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1715),
.B(n_1760),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1761),
.Y(n_1865)
);

CKINVDCx6p67_ASAP7_75t_R g1866 ( 
.A(n_1715),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1607),
.B(n_1762),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1670),
.Y(n_1868)
);

NOR2x1_ASAP7_75t_SL g1869 ( 
.A(n_1576),
.B(n_1762),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_SL g1870 ( 
.A1(n_1694),
.A2(n_1696),
.B(n_1670),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1607),
.B(n_1653),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1694),
.A2(n_1725),
.B1(n_1728),
.B2(n_1659),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1607),
.B(n_1653),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1770),
.B(n_1576),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1694),
.A2(n_1728),
.B1(n_1725),
.B2(n_1659),
.Y(n_1875)
);

O2A1O1Ixp5_ASAP7_75t_L g1876 ( 
.A1(n_1630),
.A2(n_1631),
.B(n_1642),
.C(n_1681),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1681),
.A2(n_1692),
.B1(n_1574),
.B2(n_1764),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1692),
.Y(n_1878)
);

O2A1O1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1576),
.A2(n_1771),
.B(n_1769),
.C(n_1735),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1579),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1652),
.B(n_1623),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1670),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1574),
.A2(n_1744),
.B1(n_1742),
.B2(n_1764),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1579),
.Y(n_1885)
);

A2O1A1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1611),
.A2(n_1627),
.B(n_1634),
.C(n_1637),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1588),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1717),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1574),
.A2(n_1744),
.B1(n_1742),
.B2(n_1764),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1717),
.Y(n_1890)
);

AND2x6_ASAP7_75t_L g1891 ( 
.A(n_1756),
.B(n_1637),
.Y(n_1891)
);

O2A1O1Ixp33_ASAP7_75t_L g1892 ( 
.A1(n_1771),
.A2(n_1754),
.B(n_1752),
.C(n_1744),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1770),
.B(n_1624),
.Y(n_1893)
);

O2A1O1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1752),
.A2(n_1754),
.B(n_1756),
.C(n_1624),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1652),
.B(n_1589),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1589),
.B(n_1729),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1770),
.B(n_1624),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1752),
.A2(n_1754),
.B(n_1687),
.Y(n_1898)
);

OA21x2_ASAP7_75t_L g1899 ( 
.A1(n_1739),
.A2(n_1763),
.B(n_1765),
.Y(n_1899)
);

OA22x2_ASAP7_75t_L g1900 ( 
.A1(n_1609),
.A2(n_1625),
.B1(n_1729),
.B2(n_1703),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1770),
.B(n_1624),
.Y(n_1901)
);

OA21x2_ASAP7_75t_L g1902 ( 
.A1(n_1740),
.A2(n_1768),
.B(n_1766),
.Y(n_1902)
);

NAND4xp25_ASAP7_75t_L g1903 ( 
.A(n_1756),
.B(n_1625),
.C(n_1609),
.D(n_1716),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1687),
.A2(n_1703),
.B(n_1766),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1716),
.Y(n_1905)
);

OAI22xp5_ASAP7_75t_L g1906 ( 
.A1(n_1724),
.A2(n_1600),
.B1(n_1605),
.B2(n_1698),
.Y(n_1906)
);

O2A1O1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1600),
.A2(n_1605),
.B(n_1610),
.C(n_1698),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1748),
.A2(n_1768),
.B(n_1655),
.Y(n_1908)
);

NOR2xp67_ASAP7_75t_L g1909 ( 
.A(n_1575),
.B(n_1610),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1655),
.B(n_1748),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1683),
.B(n_1591),
.Y(n_1911)
);

O2A1O1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1595),
.A2(n_1594),
.B(n_1772),
.C(n_1636),
.Y(n_1912)
);

AOI21x1_ASAP7_75t_SL g1913 ( 
.A1(n_1595),
.A2(n_1683),
.B(n_1591),
.Y(n_1913)
);

O2A1O1Ixp33_ASAP7_75t_L g1914 ( 
.A1(n_1594),
.A2(n_1772),
.B(n_1636),
.C(n_1487),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1667),
.B(n_1661),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1747),
.A2(n_1145),
.B1(n_1636),
.B2(n_1622),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1645),
.Y(n_1917)
);

AOI21x1_ASAP7_75t_SL g1918 ( 
.A1(n_1596),
.A2(n_1547),
.B(n_1557),
.Y(n_1918)
);

OAI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1747),
.A2(n_1145),
.B1(n_1636),
.B2(n_1622),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1622),
.A2(n_1398),
.B(n_1314),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1667),
.B(n_1661),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1622),
.A2(n_1398),
.B(n_1314),
.Y(n_1922)
);

AND2x4_ASAP7_75t_L g1923 ( 
.A(n_1667),
.B(n_1708),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1601),
.Y(n_1924)
);

AOI21x1_ASAP7_75t_SL g1925 ( 
.A1(n_1596),
.A2(n_1547),
.B(n_1557),
.Y(n_1925)
);

O2A1O1Ixp5_ASAP7_75t_L g1926 ( 
.A1(n_1594),
.A2(n_1636),
.B(n_1646),
.C(n_1668),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1660),
.B(n_1749),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1667),
.B(n_1708),
.Y(n_1928)
);

OA21x2_ASAP7_75t_L g1929 ( 
.A1(n_1663),
.A2(n_1685),
.B(n_1534),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1622),
.A2(n_1398),
.B(n_1314),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1747),
.A2(n_1145),
.B1(n_1636),
.B2(n_1622),
.Y(n_1931)
);

AND2x2_ASAP7_75t_SL g1932 ( 
.A(n_1757),
.B(n_1747),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1661),
.B(n_1675),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1661),
.B(n_1679),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1667),
.B(n_1661),
.Y(n_1935)
);

AOI21x1_ASAP7_75t_SL g1936 ( 
.A1(n_1596),
.A2(n_1547),
.B(n_1557),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1661),
.B(n_1679),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1661),
.B(n_1675),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1594),
.A2(n_1398),
.B(n_1145),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1601),
.Y(n_1940)
);

OA21x2_ASAP7_75t_L g1941 ( 
.A1(n_1663),
.A2(n_1685),
.B(n_1534),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1601),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1660),
.B(n_1749),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1789),
.B(n_1933),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1887),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1775),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1797),
.B(n_1782),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1821),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1838),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1797),
.B(n_1786),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1858),
.B(n_1943),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1849),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1833),
.B(n_1847),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1792),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1916),
.A2(n_1919),
.B1(n_1931),
.B2(n_1784),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1822),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1914),
.A2(n_1813),
.B(n_1926),
.Y(n_1957)
);

HB1xp67_ASAP7_75t_L g1958 ( 
.A(n_1778),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1782),
.B(n_1927),
.Y(n_1959)
);

OR2x6_ASAP7_75t_L g1960 ( 
.A(n_1814),
.B(n_1920),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1943),
.B(n_1927),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1913),
.A2(n_1908),
.B(n_1904),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1796),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1923),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1938),
.B(n_1934),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1871),
.B(n_1873),
.Y(n_1966)
);

OA21x2_ASAP7_75t_L g1967 ( 
.A1(n_1898),
.A2(n_1818),
.B(n_1807),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1937),
.B(n_1774),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1887),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1783),
.B(n_1915),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1848),
.B(n_1867),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1900),
.A2(n_1907),
.B(n_1906),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1776),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1921),
.B(n_1935),
.Y(n_1974)
);

OR2x6_ASAP7_75t_L g1975 ( 
.A(n_1922),
.B(n_1930),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1939),
.A2(n_1779),
.B(n_1916),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1803),
.B(n_1835),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1878),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1794),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1924),
.Y(n_1980)
);

INVx2_ASAP7_75t_SL g1981 ( 
.A(n_1940),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1942),
.Y(n_1982)
);

AO21x2_ASAP7_75t_L g1983 ( 
.A1(n_1886),
.A2(n_1826),
.B(n_1823),
.Y(n_1983)
);

INVx3_ASAP7_75t_L g1984 ( 
.A(n_1853),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1865),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1781),
.B(n_1773),
.Y(n_1986)
);

OAI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1919),
.A2(n_1931),
.B(n_1788),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1777),
.B(n_1888),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1890),
.B(n_1805),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1849),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1905),
.Y(n_1991)
);

OR2x6_ASAP7_75t_L g1992 ( 
.A(n_1824),
.B(n_1870),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1876),
.Y(n_1993)
);

AO21x2_ASAP7_75t_L g1994 ( 
.A1(n_1859),
.A2(n_1909),
.B(n_1889),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1874),
.B(n_1901),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1799),
.B(n_1809),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1855),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1812),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1893),
.B(n_1897),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1860),
.Y(n_2000)
);

AOI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1843),
.A2(n_1791),
.B(n_1787),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1790),
.B(n_1798),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1860),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1842),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1842),
.Y(n_2005)
);

BUFx2_ASAP7_75t_L g2006 ( 
.A(n_1923),
.Y(n_2006)
);

BUFx2_ASAP7_75t_L g2007 ( 
.A(n_1928),
.Y(n_2007)
);

AO21x2_ASAP7_75t_L g2008 ( 
.A1(n_1884),
.A2(n_1889),
.B(n_1879),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1810),
.B(n_1895),
.Y(n_2009)
);

NAND2x1_ASAP7_75t_L g2010 ( 
.A(n_1853),
.B(n_1857),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1793),
.B(n_1806),
.Y(n_2011)
);

OR2x2_ASAP7_75t_L g2012 ( 
.A(n_1893),
.B(n_1897),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1791),
.B(n_1815),
.Y(n_2013)
);

OAI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1912),
.A2(n_1787),
.B(n_1804),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1877),
.B(n_1881),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1834),
.Y(n_2016)
);

INVx4_ASAP7_75t_L g2017 ( 
.A(n_1866),
.Y(n_2017)
);

INVx2_ASAP7_75t_SL g2018 ( 
.A(n_1812),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1834),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1896),
.B(n_1869),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1801),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1877),
.B(n_1885),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1829),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1872),
.B(n_1875),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1872),
.B(n_1875),
.Y(n_2025)
);

OR2x6_ASAP7_75t_L g2026 ( 
.A(n_1841),
.B(n_1836),
.Y(n_2026)
);

AO21x2_ASAP7_75t_L g2027 ( 
.A1(n_1906),
.A2(n_1892),
.B(n_1911),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1883),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1928),
.Y(n_2029)
);

NAND2x1_ASAP7_75t_L g2030 ( 
.A(n_1857),
.B(n_1864),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1829),
.Y(n_2031)
);

BUFx3_ASAP7_75t_L g2032 ( 
.A(n_1917),
.Y(n_2032)
);

OAI21x1_ASAP7_75t_L g2033 ( 
.A1(n_1900),
.A2(n_1852),
.B(n_1861),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1932),
.B(n_1941),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1801),
.B(n_1827),
.Y(n_2035)
);

OAI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1784),
.A2(n_1795),
.B(n_1827),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1817),
.B(n_1862),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1817),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1819),
.Y(n_2039)
);

AOI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1843),
.A2(n_1819),
.B(n_1844),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1863),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1840),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1861),
.Y(n_2043)
);

OA21x2_ASAP7_75t_L g2044 ( 
.A1(n_1882),
.A2(n_1880),
.B(n_1854),
.Y(n_2044)
);

INVx1_ASAP7_75t_SL g2045 ( 
.A(n_1825),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1831),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1846),
.Y(n_2047)
);

OA21x2_ASAP7_75t_L g2048 ( 
.A1(n_1854),
.A2(n_1856),
.B(n_1903),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1894),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_1929),
.B(n_1941),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1948),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_2005),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1991),
.Y(n_2053)
);

AND2x4_ASAP7_75t_L g2054 ( 
.A(n_2020),
.B(n_1910),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1949),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_2004),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2047),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_2020),
.B(n_1864),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_1953),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2047),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1945),
.B(n_1851),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1951),
.B(n_1966),
.Y(n_2062)
);

OAI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1955),
.A2(n_2036),
.B1(n_1976),
.B2(n_1987),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1958),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2009),
.B(n_1961),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1989),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2009),
.B(n_1856),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2050),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1946),
.Y(n_2069)
);

OR2x2_ASAP7_75t_L g2070 ( 
.A(n_1995),
.B(n_1800),
.Y(n_2070)
);

AO21x2_ASAP7_75t_L g2071 ( 
.A1(n_1962),
.A2(n_1957),
.B(n_2008),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1959),
.B(n_1802),
.Y(n_2072)
);

BUFx6f_ASAP7_75t_L g2073 ( 
.A(n_1992),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2050),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_1995),
.B(n_1832),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1946),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1950),
.B(n_1800),
.Y(n_2077)
);

A2O1A1Ixp33_ASAP7_75t_L g2078 ( 
.A1(n_2014),
.A2(n_1816),
.B(n_1811),
.C(n_1883),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1971),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1969),
.B(n_1891),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2011),
.B(n_1828),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1965),
.B(n_1839),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1950),
.B(n_1837),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1971),
.Y(n_2084)
);

NAND2x1_ASAP7_75t_L g2085 ( 
.A(n_1992),
.B(n_1891),
.Y(n_2085)
);

OAI33xp33_ASAP7_75t_L g2086 ( 
.A1(n_2035),
.A2(n_1785),
.A3(n_1850),
.B1(n_1780),
.B2(n_1936),
.B3(n_1925),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_1947),
.B(n_1902),
.Y(n_2087)
);

OR2x2_ASAP7_75t_L g2088 ( 
.A(n_2015),
.B(n_1902),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2015),
.B(n_1899),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1978),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1988),
.B(n_1845),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2034),
.B(n_1986),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1960),
.A2(n_1868),
.B1(n_1830),
.B2(n_1918),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1975),
.A2(n_1820),
.B1(n_1891),
.B2(n_1808),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2022),
.B(n_2043),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_1963),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1984),
.B(n_1820),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_1999),
.B(n_2012),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1944),
.B(n_2013),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2034),
.B(n_1986),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2053),
.Y(n_2101)
);

NOR3xp33_ASAP7_75t_L g2102 ( 
.A(n_2063),
.B(n_2001),
.C(n_2040),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2057),
.Y(n_2103)
);

NAND4xp25_ASAP7_75t_L g2104 ( 
.A(n_2078),
.B(n_2037),
.C(n_2049),
.D(n_2041),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2092),
.B(n_2044),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_2086),
.A2(n_1975),
.B1(n_1960),
.B2(n_2039),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_2094),
.A2(n_1960),
.B1(n_1975),
.B2(n_2021),
.Y(n_2107)
);

AND2x2_ASAP7_75t_SL g2108 ( 
.A(n_2073),
.B(n_2048),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2057),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2057),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2092),
.B(n_2100),
.Y(n_2111)
);

NAND3xp33_ASAP7_75t_L g2112 ( 
.A(n_2093),
.B(n_2026),
.C(n_2038),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2100),
.B(n_2044),
.Y(n_2113)
);

INVxp67_ASAP7_75t_L g2114 ( 
.A(n_2096),
.Y(n_2114)
);

AOI221xp5_ASAP7_75t_L g2115 ( 
.A1(n_2064),
.A2(n_2002),
.B1(n_2046),
.B2(n_1963),
.C(n_1956),
.Y(n_2115)
);

NOR3xp33_ASAP7_75t_SL g2116 ( 
.A(n_2099),
.B(n_2042),
.C(n_2031),
.Y(n_2116)
);

BUFx2_ASAP7_75t_L g2117 ( 
.A(n_2054),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2052),
.B(n_1979),
.Y(n_2118)
);

INVxp67_ASAP7_75t_SL g2119 ( 
.A(n_2059),
.Y(n_2119)
);

AOI31xp33_ASAP7_75t_L g2120 ( 
.A1(n_2097),
.A2(n_2042),
.A3(n_1954),
.B(n_2045),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2079),
.Y(n_2121)
);

AOI222xp33_ASAP7_75t_L g2122 ( 
.A1(n_2072),
.A2(n_1996),
.B1(n_1968),
.B2(n_2023),
.C1(n_2016),
.C2(n_2019),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_2097),
.A2(n_1975),
.B1(n_1960),
.B2(n_2026),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2054),
.B(n_2044),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2051),
.Y(n_2125)
);

NAND3xp33_ASAP7_75t_L g2126 ( 
.A(n_2056),
.B(n_2026),
.C(n_2048),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2054),
.B(n_1979),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2081),
.A2(n_1996),
.B1(n_2003),
.B2(n_2000),
.C(n_1997),
.Y(n_2128)
);

OAI211xp5_ASAP7_75t_SL g2129 ( 
.A1(n_2095),
.A2(n_2024),
.B(n_2025),
.C(n_2018),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_2051),
.A2(n_1970),
.B1(n_1974),
.B2(n_1982),
.C(n_1980),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2097),
.A2(n_2026),
.B1(n_1992),
.B2(n_2017),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2054),
.B(n_2062),
.Y(n_2132)
);

OAI33xp33_ASAP7_75t_L g2133 ( 
.A1(n_2095),
.A2(n_2012),
.A3(n_1999),
.B1(n_2024),
.B2(n_2025),
.B3(n_1973),
.Y(n_2133)
);

AO21x2_ASAP7_75t_L g2134 ( 
.A1(n_2071),
.A2(n_2008),
.B(n_1983),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2062),
.B(n_2048),
.Y(n_2135)
);

OAI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_2097),
.A2(n_1992),
.B1(n_2017),
.B2(n_2032),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2060),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2084),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2060),
.Y(n_2139)
);

NAND4xp25_ASAP7_75t_L g2140 ( 
.A(n_2082),
.B(n_2032),
.C(n_1993),
.D(n_2017),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2065),
.B(n_2033),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2098),
.B(n_1993),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_2058),
.B(n_2080),
.Y(n_2143)
);

OAI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_2085),
.A2(n_1972),
.B(n_2033),
.Y(n_2144)
);

AO21x2_ASAP7_75t_L g2145 ( 
.A1(n_2071),
.A2(n_2008),
.B(n_1983),
.Y(n_2145)
);

OAI211xp5_ASAP7_75t_SL g2146 ( 
.A1(n_2070),
.A2(n_2018),
.B(n_1984),
.C(n_1981),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2065),
.B(n_1984),
.Y(n_2147)
);

CKINVDCx16_ASAP7_75t_R g2148 ( 
.A(n_2061),
.Y(n_2148)
);

OAI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2073),
.A2(n_2085),
.B1(n_2030),
.B2(n_2010),
.Y(n_2149)
);

AND2x4_ASAP7_75t_L g2150 ( 
.A(n_2058),
.B(n_1977),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2060),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_2061),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2069),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2069),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2076),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2098),
.B(n_2027),
.Y(n_2156)
);

BUFx3_ASAP7_75t_L g2157 ( 
.A(n_2061),
.Y(n_2157)
);

AOI222xp33_ASAP7_75t_L g2158 ( 
.A1(n_2067),
.A2(n_1974),
.B1(n_1970),
.B2(n_2006),
.C1(n_1964),
.C2(n_2007),
.Y(n_2158)
);

AOI221xp5_ASAP7_75t_L g2159 ( 
.A1(n_2055),
.A2(n_1981),
.B1(n_2029),
.B2(n_1983),
.C(n_1998),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2076),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2090),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2055),
.Y(n_2162)
);

NAND3xp33_ASAP7_75t_SL g2163 ( 
.A(n_2067),
.B(n_1985),
.C(n_1994),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2066),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2153),
.Y(n_2165)
);

OA21x2_ASAP7_75t_L g2166 ( 
.A1(n_2144),
.A2(n_2126),
.B(n_2159),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2153),
.Y(n_2167)
);

INVx2_ASAP7_75t_SL g2168 ( 
.A(n_2143),
.Y(n_2168)
);

NOR2x1_ASAP7_75t_SL g2169 ( 
.A(n_2163),
.B(n_2073),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2154),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2154),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2155),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2155),
.Y(n_2173)
);

OR2x6_ASAP7_75t_L g2174 ( 
.A(n_2131),
.B(n_2073),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2160),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2160),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2103),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2103),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2117),
.B(n_2135),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2142),
.B(n_2087),
.Y(n_2180)
);

INVxp67_ASAP7_75t_L g2181 ( 
.A(n_2121),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2161),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2109),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2161),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2109),
.Y(n_2185)
);

OA21x2_ASAP7_75t_L g2186 ( 
.A1(n_2156),
.A2(n_1972),
.B(n_1962),
.Y(n_2186)
);

INVx1_ASAP7_75t_SL g2187 ( 
.A(n_2108),
.Y(n_2187)
);

CKINVDCx16_ASAP7_75t_R g2188 ( 
.A(n_2148),
.Y(n_2188)
);

INVx11_ASAP7_75t_L g2189 ( 
.A(n_2120),
.Y(n_2189)
);

BUFx2_ASAP7_75t_L g2190 ( 
.A(n_2143),
.Y(n_2190)
);

INVx1_ASAP7_75t_SL g2191 ( 
.A(n_2108),
.Y(n_2191)
);

OR2x6_ASAP7_75t_L g2192 ( 
.A(n_2136),
.B(n_2073),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2110),
.Y(n_2193)
);

INVx4_ASAP7_75t_L g2194 ( 
.A(n_2134),
.Y(n_2194)
);

NAND3xp33_ASAP7_75t_L g2195 ( 
.A(n_2102),
.B(n_2073),
.C(n_1967),
.Y(n_2195)
);

OR2x2_ASAP7_75t_L g2196 ( 
.A(n_2142),
.B(n_2156),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2138),
.Y(n_2197)
);

INVx5_ASAP7_75t_L g2198 ( 
.A(n_2124),
.Y(n_2198)
);

BUFx8_ASAP7_75t_L g2199 ( 
.A(n_2117),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2137),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2164),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2125),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2104),
.B(n_2058),
.Y(n_2203)
);

OA21x2_ASAP7_75t_L g2204 ( 
.A1(n_2124),
.A2(n_2068),
.B(n_2074),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2162),
.Y(n_2205)
);

HB1xp67_ASAP7_75t_L g2206 ( 
.A(n_2119),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_2139),
.A2(n_2088),
.B(n_2089),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_2149),
.B(n_2058),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2101),
.Y(n_2209)
);

INVx2_ASAP7_75t_SL g2210 ( 
.A(n_2143),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2135),
.B(n_2077),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2151),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2101),
.Y(n_2213)
);

INVx3_ASAP7_75t_L g2214 ( 
.A(n_2199),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2207),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2181),
.B(n_2122),
.Y(n_2216)
);

INVxp67_ASAP7_75t_SL g2217 ( 
.A(n_2199),
.Y(n_2217)
);

AOI221xp5_ASAP7_75t_L g2218 ( 
.A1(n_2195),
.A2(n_2133),
.B1(n_2128),
.B2(n_2115),
.C(n_2130),
.Y(n_2218)
);

INVx1_ASAP7_75t_SL g2219 ( 
.A(n_2188),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2197),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2188),
.B(n_2105),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2165),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2190),
.B(n_2105),
.Y(n_2223)
);

NOR2x1_ASAP7_75t_L g2224 ( 
.A(n_2195),
.B(n_2112),
.Y(n_2224)
);

AOI211x1_ASAP7_75t_L g2225 ( 
.A1(n_2208),
.A2(n_2140),
.B(n_2189),
.C(n_2179),
.Y(n_2225)
);

OAI31xp33_ASAP7_75t_L g2226 ( 
.A1(n_2187),
.A2(n_2107),
.A3(n_2129),
.B(n_2146),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2203),
.B(n_2111),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_2206),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2190),
.B(n_2113),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2201),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_SL g2231 ( 
.A1(n_2166),
.A2(n_2071),
.B1(n_2145),
.B2(n_2134),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2187),
.B(n_2111),
.Y(n_2232)
);

AOI22x1_ASAP7_75t_L g2233 ( 
.A1(n_2191),
.A2(n_2189),
.B1(n_2194),
.B2(n_2158),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2191),
.B(n_2113),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2166),
.Y(n_2235)
);

NAND2x1_ASAP7_75t_L g2236 ( 
.A(n_2192),
.B(n_2150),
.Y(n_2236)
);

OR2x2_ASAP7_75t_L g2237 ( 
.A(n_2196),
.B(n_2087),
.Y(n_2237)
);

OAI211xp5_ASAP7_75t_L g2238 ( 
.A1(n_2166),
.A2(n_2106),
.B(n_2194),
.C(n_2116),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2168),
.B(n_2132),
.Y(n_2239)
);

NAND3xp33_ASAP7_75t_L g2240 ( 
.A(n_2166),
.B(n_2123),
.C(n_2114),
.Y(n_2240)
);

NAND4xp25_ASAP7_75t_L g2241 ( 
.A(n_2194),
.B(n_2118),
.C(n_2141),
.D(n_2091),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2165),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2167),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2207),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_2196),
.B(n_2070),
.Y(n_2245)
);

NOR2xp67_ASAP7_75t_L g2246 ( 
.A(n_2198),
.B(n_2150),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2168),
.B(n_2132),
.Y(n_2247)
);

NAND2x1p5_ASAP7_75t_L g2248 ( 
.A(n_2194),
.B(n_2080),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2210),
.B(n_2141),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2167),
.Y(n_2250)
);

OAI222xp33_ASAP7_75t_L g2251 ( 
.A1(n_2192),
.A2(n_2174),
.B1(n_2210),
.B2(n_2198),
.C1(n_2179),
.C2(n_2201),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2198),
.B(n_2150),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2170),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2170),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2180),
.B(n_2075),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2171),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2198),
.B(n_2152),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2198),
.B(n_2152),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2171),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2198),
.B(n_2157),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2198),
.B(n_2157),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_L g2262 ( 
.A1(n_2199),
.A2(n_2145),
.B1(n_2134),
.B2(n_2080),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2172),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2202),
.B(n_2147),
.Y(n_2264)
);

OR2x2_ASAP7_75t_L g2265 ( 
.A(n_2180),
.B(n_2075),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2223),
.Y(n_2266)
);

INVx1_ASAP7_75t_SL g2267 ( 
.A(n_2219),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2223),
.Y(n_2268)
);

OAI322xp33_ASAP7_75t_L g2269 ( 
.A1(n_2235),
.A2(n_2205),
.A3(n_2202),
.B1(n_2173),
.B2(n_2175),
.C1(n_2184),
.C2(n_2172),
.Y(n_2269)
);

OAI21xp33_ASAP7_75t_L g2270 ( 
.A1(n_2224),
.A2(n_2174),
.B(n_2192),
.Y(n_2270)
);

INVx1_ASAP7_75t_SL g2271 ( 
.A(n_2214),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2222),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2221),
.B(n_2192),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2224),
.B(n_2199),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2222),
.Y(n_2275)
);

OR2x6_ASAP7_75t_L g2276 ( 
.A(n_2214),
.B(n_2174),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2218),
.B(n_2205),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2242),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2220),
.B(n_2216),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2221),
.B(n_2192),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2242),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2243),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_2228),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2243),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2250),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2217),
.B(n_2211),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2214),
.B(n_2174),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_2236),
.Y(n_2288)
);

INVxp67_ASAP7_75t_SL g2289 ( 
.A(n_2246),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2239),
.B(n_2174),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_2227),
.B(n_2083),
.Y(n_2291)
);

AOI21xp33_ASAP7_75t_L g2292 ( 
.A1(n_2238),
.A2(n_2145),
.B(n_2186),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2232),
.B(n_2173),
.Y(n_2293)
);

OAI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_2233),
.A2(n_2175),
.B(n_2176),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2225),
.B(n_2211),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2250),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2253),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2230),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2264),
.B(n_2176),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2239),
.B(n_2169),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2225),
.B(n_2147),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2253),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_L g2303 ( 
.A(n_2240),
.B(n_2127),
.Y(n_2303)
);

INVx2_ASAP7_75t_SL g2304 ( 
.A(n_2236),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2229),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2229),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2254),
.Y(n_2307)
);

AOI22xp33_ASAP7_75t_L g2308 ( 
.A1(n_2274),
.A2(n_2233),
.B1(n_2226),
.B2(n_2231),
.Y(n_2308)
);

INVx1_ASAP7_75t_SL g2309 ( 
.A(n_2267),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2298),
.B(n_2254),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2307),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2288),
.B(n_2246),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2273),
.B(n_2247),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2273),
.B(n_2247),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2272),
.Y(n_2315)
);

AOI222xp33_ASAP7_75t_L g2316 ( 
.A1(n_2277),
.A2(n_2251),
.B1(n_2169),
.B2(n_2262),
.C1(n_2234),
.C2(n_2252),
.Y(n_2316)
);

INVx1_ASAP7_75t_SL g2317 ( 
.A(n_2271),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_2283),
.B(n_2256),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2288),
.Y(n_2319)
);

NAND3xp33_ASAP7_75t_L g2320 ( 
.A(n_2279),
.B(n_2215),
.C(n_2244),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2272),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2303),
.B(n_2234),
.Y(n_2322)
);

BUFx2_ASAP7_75t_L g2323 ( 
.A(n_2304),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2275),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2275),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2278),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2278),
.Y(n_2327)
);

NOR2xp33_ASAP7_75t_SL g2328 ( 
.A(n_2270),
.B(n_2252),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2304),
.Y(n_2329)
);

OAI21x1_ASAP7_75t_L g2330 ( 
.A1(n_2294),
.A2(n_2289),
.B(n_2300),
.Y(n_2330)
);

OR2x2_ASAP7_75t_L g2331 ( 
.A(n_2266),
.B(n_2256),
.Y(n_2331)
);

NOR2x1_ASAP7_75t_L g2332 ( 
.A(n_2276),
.B(n_2257),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2266),
.Y(n_2333)
);

AND3x1_ASAP7_75t_L g2334 ( 
.A(n_2287),
.B(n_2257),
.C(n_2261),
.Y(n_2334)
);

INVxp67_ASAP7_75t_L g2335 ( 
.A(n_2286),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2281),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2307),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2281),
.Y(n_2338)
);

OAI21xp33_ASAP7_75t_L g2339 ( 
.A1(n_2308),
.A2(n_2295),
.B(n_2301),
.Y(n_2339)
);

O2A1O1Ixp33_ASAP7_75t_L g2340 ( 
.A1(n_2309),
.A2(n_2316),
.B(n_2317),
.C(n_2292),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2311),
.Y(n_2341)
);

OAI21xp33_ASAP7_75t_SL g2342 ( 
.A1(n_2330),
.A2(n_2300),
.B(n_2280),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2311),
.Y(n_2343)
);

OAI322xp33_ASAP7_75t_L g2344 ( 
.A1(n_2328),
.A2(n_2306),
.A3(n_2305),
.B1(n_2268),
.B2(n_2297),
.C1(n_2296),
.C2(n_2282),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_2322),
.B(n_2268),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2332),
.A2(n_2276),
.B1(n_2306),
.B2(n_2305),
.Y(n_2346)
);

AOI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2334),
.A2(n_2287),
.B1(n_2276),
.B2(n_2280),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2315),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2313),
.A2(n_2276),
.B1(n_2290),
.B2(n_2261),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2323),
.Y(n_2350)
);

AOI221xp5_ASAP7_75t_L g2351 ( 
.A1(n_2320),
.A2(n_2269),
.B1(n_2282),
.B2(n_2297),
.C(n_2296),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2335),
.B(n_2291),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_L g2353 ( 
.A1(n_2313),
.A2(n_2290),
.B1(n_2293),
.B2(n_2248),
.Y(n_2353)
);

AOI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2314),
.A2(n_2330),
.B1(n_2329),
.B2(n_2319),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2315),
.Y(n_2355)
);

AOI221xp5_ASAP7_75t_L g2356 ( 
.A1(n_2321),
.A2(n_2302),
.B1(n_2284),
.B2(n_2285),
.C(n_2244),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2327),
.Y(n_2357)
);

AO21x1_ASAP7_75t_L g2358 ( 
.A1(n_2319),
.A2(n_2248),
.B(n_2260),
.Y(n_2358)
);

INVxp67_ASAP7_75t_SL g2359 ( 
.A(n_2323),
.Y(n_2359)
);

OAI322xp33_ASAP7_75t_L g2360 ( 
.A1(n_2318),
.A2(n_2293),
.A3(n_2299),
.B1(n_2248),
.B2(n_2263),
.C1(n_2259),
.C2(n_2215),
.Y(n_2360)
);

AOI22xp33_ASAP7_75t_R g2361 ( 
.A1(n_2350),
.A2(n_2339),
.B1(n_2340),
.B2(n_2344),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2359),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2341),
.Y(n_2363)
);

NAND2x1_ASAP7_75t_L g2364 ( 
.A(n_2346),
.B(n_2312),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2343),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2345),
.Y(n_2366)
);

INVx2_ASAP7_75t_SL g2367 ( 
.A(n_2346),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_2352),
.B(n_2314),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2347),
.B(n_2329),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2351),
.B(n_2333),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2348),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2355),
.B(n_2333),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2357),
.Y(n_2373)
);

OR2x6_ASAP7_75t_L g2374 ( 
.A(n_2358),
.B(n_2318),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_2368),
.B(n_2349),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2370),
.A2(n_2342),
.B1(n_2354),
.B2(n_2353),
.Y(n_2376)
);

AOI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2370),
.A2(n_2356),
.B1(n_2312),
.B2(n_2258),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2367),
.B(n_2324),
.Y(n_2378)
);

OAI211xp5_ASAP7_75t_SL g2379 ( 
.A1(n_2366),
.A2(n_2338),
.B(n_2336),
.C(n_2325),
.Y(n_2379)
);

AOI21xp33_ASAP7_75t_L g2380 ( 
.A1(n_2364),
.A2(n_2374),
.B(n_2362),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2369),
.B(n_2326),
.Y(n_2381)
);

AOI211x1_ASAP7_75t_L g2382 ( 
.A1(n_2372),
.A2(n_2337),
.B(n_2327),
.C(n_2258),
.Y(n_2382)
);

O2A1O1Ixp33_ASAP7_75t_L g2383 ( 
.A1(n_2374),
.A2(n_2360),
.B(n_2337),
.C(n_2310),
.Y(n_2383)
);

NOR3xp33_ASAP7_75t_L g2384 ( 
.A(n_2372),
.B(n_2310),
.C(n_2331),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_SL g2385 ( 
.A(n_2374),
.B(n_2312),
.Y(n_2385)
);

OAI221xp5_ASAP7_75t_SL g2386 ( 
.A1(n_2361),
.A2(n_2331),
.B1(n_2260),
.B2(n_2299),
.C(n_2241),
.Y(n_2386)
);

AOI22x1_ASAP7_75t_SL g2387 ( 
.A1(n_2380),
.A2(n_2373),
.B1(n_2365),
.B2(n_2363),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2378),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2382),
.Y(n_2389)
);

AOI31xp33_ASAP7_75t_R g2390 ( 
.A1(n_2385),
.A2(n_2361),
.A3(n_2371),
.B(n_2028),
.Y(n_2390)
);

NOR2x1_ASAP7_75t_L g2391 ( 
.A(n_2383),
.B(n_2259),
.Y(n_2391)
);

OAI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2376),
.A2(n_2263),
.B(n_2249),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_2381),
.B(n_2245),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2377),
.Y(n_2394)
);

O2A1O1Ixp5_ASAP7_75t_L g2395 ( 
.A1(n_2386),
.A2(n_2249),
.B(n_2245),
.C(n_2237),
.Y(n_2395)
);

XNOR2xp5_ASAP7_75t_L g2396 ( 
.A(n_2387),
.B(n_2394),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2391),
.B(n_2375),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2389),
.B(n_2384),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2392),
.B(n_2237),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2392),
.B(n_2255),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2393),
.Y(n_2401)
);

NOR3x1_ASAP7_75t_L g2402 ( 
.A(n_2388),
.B(n_2379),
.C(n_2265),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2395),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_R g2404 ( 
.A(n_2396),
.B(n_2390),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2401),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2397),
.Y(n_2406)
);

AOI222xp33_ASAP7_75t_L g2407 ( 
.A1(n_2403),
.A2(n_2184),
.B1(n_2182),
.B2(n_2209),
.C1(n_2213),
.C2(n_2183),
.Y(n_2407)
);

OR2x2_ASAP7_75t_L g2408 ( 
.A(n_2399),
.B(n_2255),
.Y(n_2408)
);

INVxp67_ASAP7_75t_L g2409 ( 
.A(n_2398),
.Y(n_2409)
);

OAI211xp5_ASAP7_75t_L g2410 ( 
.A1(n_2404),
.A2(n_2400),
.B(n_2402),
.C(n_2265),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2405),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2406),
.A2(n_2200),
.B(n_2177),
.Y(n_2412)
);

BUFx2_ASAP7_75t_L g2413 ( 
.A(n_2408),
.Y(n_2413)
);

XNOR2x1_ASAP7_75t_L g2414 ( 
.A(n_2411),
.B(n_2413),
.Y(n_2414)
);

OAI22xp33_ASAP7_75t_SL g2415 ( 
.A1(n_2414),
.A2(n_2409),
.B1(n_2412),
.B2(n_2410),
.Y(n_2415)
);

HB1xp67_ASAP7_75t_L g2416 ( 
.A(n_2415),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_2415),
.B(n_2407),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2416),
.B(n_2177),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2417),
.Y(n_2419)
);

INVx3_ASAP7_75t_L g2420 ( 
.A(n_2419),
.Y(n_2420)
);

OAI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2418),
.A2(n_2193),
.B1(n_2178),
.B2(n_2212),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2420),
.Y(n_2422)
);

AOI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_2422),
.A2(n_2421),
.B1(n_2028),
.B2(n_2186),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2423),
.B(n_2204),
.Y(n_2424)
);

NAND3xp33_ASAP7_75t_L g2425 ( 
.A(n_2424),
.B(n_2028),
.C(n_2182),
.Y(n_2425)
);

AOI22xp5_ASAP7_75t_L g2426 ( 
.A1(n_2425),
.A2(n_2185),
.B1(n_2193),
.B2(n_2212),
.Y(n_2426)
);

AOI211xp5_ASAP7_75t_L g2427 ( 
.A1(n_2426),
.A2(n_2028),
.B(n_1952),
.C(n_1990),
.Y(n_2427)
);


endmodule