module fake_ariane_836_n_176 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_176);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_176;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_156;
wire n_96;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_128;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_121;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_26),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx2_ASAP7_75t_SL g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_12),
.B(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_34),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_0),
.Y(n_52)
);

NOR2x1p5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_1),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_4),
.Y(n_54)
);

BUFx8_ASAP7_75t_SL g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_27),
.B(n_4),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_5),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_8),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_10),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_12),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_13),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_48),
.B(n_45),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_54),
.B(n_52),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_30),
.B(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_30),
.Y(n_80)
);

NAND2x1p5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_32),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_32),
.B(n_16),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_50),
.B(n_68),
.C(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_13),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_51),
.B1(n_63),
.B2(n_53),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_62),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AOI21x1_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_58),
.B(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_56),
.B1(n_51),
.B2(n_68),
.Y(n_98)
);

CKINVDCx6p67_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

AO21x2_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_76),
.B(n_77),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_86),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_81),
.B(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_98),
.B1(n_87),
.B2(n_72),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_78),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_90),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_57),
.B1(n_56),
.B2(n_49),
.C(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_90),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_80),
.B(n_82),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_101),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_118),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_107),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_107),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_103),
.Y(n_127)
);

AOI222xp33_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_111),
.B1(n_57),
.B2(n_49),
.C1(n_54),
.C2(n_52),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_84),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_102),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_85),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_102),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_55),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_55),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_129),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_59),
.C(n_66),
.Y(n_139)
);

AOI211xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_59),
.B(n_66),
.C(n_52),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_120),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NOR3x1_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_66),
.C(n_64),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_128),
.C(n_81),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_128),
.C(n_81),
.Y(n_146)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_142),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_133),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_120),
.B1(n_102),
.B2(n_64),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_122),
.Y(n_150)
);

AND3x1_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_61),
.C(n_60),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_102),
.B1(n_61),
.B2(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_100),
.C(n_105),
.Y(n_156)
);

NAND4xp75_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_100),
.C(n_105),
.D(n_97),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_104),
.Y(n_158)
);

NOR2x1p5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_99),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_104),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_100),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_102),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

AND3x4_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_94),
.C(n_104),
.Y(n_166)
);

NAND5xp2_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_105),
.C(n_100),
.D(n_77),
.E(n_95),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_99),
.B1(n_104),
.B2(n_93),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_93),
.A3(n_97),
.B1(n_96),
.B2(n_89),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_93),
.C(n_96),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_93),
.C(n_99),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_166),
.B1(n_162),
.B2(n_158),
.Y(n_172)
);

OAI21x1_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_161),
.B(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_162),
.Y(n_174)
);

OAI21x1_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_174),
.B(n_172),
.Y(n_175)
);

OAI221xp5_ASAP7_75t_R g176 ( 
.A1(n_175),
.A2(n_171),
.B1(n_169),
.B2(n_159),
.C(n_163),
.Y(n_176)
);


endmodule