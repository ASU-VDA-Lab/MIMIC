module fake_aes_8207_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
INVx4_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
CKINVDCx5p33_ASAP7_75t_R g4 ( .A(n_1), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
AOI22xp5_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_4), .B1(n_3), .B2(n_1), .Y(n_8) );
AOI22xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_3), .B1(n_6), .B2(n_0), .Y(n_9) );
AOI211xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_6), .B(n_7), .C(n_3), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
AOI22xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_2), .B1(n_10), .B2(n_9), .Y(n_12) );
endmodule