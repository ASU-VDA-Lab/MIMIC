module real_jpeg_26492_n_16 (n_5, n_4, n_8, n_0, n_12, n_339, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_339;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_46),
.B1(n_57),
.B2(n_60),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_0),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_46),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_1),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_115),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_57),
.B1(n_60),
.B2(n_115),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_115),
.Y(n_253)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_2),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_2),
.A2(n_135),
.B(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_2),
.Y(n_213)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_4),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_120),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_120),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_4),
.A2(n_57),
.B1(n_60),
.B2(n_120),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_6),
.A2(n_24),
.B1(n_51),
.B2(n_52),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_6),
.A2(n_24),
.B1(n_57),
.B2(n_60),
.Y(n_157)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_8),
.A2(n_11),
.B(n_57),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_44),
.B1(n_57),
.B2(n_60),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_10),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_35),
.B1(n_57),
.B2(n_60),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_11),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_11),
.B(n_29),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_11),
.A2(n_29),
.B(n_161),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_118),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_77),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_99),
.B1(n_100),
.B2(n_212),
.Y(n_215)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_67),
.Y(n_73)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_14),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_15),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_15),
.A2(n_22),
.B1(n_23),
.B2(n_113),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_15),
.A2(n_51),
.B1(n_52),
.B2(n_113),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_15),
.A2(n_57),
.B1(n_60),
.B2(n_113),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_84),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_20),
.A2(n_42),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_21),
.A2(n_31),
.B(n_81),
.Y(n_297)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_25),
.B(n_26),
.C(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_22),
.B(n_118),
.CON(n_117),
.SN(n_117)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_25),
.A2(n_31),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_26),
.B(n_29),
.Y(n_132)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_28),
.A2(n_32),
.B1(n_117),
.B2(n_132),
.Y(n_131)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_51),
.A3(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_30),
.A2(n_43),
.B(n_47),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_31),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_47),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_74),
.C(n_79),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_38),
.A2(n_39),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_48),
.C(n_63),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_40),
.A2(n_41),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_42),
.A2(n_47),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_42),
.A2(n_47),
.B1(n_126),
.B2(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_47),
.B(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_48),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_48),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_48),
.A2(n_63),
.B1(n_306),
.B2(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_56),
.B(n_61),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_49),
.A2(n_61),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_49),
.A2(n_56),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_49),
.A2(n_169),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_49),
.A2(n_56),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_49),
.A2(n_56),
.B1(n_168),
.B2(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_49),
.A2(n_56),
.B1(n_94),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_49),
.A2(n_108),
.B(n_246),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_52),
.B(n_66),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_52),
.A2(n_55),
.B(n_118),
.C(n_189),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_60),
.Y(n_56)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_56),
.B(n_118),
.Y(n_210)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_100),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_60),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_62),
.B(n_109),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_63),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_64),
.A2(n_76),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_72),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_65),
.A2(n_72),
.B1(n_112),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_65),
.A2(n_72),
.B1(n_144),
.B2(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_65),
.B(n_71),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_65),
.A2(n_72),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_70),
.A2(n_77),
.B(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_76),
.A2(n_78),
.B(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_76),
.A2(n_256),
.B(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_79),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_331),
.B(n_337),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_301),
.A3(n_323),
.B1(n_329),
.B2(n_330),
.C(n_339),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_282),
.B(n_300),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_260),
.B(n_281),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_149),
.B(n_236),
.C(n_259),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_136),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_90),
.B(n_136),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_121),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_105),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_92),
.B(n_105),
.C(n_121),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_93),
.B(n_98),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_95),
.B(n_179),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B(n_102),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_99),
.A2(n_197),
.B(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_99),
.A2(n_204),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_99),
.A2(n_213),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_104),
.Y(n_103)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_100),
.B(n_118),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_130),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_123),
.B(n_128),
.C(n_130),
.Y(n_257)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_133),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_137),
.A2(n_138),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_148),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_235),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_228),
.B(n_234),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_180),
.B(n_227),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_170),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_153),
.B(n_170),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.C(n_166),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_154),
.A2(n_155),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_199),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_177),
.C(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_221),
.B(n_226),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_200),
.B(n_220),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_183),
.B(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_208),
.B(n_219),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_206),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_214),
.B(n_218),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_222),
.B(n_223),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_229),
.B(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_238),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_257),
.B2(n_258),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_248),
.C(n_258),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_251),
.C(n_255),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_262),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_280),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_274),
.C(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_269),
.C(n_271),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_275),
.A2(n_276),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_278),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_294),
.B(n_297),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_284),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_298),
.B2(n_299),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_293),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_293),
.C(n_299),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B(n_292),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_291),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_303),
.C(n_313),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_303),
.B1(n_304),
.B2(n_328),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_292),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_315),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_315),
.Y(n_330)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_304)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_310),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_312),
.B1(n_317),
.B2(n_321),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_321),
.C(n_322),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_314),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_322),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);


endmodule