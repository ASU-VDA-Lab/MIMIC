module fake_jpeg_14375_n_426 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_65),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_7),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_48),
.B(n_50),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_14),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_49),
.B(n_75),
.C(n_44),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_16),
.B(n_6),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_52),
.Y(n_138)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_6),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_6),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_61),
.B(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_66),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_9),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_30),
.B(n_5),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_69),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_5),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_10),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_2),
.C(n_3),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_32),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_13),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_31),
.B1(n_40),
.B2(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_89),
.A2(n_98),
.B1(n_109),
.B2(n_27),
.Y(n_158)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_38),
.B1(n_40),
.B2(n_44),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_116),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_66),
.B1(n_70),
.B2(n_60),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_102),
.A2(n_111),
.B1(n_117),
.B2(n_130),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_57),
.A2(n_40),
.B1(n_27),
.B2(n_26),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_59),
.A2(n_40),
.B1(n_21),
.B2(n_37),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_62),
.A2(n_81),
.B1(n_85),
.B2(n_84),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_45),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_79),
.B1(n_64),
.B2(n_73),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_33),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_76),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_55),
.B(n_41),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_29),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_49),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_140),
.B(n_147),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_27),
.B(n_26),
.C(n_44),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_141),
.A2(n_96),
.B(n_113),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_142),
.B(n_153),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_157),
.C(n_159),
.Y(n_194)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_33),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_82),
.B1(n_80),
.B2(n_78),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_151),
.A2(n_108),
.B1(n_92),
.B2(n_107),
.Y(n_192)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_95),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_89),
.A2(n_36),
.B1(n_43),
.B2(n_35),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_178),
.B1(n_101),
.B2(n_106),
.Y(n_201)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_35),
.C(n_32),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_180),
.B1(n_187),
.B2(n_107),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_33),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_26),
.B1(n_39),
.B2(n_29),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_160),
.A2(n_186),
.B1(n_96),
.B2(n_113),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_0),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_0),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_164),
.B(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_29),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_166),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_0),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_2),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_177),
.C(n_182),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_39),
.B(n_3),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_105),
.A2(n_28),
.B1(n_4),
.B2(n_11),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_170),
.A2(n_178),
.B(n_177),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_98),
.A2(n_2),
.B(n_4),
.C(n_11),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_173),
.Y(n_198)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_12),
.B(n_13),
.C(n_28),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_12),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_115),
.A2(n_28),
.B1(n_12),
.B2(n_13),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_28),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_115),
.A2(n_28),
.B1(n_123),
.B2(n_124),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_127),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_112),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_183),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_129),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_96),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_108),
.A2(n_124),
.B1(n_106),
.B2(n_92),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_192),
.A2(n_201),
.B1(n_204),
.B2(n_210),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_199),
.A2(n_213),
.B1(n_214),
.B2(n_221),
.Y(n_247)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_200),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_148),
.A2(n_101),
.B1(n_119),
.B2(n_131),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_208),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_209),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_148),
.A2(n_119),
.B1(n_131),
.B2(n_132),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_158),
.A2(n_119),
.B1(n_131),
.B2(n_132),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_179),
.B(n_177),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_154),
.A2(n_164),
.B1(n_165),
.B2(n_140),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_173),
.Y(n_238)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

AO21x2_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_113),
.B(n_171),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_180),
.A2(n_181),
.B1(n_176),
.B2(n_172),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_152),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_228),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_162),
.A2(n_155),
.B1(n_170),
.B2(n_163),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_155),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_231),
.B(n_233),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_143),
.C(n_159),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_243),
.C(n_248),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_216),
.B(n_143),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_153),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_234),
.B(n_239),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_235),
.A2(n_219),
.B(n_196),
.Y(n_293)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_238),
.B(n_226),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_191),
.B(n_157),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_221),
.A2(n_149),
.B1(n_144),
.B2(n_187),
.Y(n_241)
);

AOI22x1_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_253),
.B1(n_201),
.B2(n_221),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_184),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_246),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_161),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_161),
.C(n_182),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_212),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_263),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_191),
.B(n_168),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_214),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_141),
.B1(n_175),
.B2(n_168),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_182),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_257),
.C(n_259),
.Y(n_291)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_197),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_SL g257 ( 
.A(n_209),
.B(n_193),
.C(n_198),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_211),
.Y(n_258)
);

INVx6_ASAP7_75t_SL g290 ( 
.A(n_258),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_174),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_205),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_146),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_220),
.B(n_142),
.Y(n_263)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_203),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_272),
.C(n_287),
.Y(n_305)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_221),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_273),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_238),
.A2(n_198),
.B(n_215),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_227),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_281),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_207),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_251),
.A2(n_189),
.B1(n_205),
.B2(n_213),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_276),
.A2(n_282),
.B1(n_254),
.B2(n_250),
.Y(n_303)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_277),
.Y(n_298)
);

CKINVDCx10_ASAP7_75t_R g280 ( 
.A(n_236),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_199),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_189),
.B1(n_223),
.B2(n_196),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_296),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_190),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_219),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_260),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_251),
.B(n_293),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_303),
.Y(n_340)
);

AOI22x1_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_247),
.B1(n_262),
.B2(n_241),
.Y(n_302)
);

AOI22x1_ASAP7_75t_SL g342 ( 
.A1(n_302),
.A2(n_279),
.B1(n_285),
.B2(n_280),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_245),
.B1(n_262),
.B2(n_250),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_306),
.A2(n_309),
.B1(n_316),
.B2(n_275),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_245),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_307),
.B(n_312),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_266),
.A2(n_245),
.B1(n_290),
.B2(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_278),
.B(n_256),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_278),
.A2(n_244),
.B1(n_248),
.B2(n_235),
.Y(n_313)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_265),
.A2(n_230),
.B1(n_264),
.B2(n_237),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_315),
.Y(n_328)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_229),
.B(n_225),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_190),
.C(n_222),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_322),
.C(n_287),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_270),
.A2(n_274),
.B1(n_265),
.B2(n_269),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_319),
.A2(n_296),
.B1(n_279),
.B2(n_267),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_222),
.C(n_225),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_271),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_325),
.B(n_332),
.Y(n_359)
);

BUFx12_ASAP7_75t_L g326 ( 
.A(n_311),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_268),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_331),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_338),
.C(n_347),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_291),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_323),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_291),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_337),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_319),
.B(n_290),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_321),
.B(n_272),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_336),
.B(n_343),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_284),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_288),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_323),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_342),
.B1(n_345),
.B2(n_309),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_346),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_301),
.B(n_285),
.Y(n_343)
);

FAx1_ASAP7_75t_SL g346 ( 
.A(n_308),
.B(n_294),
.CI(n_174),
.CON(n_346),
.SN(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_310),
.C(n_320),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_300),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_345),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_367),
.Y(n_369)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_358),
.Y(n_376)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_327),
.Y(n_361)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_361),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_306),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_365),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_336),
.B(n_317),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_363),
.B(n_337),
.Y(n_370)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_300),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_299),
.B1(n_316),
.B2(n_320),
.Y(n_366)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_366),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_298),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_347),
.A2(n_299),
.B1(n_297),
.B2(n_302),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_368),
.A2(n_341),
.B1(n_340),
.B2(n_342),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_374),
.Y(n_390)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_371),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_329),
.C(n_331),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_375),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_338),
.C(n_340),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_363),
.B(n_340),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_360),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_351),
.A2(n_346),
.B(n_302),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_382),
.A2(n_349),
.B(n_367),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_368),
.A2(n_298),
.B1(n_324),
.B2(n_315),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_381),
.B(n_356),
.C(n_354),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_386),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_371),
.Y(n_385)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_377),
.B(n_350),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_356),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_362),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_375),
.A2(n_359),
.B(n_355),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_393),
.Y(n_397)
);

OAI221xp5_ASAP7_75t_L g396 ( 
.A1(n_391),
.A2(n_395),
.B1(n_372),
.B2(n_380),
.C(n_379),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g395 ( 
.A1(n_369),
.A2(n_349),
.B(n_365),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_396),
.A2(n_326),
.B1(n_346),
.B2(n_304),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_373),
.C(n_354),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_400),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_387),
.A2(n_374),
.B(n_383),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_403),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_376),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_370),
.C(n_378),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_229),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_392),
.B(n_311),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_405),
.A2(n_240),
.B1(n_146),
.B2(n_200),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_404),
.A2(n_392),
.B1(n_390),
.B2(n_382),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_412),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_397),
.A2(n_390),
.B(n_393),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_409),
.A2(n_411),
.B(n_413),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_410),
.Y(n_417)
);

OAI322xp33_ASAP7_75t_L g411 ( 
.A1(n_399),
.A2(n_360),
.A3(n_326),
.B1(n_294),
.B2(n_304),
.C1(n_237),
.C2(n_195),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_406),
.B(n_398),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_414),
.A2(n_407),
.B(n_409),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_397),
.C(n_402),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_412),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_419),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_421),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_417),
.A2(n_240),
.B(n_206),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g424 ( 
.A1(n_423),
.A2(n_417),
.A3(n_416),
.B1(n_418),
.B2(n_218),
.C1(n_174),
.C2(n_240),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_424),
.A2(n_422),
.B(n_206),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_195),
.Y(n_426)
);


endmodule