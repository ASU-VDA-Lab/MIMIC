module fake_netlist_5_890_n_794 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_794);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_794;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_679;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_45),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_51),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_44),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_34),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_38),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_54),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_96),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_122),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_52),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_80),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_7),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_95),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_107),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_74),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_128),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_126),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_81),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_148),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_63),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_13),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_124),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_5),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_97),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_37),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_90),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_10),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_75),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_69),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_93),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_151),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_121),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_19),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_98),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_144),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_113),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_116),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_53),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_117),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_162),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_170),
.B(n_0),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_177),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_161),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_163),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_188),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_165),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_166),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_169),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_172),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_167),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_174),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_175),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_179),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_180),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_182),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_183),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_215),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_189),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_217),
.B(n_199),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_223),
.Y(n_279)
);

BUFx8_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

AND2x6_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_18),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_247),
.A2(n_216),
.B1(n_214),
.B2(n_213),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_184),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_256),
.B(n_185),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_258),
.B(n_186),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_218),
.A2(n_212),
.B1(n_211),
.B2(n_208),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_218),
.A2(n_207),
.B(n_205),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_219),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_219),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_221),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_222),
.B(n_190),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_225),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_232),
.B(n_20),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

INVx4_ASAP7_75t_SL g309 ( 
.A(n_307),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

NAND3x1_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_238),
.C(n_2),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_263),
.B(n_193),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_262),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_194),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_306),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_196),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_267),
.A2(n_283),
.B1(n_307),
.B2(n_282),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_265),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_21),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_267),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_198),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_267),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_204),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_284),
.B(n_203),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_1),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_279),
.B(n_22),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_1),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_2),
.C(n_3),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_292),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_264),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_283),
.B(n_3),
.Y(n_340)
);

INVx4_ASAP7_75t_SL g341 ( 
.A(n_307),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_4),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_287),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_264),
.B(n_159),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_268),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_4),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_303),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_SL g349 ( 
.A(n_297),
.B(n_5),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_6),
.Y(n_350)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_281),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_270),
.Y(n_352)
);

NAND2xp33_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_6),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_303),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_288),
.B(n_7),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_8),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_277),
.Y(n_358)
);

INVx6_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_295),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_291),
.B(n_8),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_277),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_266),
.B(n_23),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_285),
.B(n_9),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_274),
.B(n_24),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_276),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_276),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_276),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_275),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_271),
.B(n_266),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_266),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_296),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_317),
.B(n_296),
.Y(n_376)
);

OAI221xp5_ASAP7_75t_L g377 ( 
.A1(n_347),
.A2(n_296),
.B1(n_305),
.B2(n_271),
.C(n_294),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_363),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_265),
.Y(n_380)
);

AO22x2_ASAP7_75t_L g381 ( 
.A1(n_336),
.A2(n_308),
.B1(n_299),
.B2(n_298),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_317),
.B(n_265),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_298),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_328),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_299),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_304),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_335),
.A2(n_281),
.B1(n_300),
.B2(n_308),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_354),
.Y(n_394)
);

OR2x2_ASAP7_75t_SL g395 ( 
.A(n_359),
.B(n_301),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_354),
.B(n_304),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_326),
.B(n_281),
.Y(n_398)
);

OR2x2_ASAP7_75t_SL g399 ( 
.A(n_359),
.B(n_302),
.Y(n_399)
);

AO22x2_ASAP7_75t_L g400 ( 
.A1(n_336),
.A2(n_302),
.B1(n_304),
.B2(n_306),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

AO22x2_ASAP7_75t_L g402 ( 
.A1(n_367),
.A2(n_306),
.B1(n_286),
.B2(n_272),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_300),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_321),
.A2(n_293),
.B1(n_11),
.B2(n_12),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_281),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_281),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_321),
.B(n_281),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_322),
.Y(n_412)
);

OAI221xp5_ASAP7_75t_L g413 ( 
.A1(n_356),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_327),
.Y(n_415)
);

NAND2x1p5_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_280),
.Y(n_416)
);

NAND2x1p5_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_280),
.Y(n_417)
);

BUFx8_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_14),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_337),
.B(n_25),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_337),
.B(n_26),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

A2O1A1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_342),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_372),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_320),
.B(n_15),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_329),
.B(n_316),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_320),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_360),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_311),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_311),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_361),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_357),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_350),
.A2(n_16),
.B1(n_17),
.B2(n_27),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_358),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_358),
.B(n_28),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_310),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g444 ( 
.A(n_361),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_375),
.B(n_309),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_376),
.B(n_309),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_394),
.B(n_341),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_316),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_394),
.B(n_341),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_384),
.B(n_351),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_411),
.B(n_351),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_414),
.B(n_351),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_318),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_392),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_390),
.B(n_362),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_333),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_415),
.B(n_345),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_412),
.B(n_345),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_389),
.B(n_349),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_397),
.B(n_368),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_388),
.B(n_387),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_380),
.B(n_368),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_404),
.B(n_313),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_404),
.B(n_385),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_419),
.B(n_332),
.Y(n_465)
);

XNOR2x2_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_314),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_438),
.B(n_334),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_410),
.B(n_323),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_378),
.B(n_353),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_422),
.B(n_426),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_396),
.B(n_323),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_405),
.B(n_323),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_405),
.B(n_323),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_393),
.B(n_30),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_401),
.B(n_17),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_393),
.B(n_442),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_442),
.B(n_403),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_408),
.B(n_31),
.Y(n_478)
);

NAND2xp33_ASAP7_75t_SL g479 ( 
.A(n_437),
.B(n_406),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_409),
.B(n_32),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_424),
.B(n_420),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_379),
.B(n_433),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_434),
.B(n_33),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_407),
.B(n_35),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_382),
.B(n_36),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_377),
.B(n_39),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_SL g487 ( 
.A(n_398),
.B(n_40),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_SL g488 ( 
.A(n_398),
.B(n_41),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_SL g489 ( 
.A(n_383),
.B(n_42),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_386),
.B(n_43),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_SL g491 ( 
.A(n_391),
.B(n_46),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_443),
.B(n_48),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_439),
.B(n_49),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_SL g494 ( 
.A(n_435),
.B(n_50),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_440),
.B(n_55),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_431),
.B(n_56),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_441),
.B(n_57),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_436),
.B(n_58),
.Y(n_498)
);

AO31x2_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_423),
.A3(n_428),
.B(n_432),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_454),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_453),
.A2(n_429),
.B(n_425),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_476),
.A2(n_402),
.B(n_381),
.Y(n_502)
);

AO31x2_ASAP7_75t_L g503 ( 
.A1(n_486),
.A2(n_381),
.A3(n_400),
.B(n_402),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_448),
.B(n_400),
.Y(n_504)
);

OAI21x1_ASAP7_75t_SL g505 ( 
.A1(n_490),
.A2(n_410),
.B(n_413),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_462),
.A2(n_410),
.B(n_417),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_444),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_455),
.B(n_418),
.Y(n_508)
);

AO31x2_ASAP7_75t_L g509 ( 
.A1(n_471),
.A2(n_410),
.A3(n_399),
.B(n_395),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_416),
.Y(n_510)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_474),
.A2(n_60),
.B(n_61),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_456),
.B(n_418),
.Y(n_512)
);

AO31x2_ASAP7_75t_L g513 ( 
.A1(n_492),
.A2(n_62),
.A3(n_64),
.B(n_65),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_456),
.B(n_158),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

OAI21x1_ASAP7_75t_SL g516 ( 
.A1(n_466),
.A2(n_66),
.B(n_67),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_458),
.B(n_68),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_459),
.B(n_70),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_468),
.A2(n_71),
.B(n_72),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_469),
.A2(n_73),
.B(n_76),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_467),
.B(n_78),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_79),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_464),
.B(n_82),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_460),
.A2(n_83),
.B(n_84),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_481),
.A2(n_85),
.B(n_86),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_463),
.A2(n_87),
.B(n_88),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_472),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_465),
.Y(n_530)
);

BUFx2_ASAP7_75t_R g531 ( 
.A(n_447),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_473),
.A2(n_493),
.B1(n_457),
.B2(n_446),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_479),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_450),
.B(n_94),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_484),
.A2(n_100),
.B(n_101),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_102),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_445),
.B(n_103),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_451),
.B(n_156),
.Y(n_540)
);

AOI21xp33_ASAP7_75t_L g541 ( 
.A1(n_452),
.A2(n_105),
.B(n_106),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_480),
.B(n_109),
.Y(n_542)
);

A2O1A1Ixp33_ASAP7_75t_L g543 ( 
.A1(n_502),
.A2(n_491),
.B(n_494),
.C(n_487),
.Y(n_543)
);

OAI221xp5_ASAP7_75t_L g544 ( 
.A1(n_508),
.A2(n_485),
.B1(n_488),
.B2(n_483),
.C(n_498),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_500),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_519),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g547 ( 
.A1(n_505),
.A2(n_497),
.B(n_495),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_530),
.Y(n_548)
);

AO31x2_ASAP7_75t_L g549 ( 
.A1(n_533),
.A2(n_110),
.A3(n_111),
.B(n_112),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_506),
.A2(n_114),
.B(n_115),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_532),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_512),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_504),
.A2(n_120),
.B1(n_125),
.B2(n_127),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_501),
.A2(n_129),
.B(n_130),
.Y(n_554)
);

AND3x2_ASAP7_75t_L g555 ( 
.A(n_512),
.B(n_518),
.C(n_507),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_525),
.A2(n_131),
.B(n_132),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_524),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_520),
.A2(n_135),
.B(n_137),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_524),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_515),
.B(n_139),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_499),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_499),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_526),
.A2(n_140),
.B(n_142),
.Y(n_563)
);

A2O1A1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_537),
.A2(n_143),
.B(n_145),
.C(n_146),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_514),
.A2(n_147),
.B(n_150),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_535),
.A2(n_152),
.B(n_153),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g567 ( 
.A1(n_516),
.A2(n_155),
.B1(n_538),
.B2(n_510),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_534),
.B(n_517),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_521),
.A2(n_527),
.B(n_528),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_522),
.A2(n_536),
.B1(n_511),
.B2(n_523),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_540),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_503),
.B(n_499),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_529),
.A2(n_542),
.B1(n_541),
.B2(n_531),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_503),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_503),
.B(n_509),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_509),
.B(n_513),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_513),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_509),
.A2(n_466),
.B1(n_493),
.B2(n_335),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_500),
.B(n_448),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_508),
.B(n_375),
.C(n_384),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_500),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_515),
.B(n_524),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_524),
.B(n_500),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_574),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_561),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_584),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_584),
.Y(n_588)
);

CKINVDCx11_ASAP7_75t_R g589 ( 
.A(n_552),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_584),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_574),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_583),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_545),
.B(n_582),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_582),
.Y(n_595)
);

AO21x2_ASAP7_75t_L g596 ( 
.A1(n_576),
.A2(n_543),
.B(n_575),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_548),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_562),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_548),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_572),
.B(n_579),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_546),
.B(n_580),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_550),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_568),
.B(n_578),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_550),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_577),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_569),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_551),
.B(n_549),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

NAND2x1p5_ASAP7_75t_L g609 ( 
.A(n_554),
.B(n_563),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_554),
.A2(n_569),
.B(n_563),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_583),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_549),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_549),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_558),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_558),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_547),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_547),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_547),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_568),
.B(n_555),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_543),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_571),
.Y(n_623)
);

AOI21xp33_ASAP7_75t_L g624 ( 
.A1(n_581),
.A2(n_573),
.B(n_544),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_557),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_571),
.Y(n_626)
);

BUFx2_ASAP7_75t_SL g627 ( 
.A(n_559),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_560),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_564),
.Y(n_631)
);

AO21x2_ASAP7_75t_L g632 ( 
.A1(n_565),
.A2(n_566),
.B(n_570),
.Y(n_632)
);

CKINVDCx6p67_ASAP7_75t_R g633 ( 
.A(n_567),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_553),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_594),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_R g636 ( 
.A(n_589),
.B(n_592),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_624),
.B(n_590),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_601),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_R g639 ( 
.A(n_621),
.B(n_587),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_R g640 ( 
.A(n_592),
.B(n_612),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_587),
.Y(n_641)
);

BUFx4f_ASAP7_75t_L g642 ( 
.A(n_621),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_588),
.B(n_601),
.Y(n_643)
);

BUFx2_ASAP7_75t_R g644 ( 
.A(n_634),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_R g645 ( 
.A(n_621),
.B(n_587),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_600),
.B(n_611),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_587),
.B(n_592),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_594),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_612),
.B(n_611),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_600),
.B(n_612),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_585),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_628),
.B(n_634),
.Y(n_652)
);

CKINVDCx12_ASAP7_75t_R g653 ( 
.A(n_628),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_R g654 ( 
.A(n_618),
.B(n_603),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_625),
.B(n_593),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_625),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_618),
.B(n_593),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g658 ( 
.A(n_603),
.B(n_626),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_595),
.B(n_597),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_622),
.B(n_595),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_R g661 ( 
.A(n_607),
.B(n_631),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_599),
.B(n_622),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_599),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_633),
.B(n_607),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_R g666 ( 
.A(n_633),
.B(n_626),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_R g667 ( 
.A(n_630),
.B(n_631),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_623),
.B(n_585),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_R g669 ( 
.A(n_630),
.B(n_623),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_627),
.B(n_634),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_627),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_591),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_591),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_598),
.B(n_586),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_R g676 ( 
.A(n_629),
.B(n_614),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_636),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_651),
.Y(n_678)
);

INVx1_ASAP7_75t_SL g679 ( 
.A(n_671),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_646),
.B(n_608),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_641),
.B(n_605),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_672),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_638),
.B(n_632),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_650),
.B(n_657),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_641),
.B(n_605),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_674),
.Y(n_686)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_643),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_675),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_675),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_664),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_657),
.B(n_614),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_668),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_668),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_637),
.B(n_632),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_659),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_635),
.B(n_613),
.Y(n_696)
);

INVxp33_ASAP7_75t_L g697 ( 
.A(n_658),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_648),
.B(n_613),
.Y(n_698)
);

AO21x2_ASAP7_75t_L g699 ( 
.A1(n_652),
.A2(n_615),
.B(n_610),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_660),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_667),
.Y(n_701)
);

AND2x4_ASAP7_75t_SL g702 ( 
.A(n_670),
.B(n_586),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_649),
.B(n_605),
.Y(n_703)
);

INVxp67_ASAP7_75t_SL g704 ( 
.A(n_669),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_644),
.B(n_629),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_665),
.B(n_596),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_640),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_678),
.Y(n_708)
);

INVx5_ASAP7_75t_SL g709 ( 
.A(n_699),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_701),
.A2(n_642),
.B1(n_647),
.B2(n_656),
.Y(n_710)
);

NOR2x1_ASAP7_75t_L g711 ( 
.A(n_707),
.B(n_662),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_677),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_682),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_686),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_690),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_694),
.A2(n_632),
.B1(n_697),
.B2(n_687),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_706),
.B(n_673),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_687),
.B(n_649),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_688),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_684),
.B(n_642),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_693),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_683),
.B(n_615),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_693),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_706),
.B(n_673),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_722),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_717),
.B(n_684),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_722),
.B(n_721),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_717),
.B(n_691),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_723),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_708),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_714),
.B(n_697),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_722),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_711),
.B(n_677),
.Y(n_733)
);

NOR2x1p5_ASAP7_75t_L g734 ( 
.A(n_712),
.B(n_704),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_724),
.B(n_691),
.Y(n_735)
);

AO221x2_ASAP7_75t_L g736 ( 
.A1(n_734),
.A2(n_710),
.B1(n_718),
.B2(n_715),
.C(n_719),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_731),
.B(n_716),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_733),
.A2(n_666),
.B1(n_731),
.B2(n_705),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_726),
.B(n_716),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_735),
.B(n_713),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_725),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_725),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_738),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_740),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_741),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_737),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_746),
.B(n_736),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_744),
.B(n_742),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_745),
.B(n_739),
.Y(n_749)
);

AOI21xp33_ASAP7_75t_SL g750 ( 
.A1(n_743),
.A2(n_732),
.B(n_727),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_748),
.B(n_732),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_749),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_747),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_751),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_752),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_751),
.Y(n_756)
);

BUFx4f_ASAP7_75t_SL g757 ( 
.A(n_753),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_754),
.B(n_750),
.Y(n_758)
);

NAND4xp25_ASAP7_75t_L g759 ( 
.A(n_756),
.B(n_712),
.C(n_679),
.D(n_639),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_757),
.B(n_730),
.Y(n_760)
);

NAND4xp25_ASAP7_75t_L g761 ( 
.A(n_755),
.B(n_645),
.C(n_661),
.D(n_654),
.Y(n_761)
);

AND4x1_ASAP7_75t_L g762 ( 
.A(n_757),
.B(n_720),
.C(n_724),
.D(n_728),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_758),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_759),
.A2(n_709),
.B1(n_722),
.B2(n_685),
.Y(n_764)
);

NOR4xp25_ASAP7_75t_L g765 ( 
.A(n_760),
.B(n_729),
.C(n_708),
.D(n_689),
.Y(n_765)
);

OAI221xp5_ASAP7_75t_L g766 ( 
.A1(n_762),
.A2(n_676),
.B1(n_723),
.B2(n_692),
.C(n_695),
.Y(n_766)
);

CKINVDCx6p67_ASAP7_75t_R g767 ( 
.A(n_761),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_758),
.A2(n_709),
.B1(n_723),
.B2(n_700),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_763),
.Y(n_769)
);

NAND4xp75_ASAP7_75t_L g770 ( 
.A(n_767),
.B(n_655),
.C(n_696),
.D(n_680),
.Y(n_770)
);

NAND4xp75_ASAP7_75t_L g771 ( 
.A(n_765),
.B(n_696),
.C(n_680),
.D(n_663),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_764),
.B(n_709),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_766),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_768),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_SL g775 ( 
.A(n_769),
.B(n_653),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_R g776 ( 
.A(n_774),
.B(n_660),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_SL g777 ( 
.A(n_773),
.B(n_772),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_771),
.B(n_681),
.Y(n_778)
);

NOR3xp33_ASAP7_75t_L g779 ( 
.A(n_777),
.B(n_770),
.C(n_606),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_775),
.Y(n_780)
);

XOR2xp5_ASAP7_75t_L g781 ( 
.A(n_778),
.B(n_685),
.Y(n_781)
);

OR4x1_ASAP7_75t_L g782 ( 
.A(n_780),
.B(n_776),
.C(n_779),
.D(n_781),
.Y(n_782)
);

AO21x2_ASAP7_75t_L g783 ( 
.A1(n_779),
.A2(n_699),
.B(n_610),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_SL g784 ( 
.A(n_780),
.B(n_609),
.C(n_698),
.Y(n_784)
);

OAI22x1_ASAP7_75t_L g785 ( 
.A1(n_780),
.A2(n_685),
.B1(n_681),
.B2(n_703),
.Y(n_785)
);

OAI22x1_ASAP7_75t_L g786 ( 
.A1(n_782),
.A2(n_681),
.B1(n_703),
.B2(n_609),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_783),
.Y(n_787)
);

AOI31xp33_ASAP7_75t_L g788 ( 
.A1(n_786),
.A2(n_784),
.A3(n_785),
.B(n_609),
.Y(n_788)
);

AOI31xp33_ASAP7_75t_L g789 ( 
.A1(n_787),
.A2(n_698),
.A3(n_703),
.B(n_616),
.Y(n_789)
);

OAI322xp33_ASAP7_75t_L g790 ( 
.A1(n_788),
.A2(n_616),
.A3(n_602),
.B1(n_604),
.B2(n_617),
.C1(n_620),
.C2(n_619),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_L g791 ( 
.A(n_790),
.B(n_789),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_791),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_R g793 ( 
.A1(n_792),
.A2(n_702),
.B1(n_699),
.B2(n_596),
.C(n_606),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_793),
.A2(n_602),
.B1(n_604),
.B2(n_619),
.Y(n_794)
);


endmodule