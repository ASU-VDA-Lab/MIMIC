module fake_netlist_1_11560_n_28 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_6), .B(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
NAND2xp5_ASAP7_75t_SL g22 ( .A(n_21), .B(n_19), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_15), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_0), .Y(n_24) );
A2O1A1Ixp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_17), .B(n_0), .C(n_3), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI322xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_2), .A3(n_5), .B1(n_7), .B2(n_10), .C1(n_11), .C2(n_13), .Y(n_28) );
endmodule