module fake_jpeg_17238_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_41),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_17),
.B1(n_20),
.B2(n_24),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_32),
.B1(n_30),
.B2(n_20),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_17),
.B1(n_24),
.B2(n_20),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_60),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_34),
.B1(n_25),
.B2(n_31),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_54),
.B(n_63),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_21),
.B(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_24),
.B1(n_20),
.B2(n_2),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_70),
.B1(n_0),
.B2(n_1),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_28),
.B1(n_31),
.B2(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g93 ( 
.A(n_65),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_26),
.B1(n_22),
.B2(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_77),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_38),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_39),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_62),
.B(n_22),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_83),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_89),
.Y(n_112)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_37),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_53),
.B1(n_56),
.B2(n_68),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_52),
.B(n_38),
.Y(n_95)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_102),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_68),
.B1(n_61),
.B2(n_48),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_86),
.B1(n_71),
.B2(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_80),
.B1(n_79),
.B2(n_95),
.Y(n_131)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_18),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_67),
.B1(n_62),
.B2(n_46),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_115),
.B1(n_116),
.B2(n_90),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_109),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_114),
.Y(n_137)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_69),
.B1(n_70),
.B2(n_26),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_69),
.B1(n_51),
.B2(n_59),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_65),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_22),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_65),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_96),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_59),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_91),
.B1(n_80),
.B2(n_75),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_138),
.B1(n_101),
.B2(n_117),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_88),
.B1(n_85),
.B2(n_75),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_131),
.B1(n_149),
.B2(n_103),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_111),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_143),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_88),
.B1(n_78),
.B2(n_89),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_71),
.C(n_79),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_139),
.C(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_93),
.C(n_81),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_100),
.B(n_19),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_99),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_27),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_81),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_81),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_96),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_108),
.B(n_109),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_26),
.B1(n_27),
.B2(n_19),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_156),
.A2(n_161),
.B1(n_176),
.B2(n_127),
.Y(n_197)
);

OA21x2_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_119),
.B(n_107),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_158),
.A2(n_159),
.B(n_18),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_103),
.B(n_119),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_160),
.A2(n_170),
.B(n_171),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_174),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_99),
.B(n_124),
.C(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_169),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_129),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_173),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_122),
.Y(n_169)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_110),
.B(n_106),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_136),
.C(n_153),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_139),
.C(n_131),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_129),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_179),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_111),
.B1(n_114),
.B2(n_102),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_114),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_2),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_148),
.B(n_142),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_192),
.A2(n_193),
.B(n_207),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_142),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_199),
.C(n_168),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_201),
.B1(n_165),
.B2(n_171),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_128),
.C(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_102),
.B(n_126),
.C(n_154),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_157),
.A2(n_156),
.B1(n_155),
.B2(n_158),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_204),
.B1(n_159),
.B2(n_182),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_155),
.A2(n_126),
.B1(n_149),
.B2(n_19),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_18),
.B(n_2),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_8),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_8),
.Y(n_212)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_174),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_222),
.C(n_226),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_221),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_177),
.B1(n_161),
.B2(n_169),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_231),
.B1(n_188),
.B2(n_201),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_SL g220 ( 
.A(n_189),
.B(n_163),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_228),
.B(n_190),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_172),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_160),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_184),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_223),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_174),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_165),
.B1(n_166),
.B2(n_175),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_201),
.B1(n_187),
.B2(n_204),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_208),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_210),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_237),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_2),
.C(n_3),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_16),
.C(n_5),
.Y(n_255)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_221),
.A2(n_201),
.B1(n_192),
.B2(n_205),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_249),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_194),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_251),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_193),
.B(n_201),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_252),
.B(n_256),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_193),
.B1(n_188),
.B2(n_190),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_227),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_207),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_206),
.B(n_4),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_3),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_218),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_233),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_4),
.B(n_6),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_213),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_219),
.C(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_232),
.C(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_270),
.B(n_257),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_223),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_274),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_227),
.C(n_235),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_239),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_230),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_286),
.C(n_287),
.Y(n_292)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_280),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_245),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_277),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_245),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_288),
.Y(n_291)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_244),
.B(n_258),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_267),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_243),
.B(n_254),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_247),
.B(n_256),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_290),
.B(n_295),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_263),
.C(n_259),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_300),
.C(n_4),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_259),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

INVx11_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_255),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_286),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_283),
.B(n_251),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_274),
.C(n_260),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_R g301 ( 
.A(n_297),
.B(n_292),
.Y(n_301)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_306),
.C(n_309),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_292),
.A2(n_267),
.B1(n_6),
.B2(n_7),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_289),
.A3(n_294),
.B1(n_296),
.B2(n_300),
.C1(n_12),
.C2(n_7),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_312),
.A3(n_13),
.B1(n_307),
.B2(n_311),
.C1(n_315),
.C2(n_313),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_9),
.B(n_10),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_9),
.C(n_10),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_13),
.B(n_14),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_317),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_313),
.B(n_318),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.Y(n_322)
);


endmodule