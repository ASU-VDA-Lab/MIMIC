module fake_jpeg_13596_n_64 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_1),
.B(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_18),
.B(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_31),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_28),
.C(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_24),
.CON(n_37),
.SN(n_37)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_22),
.B1(n_23),
.B2(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_15),
.B1(n_27),
.B2(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_41),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_31),
.B(n_9),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_16),
.C(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_27),
.B1(n_16),
.B2(n_14),
.Y(n_45)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

AO221x1_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_37),
.B1(n_9),
.B2(n_20),
.C(n_3),
.Y(n_49)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_47),
.B1(n_48),
.B2(n_3),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_51),
.B(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

AOI322xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_61),
.A3(n_51),
.B1(n_56),
.B2(n_54),
.C1(n_53),
.C2(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);


endmodule