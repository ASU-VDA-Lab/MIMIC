module fake_jpeg_20447_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_42),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_55),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_28),
.B1(n_20),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_51),
.B1(n_61),
.B2(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_28),
.B1(n_20),
.B2(n_33),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_26),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_26),
.Y(n_90)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_45),
.B1(n_41),
.B2(n_40),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_43),
.B1(n_37),
.B2(n_30),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_64),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_66),
.B(n_69),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_43),
.B1(n_37),
.B2(n_18),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_67),
.A2(n_83),
.B1(n_84),
.B2(n_89),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_74),
.B(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_44),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_38),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_98),
.B(n_99),
.Y(n_107)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_38),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_93),
.B(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_45),
.B1(n_41),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_55),
.B1(n_41),
.B2(n_40),
.Y(n_104)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_78),
.B(n_85),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_87),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_82),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_27),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_101),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_27),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_27),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_21),
.C(n_32),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_97),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_25),
.B(n_19),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_24),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_55),
.B1(n_63),
.B2(n_45),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_112),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_55),
.B1(n_39),
.B2(n_25),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_55),
.C(n_26),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_116),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_34),
.B1(n_31),
.B2(n_23),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_127),
.B1(n_122),
.B2(n_109),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_26),
.C(n_24),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_86),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_89),
.B(n_79),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_31),
.B1(n_23),
.B2(n_34),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_26),
.C(n_24),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_135),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_155),
.B1(n_77),
.B2(n_130),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_94),
.B(n_95),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_145),
.B(n_112),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_94),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_76),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_98),
.B(n_76),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_81),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_149),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_81),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_71),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_97),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_157),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_72),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_106),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_159),
.B(n_168),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_160),
.A2(n_178),
.B(n_128),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_185),
.B(n_149),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_116),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_134),
.B(n_133),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_113),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_131),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_170),
.B(n_175),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_103),
.C(n_106),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_135),
.C(n_144),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_126),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_126),
.B1(n_104),
.B2(n_105),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_180),
.B1(n_138),
.B2(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_125),
.B1(n_82),
.B2(n_119),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_195),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_207),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_155),
.B1(n_145),
.B2(n_139),
.C(n_135),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_203),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_209),
.C(n_169),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_194),
.B1(n_196),
.B2(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_139),
.B1(n_151),
.B2(n_136),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_154),
.Y(n_195)
);

OAI321xp33_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_151),
.A3(n_143),
.B1(n_153),
.B2(n_132),
.C(n_129),
.Y(n_196)
);

OAI322xp33_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_153),
.A3(n_19),
.B1(n_34),
.B2(n_31),
.C1(n_23),
.C2(n_5),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_206),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_204),
.Y(n_226)
);

AOI221xp5_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_19),
.B1(n_34),
.B2(n_31),
.C(n_102),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

OAI322xp33_ASAP7_75t_L g206 ( 
.A1(n_186),
.A2(n_10),
.A3(n_16),
.B1(n_15),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_102),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_187),
.A2(n_171),
.B1(n_160),
.B2(n_174),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_210),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_172),
.C(n_161),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_217),
.C(n_221),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_172),
.C(n_161),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_163),
.B1(n_162),
.B2(n_183),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_175),
.C(n_174),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_160),
.B1(n_170),
.B2(n_179),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_197),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_205),
.B(n_183),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_188),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_176),
.C(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.C(n_202),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_176),
.C(n_173),
.Y(n_229)
);

NAND4xp25_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_204),
.C(n_200),
.D(n_163),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_247),
.B(n_230),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_236),
.C(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_240),
.Y(n_260)
);

NOR3xp33_ASAP7_75t_SL g237 ( 
.A(n_224),
.B(n_207),
.C(n_202),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_243),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_189),
.C(n_195),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_238),
.A2(n_217),
.B(n_221),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_227),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_10),
.Y(n_257)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_244),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_173),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_218),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_198),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_0),
.B(n_1),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_249),
.B(n_250),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_228),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_213),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_254),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_232),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_242),
.A2(n_218),
.B1(n_75),
.B2(n_2),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_239),
.B1(n_246),
.B2(n_2),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_259),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_247),
.C(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_11),
.C(n_3),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_238),
.B(n_239),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.C(n_269),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_240),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_237),
.B(n_233),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_255),
.B1(n_258),
.B2(n_250),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_6),
.B(n_7),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_6),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_275),
.C(n_270),
.Y(n_278)
);

NOR2x1_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_8),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_277),
.B(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_280),
.A2(n_281),
.B(n_13),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_272),
.B(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_9),
.C(n_12),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_12),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_286),
.B(n_279),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_14),
.B(n_15),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_16),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_287),
.B(n_15),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_291),
.Y(n_292)
);


endmodule