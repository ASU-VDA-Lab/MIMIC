module fake_jpeg_16743_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx4f_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_2),
.B(n_5),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_19),
.B1(n_22),
.B2(n_23),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.C(n_1),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.Y(n_24)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_11),
.B(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_7),
.B1(n_3),
.B2(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_9),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_12),
.B1(n_14),
.B2(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_31),
.B1(n_26),
.B2(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_27),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_24),
.C(n_20),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_24),
.B1(n_22),
.B2(n_29),
.Y(n_39)
);

AOI221xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.C(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_10),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_36),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_35),
.C(n_34),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_24),
.B1(n_29),
.B2(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_37),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_41),
.B(n_39),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_13),
.C(n_8),
.Y(n_47)
);

AOI322xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_8),
.A3(n_29),
.B1(n_16),
.B2(n_13),
.C1(n_45),
.C2(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_5),
.Y(n_49)
);


endmodule