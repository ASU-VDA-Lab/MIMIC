module fake_netlist_1_12637_n_692 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_692);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_692;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_42), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_17), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_63), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_93), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_30), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_90), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_31), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_98), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_95), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_91), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_35), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_105), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_104), .Y(n_120) );
CKINVDCx14_ASAP7_75t_R g121 ( .A(n_15), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_1), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_97), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_100), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_34), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_11), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_6), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_0), .Y(n_128) );
BUFx10_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_0), .Y(n_130) );
BUFx10_ASAP7_75t_L g131 ( .A(n_50), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_96), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_59), .B(n_18), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_64), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_7), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_18), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_47), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_54), .Y(n_138) );
INVxp67_ASAP7_75t_SL g139 ( .A(n_65), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_46), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_4), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_86), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_41), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_49), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_52), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_8), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_21), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_4), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_33), .Y(n_149) );
INVx2_ASAP7_75t_SL g150 ( .A(n_66), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_5), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_121), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
INVx2_ASAP7_75t_SL g155 ( .A(n_129), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_138), .Y(n_156) );
INVx6_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_138), .Y(n_159) );
BUFx8_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_147), .B(n_2), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_109), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_112), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_150), .B(n_3), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_114), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_117), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_119), .Y(n_168) );
BUFx8_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_136), .B(n_5), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_161), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_161), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
INVx6_ASAP7_75t_L g176 ( .A(n_160), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_160), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
OAI22xp33_ASAP7_75t_L g181 ( .A1(n_152), .A2(n_128), .B1(n_146), .B2(n_122), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
XNOR2x1_ASAP7_75t_L g183 ( .A(n_170), .B(n_148), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_153), .B(n_154), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_158), .B(n_131), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_158), .B(n_120), .Y(n_187) );
OR2x6_ASAP7_75t_L g188 ( .A(n_158), .B(n_127), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_160), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_153), .B(n_132), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_158), .B(n_131), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_156), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_156), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_157), .B(n_144), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
BUFx10_ASAP7_75t_L g197 ( .A(n_157), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_179), .A2(n_164), .B(n_155), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_186), .B(n_157), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_174), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_186), .B(n_191), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_179), .B(n_169), .Y(n_203) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_183), .A2(n_128), .B1(n_146), .B2(n_122), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_174), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g206 ( .A1(n_183), .A2(n_169), .B1(n_157), .B2(n_113), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_186), .B(n_191), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_176), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_191), .B(n_172), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_172), .B(n_173), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_173), .B(n_175), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_179), .B(n_169), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_194), .B(n_155), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_189), .B(n_169), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_176), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_175), .A2(n_171), .B1(n_168), .B2(n_167), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_174), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_194), .B(n_160), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_174), .A2(n_171), .B(n_168), .C(n_167), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_163), .B(n_162), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_188), .A2(n_163), .B1(n_162), .B2(n_165), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_187), .B(n_165), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_184), .Y(n_225) );
AND2x2_ASAP7_75t_L g226 ( .A(n_188), .B(n_154), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_185), .A2(n_166), .B(n_159), .C(n_151), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_185), .B(n_182), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_188), .B(n_166), .Y(n_229) );
OR2x6_ASAP7_75t_L g230 ( .A(n_188), .B(n_166), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_180), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_180), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_182), .B(n_111), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_223), .B(n_189), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_204), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_230), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_230), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_202), .B(n_188), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_202), .B(n_188), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_207), .B(n_183), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_209), .B(n_182), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_228), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
NAND3xp33_ASAP7_75t_L g244 ( .A(n_206), .B(n_181), .C(n_190), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_230), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_190), .B(n_176), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_211), .A2(n_176), .B(n_196), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_211), .A2(n_176), .B(n_196), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_212), .A2(n_176), .B(n_195), .Y(n_249) );
AOI33xp33_ASAP7_75t_L g250 ( .A1(n_217), .A2(n_181), .A3(n_135), .B1(n_130), .B2(n_141), .B3(n_149), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_201), .A2(n_198), .B(n_177), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_220), .A2(n_198), .B(n_133), .C(n_139), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_230), .A2(n_198), .B1(n_113), .B2(n_118), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_209), .B(n_197), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_230), .A2(n_118), .B1(n_197), .B2(n_148), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_200), .B(n_197), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_210), .B(n_197), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_212), .A2(n_198), .B(n_108), .C(n_126), .Y(n_258) );
NOR2x1p5_ASAP7_75t_SL g259 ( .A(n_210), .B(n_201), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
NOR3xp33_ASAP7_75t_L g261 ( .A(n_200), .B(n_111), .C(n_115), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_229), .A2(n_198), .B1(n_115), .B2(n_143), .Y(n_262) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_226), .B(n_140), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_258), .A2(n_227), .B(n_214), .C(n_224), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_246), .A2(n_229), .B(n_218), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_240), .B(n_226), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_252), .A2(n_213), .B(n_215), .C(n_203), .Y(n_268) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_249), .A2(n_199), .B(n_232), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_251), .A2(n_232), .B(n_231), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_236), .B(n_205), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_218), .B(n_221), .C(n_225), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_247), .A2(n_232), .B(n_231), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_248), .A2(n_231), .B(n_221), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_260), .A2(n_253), .B1(n_255), .B2(n_238), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_245), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_244), .A2(n_225), .B(n_219), .C(n_233), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_240), .B(n_197), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_234), .A2(n_195), .B(n_177), .Y(n_279) );
AOI21x1_ASAP7_75t_SL g280 ( .A1(n_239), .A2(n_131), .B(n_208), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_236), .Y(n_281) );
NOR2xp33_ASAP7_75t_SL g282 ( .A(n_245), .B(n_216), .Y(n_282) );
AOI221x1_ASAP7_75t_L g283 ( .A1(n_261), .A2(n_180), .B1(n_192), .B2(n_177), .C(n_178), .Y(n_283) );
BUFx10_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_250), .B(n_180), .C(n_192), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_253), .B(n_6), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_263), .B(n_216), .Y(n_287) );
OAI22x1_ASAP7_75t_L g288 ( .A1(n_235), .A2(n_107), .B1(n_110), .B2(n_125), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_272), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_281), .B(n_236), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_273), .Y(n_291) );
OA21x2_ASAP7_75t_L g292 ( .A1(n_277), .A2(n_178), .B(n_195), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_286), .A2(n_237), .B1(n_263), .B2(n_236), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_279), .A2(n_234), .B(n_257), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_275), .A2(n_237), .B1(n_243), .B2(n_241), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_277), .A2(n_254), .B(n_243), .Y(n_296) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_265), .A2(n_272), .B(n_278), .C(n_268), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_281), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_281), .Y(n_299) );
AO21x1_ASAP7_75t_L g300 ( .A1(n_266), .A2(n_257), .B(n_256), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_281), .B(n_259), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_273), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_267), .B(n_262), .Y(n_303) );
BUFx2_ASAP7_75t_L g304 ( .A(n_276), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_278), .A2(n_134), .B1(n_137), .B2(n_142), .C(n_145), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_285), .A2(n_208), .B(n_178), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_279), .A2(n_180), .B(n_192), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_284), .Y(n_310) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_297), .A2(n_274), .B(n_269), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_297), .A2(n_269), .B(n_270), .Y(n_312) );
OA21x2_ASAP7_75t_L g313 ( .A1(n_302), .A2(n_291), .B(n_294), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_289), .B(n_276), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_302), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_302), .Y(n_316) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_302), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_289), .B(n_271), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_301), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_291), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_295), .B(n_271), .Y(n_322) );
OAI21x1_ASAP7_75t_L g323 ( .A1(n_294), .A2(n_280), .B(n_283), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_301), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_292), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_301), .B(n_271), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_292), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_301), .B(n_287), .Y(n_328) );
AO31x2_ASAP7_75t_L g329 ( .A1(n_300), .A2(n_287), .A3(n_288), .B(n_282), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_292), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_292), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_292), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_301), .B(n_7), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_303), .B(n_293), .Y(n_334) );
AO21x2_ASAP7_75t_L g335 ( .A1(n_296), .A2(n_180), .B(n_192), .Y(n_335) );
AO21x2_ASAP7_75t_L g336 ( .A1(n_296), .A2(n_180), .B(n_192), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_316), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_333), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_320), .B(n_299), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_316), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_320), .B(n_299), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_316), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_324), .B(n_299), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_318), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_324), .B(n_298), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_333), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_320), .B(n_298), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_317), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_324), .B(n_304), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_300), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_321), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_321), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_334), .B(n_303), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_334), .B(n_293), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_320), .B(n_304), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_314), .B(n_307), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_328), .B(n_300), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_321), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_326), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_314), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_333), .B(n_304), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_313), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_314), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_337), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_326), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_328), .B(n_295), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_328), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_326), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_326), .B(n_294), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_326), .B(n_305), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_367), .B(n_325), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_374), .B(n_331), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_338), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_367), .B(n_325), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_363), .B(n_319), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_372), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_349), .B(n_307), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_374), .B(n_331), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_341), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_325), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_381), .B(n_8), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_370), .B(n_327), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_373), .B(n_327), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_373), .B(n_327), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_355), .B(n_330), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_356), .B(n_330), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_356), .B(n_330), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_339), .B(n_319), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_380), .B(n_337), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_345), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_354), .B(n_307), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_345), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_347), .Y(n_406) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_354), .B(n_307), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_348), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_380), .B(n_337), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_346), .Y(n_410) );
NOR2xp33_ASAP7_75t_R g411 ( .A(n_374), .B(n_307), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_341), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_369), .B(n_331), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_343), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_348), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_353), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_378), .B(n_329), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_347), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_354), .B(n_331), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_369), .B(n_332), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_351), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_364), .B(n_329), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_375), .B(n_332), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_351), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_352), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_355), .B(n_332), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_375), .B(n_377), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_344), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_371), .B(n_329), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_371), .B(n_329), .Y(n_430) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_357), .B(n_305), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_343), .B(n_329), .Y(n_432) );
NOR2x1_ASAP7_75t_SL g433 ( .A(n_365), .B(n_310), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_352), .B(n_329), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_379), .B(n_332), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_365), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_376), .B(n_311), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_357), .B(n_311), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_358), .B(n_311), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_358), .B(n_311), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_359), .B(n_311), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_359), .B(n_311), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_376), .B(n_312), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_361), .Y(n_444) );
INVx3_ASAP7_75t_L g445 ( .A(n_360), .Y(n_445) );
AND2x4_ASAP7_75t_SL g446 ( .A(n_406), .B(n_366), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_403), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_418), .B(n_361), .Y(n_448) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_431), .B(n_310), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_383), .B(n_362), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_433), .B(n_350), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_433), .B(n_350), .Y(n_452) );
NOR4xp25_ASAP7_75t_L g453 ( .A(n_393), .B(n_322), .C(n_340), .D(n_342), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_383), .B(n_362), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g455 ( .A(n_389), .B(n_310), .Y(n_455) );
OR2x6_ASAP7_75t_L g456 ( .A(n_404), .B(n_366), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_382), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_405), .Y(n_458) );
OR2x6_ASAP7_75t_L g459 ( .A(n_404), .B(n_407), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_382), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_416), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_416), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_410), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_428), .B(n_368), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_386), .B(n_342), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_411), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_397), .B(n_360), .Y(n_468) );
BUFx2_ASAP7_75t_SL g469 ( .A(n_416), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_401), .B(n_366), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_388), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_422), .B(n_329), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_445), .Y(n_473) );
NAND2xp67_ASAP7_75t_L g474 ( .A(n_392), .B(n_322), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_427), .B(n_329), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_425), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_401), .B(n_329), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_409), .B(n_312), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_409), .B(n_312), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_398), .B(n_312), .Y(n_480) );
NAND2x1p5_ASAP7_75t_L g481 ( .A(n_445), .B(n_419), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_385), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_398), .B(n_312), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_397), .B(n_313), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_391), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_412), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_388), .Y(n_487) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_417), .B(n_306), .C(n_10), .D(n_11), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_399), .B(n_312), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_414), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_426), .B(n_313), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_404), .B(n_290), .Y(n_492) );
NOR2x2_ASAP7_75t_L g493 ( .A(n_402), .B(n_9), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_444), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_402), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_445), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_436), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_426), .B(n_313), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_399), .B(n_313), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_435), .B(n_313), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_435), .B(n_335), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_394), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_413), .B(n_335), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_394), .B(n_335), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_395), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_395), .B(n_335), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_396), .B(n_335), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_413), .B(n_335), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_396), .B(n_336), .Y(n_509) );
NAND2xp33_ASAP7_75t_L g510 ( .A(n_407), .B(n_290), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_423), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_423), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_407), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_408), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_420), .B(n_387), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_420), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_408), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_432), .B(n_336), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_443), .B(n_336), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_443), .B(n_336), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_502), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_475), .B(n_434), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_505), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_473), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_449), .A2(n_429), .B1(n_430), .B2(n_390), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_500), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_475), .B(n_441), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_497), .B(n_400), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g529 ( .A(n_488), .B(n_438), .C(n_440), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_470), .B(n_437), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_488), .B(n_438), .C(n_440), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_515), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_466), .B(n_437), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_482), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_512), .B(n_439), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_487), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_448), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_485), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_472), .B(n_441), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_516), .B(n_384), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_472), .B(n_439), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_451), .B(n_384), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_451), .B(n_384), .Y(n_543) );
AO22x1_ASAP7_75t_L g544 ( .A1(n_467), .A2(n_390), .B1(n_419), .B2(n_421), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_486), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_490), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_465), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_495), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_452), .B(n_390), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_494), .Y(n_551) );
OAI32xp33_ASAP7_75t_L g552 ( .A1(n_449), .A2(n_442), .A3(n_290), .B1(n_421), .B2(n_415), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_452), .B(n_419), .Y(n_553) );
OAI21xp33_ASAP7_75t_SL g554 ( .A1(n_453), .A2(n_442), .B(n_424), .Y(n_554) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_459), .B(n_415), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_477), .B(n_424), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_447), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_512), .B(n_336), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_495), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_458), .Y(n_560) );
AOI222xp33_ASAP7_75t_L g561 ( .A1(n_480), .A2(n_306), .B1(n_10), .B2(n_12), .C1(n_13), .C2(n_14), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_483), .B(n_489), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_463), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_464), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_499), .B(n_336), .Y(n_565) );
AOI21xp33_ASAP7_75t_L g566 ( .A1(n_518), .A2(n_9), .B(n_12), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_480), .B(n_323), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_446), .B(n_323), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_453), .A2(n_290), .B(n_323), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_517), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_511), .B(n_323), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_450), .B(n_13), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_491), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_510), .A2(n_308), .B(n_309), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_450), .B(n_14), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_469), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_476), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_454), .B(n_15), .Y(n_578) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_457), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g580 ( .A1(n_474), .A2(n_308), .B(n_192), .Y(n_580) );
AND2x2_ASAP7_75t_SL g581 ( .A(n_493), .B(n_309), .Y(n_581) );
OA21x2_ASAP7_75t_L g582 ( .A1(n_518), .A2(n_309), .B(n_17), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_478), .B(n_479), .Y(n_583) );
INVx2_ASAP7_75t_SL g584 ( .A(n_468), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_460), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_484), .B(n_16), .Y(n_586) );
OAI322xp33_ASAP7_75t_L g587 ( .A1(n_503), .A2(n_16), .A3(n_19), .B1(n_20), .B2(n_21), .C1(n_192), .C2(n_193), .Y(n_587) );
NOR2xp33_ASAP7_75t_SL g588 ( .A(n_581), .B(n_459), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_534), .Y(n_589) );
OA22x2_ASAP7_75t_L g590 ( .A1(n_576), .A2(n_459), .B1(n_456), .B2(n_492), .Y(n_590) );
OAI21xp5_ASAP7_75t_SL g591 ( .A1(n_561), .A2(n_455), .B(n_481), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_554), .A2(n_456), .B(n_492), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_533), .B(n_519), .Y(n_594) );
OAI32xp33_ASAP7_75t_L g595 ( .A1(n_529), .A2(n_455), .A3(n_481), .B1(n_513), .B2(n_498), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_522), .B(n_520), .Y(n_596) );
NOR3xp33_ASAP7_75t_SL g597 ( .A(n_586), .B(n_514), .C(n_20), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_509), .B1(n_504), .B2(n_507), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_584), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_506), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_522), .B(n_471), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_539), .A2(n_508), .B(n_501), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_545), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_537), .B(n_456), .Y(n_604) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_561), .A2(n_462), .B(n_461), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_547), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_551), .Y(n_607) );
OAI32xp33_ASAP7_75t_L g608 ( .A1(n_531), .A2(n_496), .A3(n_492), .B1(n_19), .B2(n_193), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_541), .B(n_309), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_553), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_579), .Y(n_611) );
AOI332xp33_ASAP7_75t_L g612 ( .A1(n_532), .A2(n_193), .A3(n_23), .B1(n_24), .B2(n_25), .B3(n_26), .C1(n_27), .C2(n_28), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_539), .B(n_309), .Y(n_613) );
NAND3xp33_ASAP7_75t_SL g614 ( .A(n_580), .B(n_22), .C(n_29), .Y(n_614) );
AOI21xp33_ASAP7_75t_SL g615 ( .A1(n_544), .A2(n_32), .B(n_36), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_566), .A2(n_193), .B(n_38), .Y(n_616) );
INVx2_ASAP7_75t_SL g617 ( .A(n_542), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_525), .A2(n_193), .B1(n_39), .B2(n_40), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_557), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_583), .B(n_37), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_560), .Y(n_621) );
NAND2xp33_ASAP7_75t_SL g622 ( .A(n_543), .B(n_43), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_572), .A2(n_44), .B1(n_45), .B2(n_48), .Y(n_623) );
CKINVDCx14_ASAP7_75t_R g624 ( .A(n_550), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_540), .B(n_51), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_563), .Y(n_626) );
AOI221x1_ASAP7_75t_L g627 ( .A1(n_578), .A2(n_53), .B1(n_55), .B2(n_56), .C(n_57), .Y(n_627) );
NAND4xp25_ASAP7_75t_SL g628 ( .A(n_555), .B(n_58), .C(n_60), .D(n_61), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_575), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_570), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_527), .A2(n_62), .B(n_67), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_528), .A2(n_587), .B1(n_548), .B2(n_541), .C(n_527), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_591), .A2(n_578), .B(n_566), .C(n_569), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_590), .A2(n_526), .B1(n_573), .B2(n_521), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_595), .A2(n_552), .B(n_569), .C(n_565), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_630), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_611), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_632), .A2(n_605), .B1(n_629), .B2(n_608), .C(n_602), .Y(n_638) );
INVx2_ASAP7_75t_SL g639 ( .A(n_599), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_592), .A2(n_524), .B(n_570), .C(n_582), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_601), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_605), .A2(n_523), .B1(n_524), .B2(n_564), .C(n_577), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_620), .B(n_582), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_615), .A2(n_568), .B(n_558), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_590), .A2(n_567), .B1(n_571), .B2(n_556), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_618), .B(n_567), .C(n_585), .Y(n_647) );
OAI21xp33_ASAP7_75t_L g648 ( .A1(n_598), .A2(n_556), .B(n_562), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_619), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_597), .A2(n_559), .B(n_549), .C(n_546), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_588), .A2(n_562), .B1(n_536), .B2(n_574), .C1(n_535), .C2(n_73), .Y(n_651) );
AO221x1_ASAP7_75t_L g652 ( .A1(n_618), .A2(n_624), .B1(n_622), .B2(n_593), .C(n_606), .Y(n_652) );
NOR2xp67_ASAP7_75t_SL g653 ( .A(n_616), .B(n_574), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_604), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_628), .A2(n_71), .B(n_74), .C(n_75), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_610), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_621), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_616), .A2(n_79), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g659 ( .A1(n_612), .A2(n_84), .B(n_85), .C(n_87), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_614), .A2(n_88), .B(n_89), .C(n_92), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_589), .A2(n_94), .B1(n_99), .B2(n_101), .C(n_102), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_627), .A2(n_216), .B(n_103), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_623), .A2(n_106), .B(n_631), .C(n_625), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_617), .A2(n_596), .B1(n_594), .B2(n_600), .Y(n_664) );
AOI221x1_ASAP7_75t_L g665 ( .A1(n_603), .A2(n_607), .B1(n_626), .B2(n_609), .C(n_613), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_632), .B(n_630), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_608), .A2(n_595), .B(n_591), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_591), .A2(n_592), .B(n_554), .Y(n_668) );
NAND4xp25_ASAP7_75t_L g669 ( .A(n_667), .B(n_668), .C(n_666), .D(n_638), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_635), .B(n_640), .C(n_643), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_633), .A2(n_650), .B(n_659), .C(n_645), .Y(n_671) );
NOR5xp2_ASAP7_75t_L g672 ( .A(n_649), .B(n_663), .C(n_648), .D(n_652), .E(n_658), .Y(n_672) );
NAND4xp25_ASAP7_75t_SL g673 ( .A(n_651), .B(n_634), .C(n_646), .D(n_643), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g674 ( .A1(n_653), .A2(n_654), .B(n_656), .C(n_639), .Y(n_674) );
NAND3xp33_ASAP7_75t_SL g675 ( .A(n_651), .B(n_655), .C(n_660), .Y(n_675) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_669), .B(n_656), .Y(n_676) );
NAND4xp75_ASAP7_75t_L g677 ( .A(n_672), .B(n_665), .C(n_662), .D(n_637), .Y(n_677) );
NAND3xp33_ASAP7_75t_SL g678 ( .A(n_671), .B(n_644), .C(n_654), .Y(n_678) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_674), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_679), .B(n_670), .Y(n_680) );
NOR3xp33_ASAP7_75t_SL g681 ( .A(n_678), .B(n_673), .C(n_675), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_676), .A2(n_636), .B1(n_664), .B2(n_647), .Y(n_682) );
INVxp67_ASAP7_75t_L g683 ( .A(n_680), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_682), .B(n_677), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_683), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_684), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_686), .B(n_681), .Y(n_687) );
INVx1_ASAP7_75t_SL g688 ( .A(n_685), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_688), .Y(n_689) );
AO21x2_ASAP7_75t_L g690 ( .A1(n_689), .A2(n_687), .B(n_661), .Y(n_690) );
AO21x2_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_641), .B(n_642), .Y(n_691) );
AOI21xp33_ASAP7_75t_SL g692 ( .A1(n_691), .A2(n_644), .B(n_657), .Y(n_692) );
endmodule