module fake_jpeg_7737_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_1),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_26),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_22),
.B1(n_35),
.B2(n_18),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_22),
.B1(n_64),
.B2(n_63),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_13),
.Y(n_105)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_87),
.Y(n_113)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_78),
.B1(n_82),
.B2(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_50),
.Y(n_101)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_89),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_25),
.B(n_17),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_84),
.Y(n_110)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_22),
.B1(n_35),
.B2(n_25),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_35),
.B1(n_52),
.B2(n_57),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_48),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_19),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_84),
.Y(n_116)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_92),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_106),
.B1(n_107),
.B2(n_115),
.Y(n_123)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_59),
.B(n_66),
.C(n_35),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_82),
.B1(n_78),
.B2(n_72),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_109),
.C(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_40),
.C(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_116),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_111),
.Y(n_142)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_70),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_118),
.B(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_28),
.B1(n_16),
.B2(n_27),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_16),
.B1(n_40),
.B2(n_42),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_82),
.B1(n_79),
.B2(n_72),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_134),
.B1(n_133),
.B2(n_130),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_137),
.B1(n_102),
.B2(n_96),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_10),
.C(n_15),
.Y(n_159)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_128),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_135),
.C(n_99),
.Y(n_152)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_134),
.B(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_77),
.C(n_69),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_68),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_91),
.C(n_81),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_125),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_94),
.A2(n_78),
.B1(n_81),
.B2(n_91),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_115),
.B1(n_106),
.B2(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_105),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_38),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_123),
.B1(n_144),
.B2(n_132),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_174),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_160),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_98),
.B(n_69),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_172),
.B(n_124),
.Y(n_182)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_159),
.B(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_158),
.B1(n_36),
.B2(n_34),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_97),
.B1(n_102),
.B2(n_49),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_42),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_38),
.C(n_37),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_165),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_164),
.B(n_169),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_42),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_170),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_34),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_38),
.C(n_37),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_103),
.Y(n_171)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_75),
.B(n_23),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_37),
.C(n_36),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_178),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_120),
.A2(n_37),
.B(n_36),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_132),
.B(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_23),
.Y(n_179)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_180),
.B(n_184),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_182),
.A2(n_183),
.B(n_167),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_153),
.B(n_164),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_198),
.B1(n_202),
.B2(n_30),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_163),
.A2(n_142),
.B1(n_144),
.B2(n_75),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_200),
.B1(n_157),
.B2(n_168),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_154),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_191),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_14),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_197),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_24),
.B1(n_142),
.B2(n_33),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_162),
.A2(n_36),
.B1(n_34),
.B2(n_24),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_204),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_34),
.B1(n_24),
.B2(n_27),
.Y(n_205)
);

AO22x2_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_30),
.B1(n_29),
.B2(n_31),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_213),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_196),
.A2(n_149),
.B1(n_175),
.B2(n_176),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_222),
.B1(n_229),
.B2(n_205),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_160),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_186),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_190),
.B(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_214),
.Y(n_252)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_152),
.C(n_166),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_218),
.C(n_219),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_221),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_161),
.C(n_169),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_167),
.C(n_9),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_183),
.B(n_30),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_204),
.B1(n_197),
.B2(n_199),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_241),
.B1(n_209),
.B2(n_229),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_235),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_186),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_193),
.C(n_195),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_200),
.B1(n_195),
.B2(n_191),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_205),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_251),
.B1(n_229),
.B2(n_215),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_31),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_246),
.C(n_250),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_31),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_230),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_210),
.A2(n_29),
.B1(n_8),
.B2(n_3),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_244),
.B1(n_242),
.B2(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_265),
.B(n_234),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_31),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_212),
.B(n_229),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_8),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_238),
.B1(n_237),
.B2(n_235),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_262),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_265),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_277),
.B(n_6),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_7),
.B1(n_14),
.B2(n_4),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_276),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_7),
.C(n_13),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_259),
.C(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_261),
.B(n_259),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_284),
.A2(n_274),
.B(n_9),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_262),
.C(n_2),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_290),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_5),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_11),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_281),
.A2(n_5),
.B(n_6),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_278),
.B(n_273),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_299),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_279),
.B1(n_269),
.B2(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_298),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_289),
.B1(n_294),
.B2(n_287),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_11),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_291),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_295),
.B(n_290),
.Y(n_304)
);

AOI31xp33_ASAP7_75t_L g313 ( 
.A1(n_304),
.A2(n_308),
.A3(n_310),
.B(n_15),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_302),
.B(n_303),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_309),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_286),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_11),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_307),
.C(n_311),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_307),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_15),
.B(n_1),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_1),
.B(n_2),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_2),
.Y(n_319)
);


endmodule