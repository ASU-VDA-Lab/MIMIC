module fake_jpeg_1659_n_495 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_495);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_495;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_9),
.B(n_11),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_50),
.Y(n_139)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_51),
.Y(n_136)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_63),
.Y(n_108)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_59),
.Y(n_149)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_7),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_8),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_34),
.Y(n_113)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_95),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_91),
.Y(n_123)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_92),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_8),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_102),
.Y(n_134)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_19),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_105),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_23),
.C(n_25),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_11),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_70),
.B(n_23),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_57),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_143),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_93),
.A2(n_32),
.B1(n_25),
.B2(n_40),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_142),
.A2(n_146),
.B1(n_39),
.B2(n_22),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_92),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_72),
.A2(n_46),
.B1(n_31),
.B2(n_36),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_76),
.B(n_32),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_161),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_71),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_46),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_40),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_162),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_35),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_45),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_168),
.Y(n_220)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_170),
.Y(n_233)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_94),
.B1(n_86),
.B2(n_77),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_126),
.B1(n_131),
.B2(n_125),
.Y(n_210)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_14),
.B1(n_15),
.B2(n_26),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_SL g244 ( 
.A1(n_174),
.A2(n_206),
.B(n_208),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_118),
.A2(n_80),
.B1(n_78),
.B2(n_73),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_178),
.A2(n_131),
.B1(n_129),
.B2(n_152),
.Y(n_222)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_184),
.Y(n_215)
);

CKINVDCx12_ASAP7_75t_R g181 ( 
.A(n_105),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_35),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_195),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_108),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_197),
.Y(n_219)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_114),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_124),
.A2(n_56),
.B1(n_68),
.B2(n_65),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_194),
.B1(n_155),
.B2(n_125),
.Y(n_213)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_49),
.B1(n_58),
.B2(n_62),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_39),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_72),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_110),
.C(n_106),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_103),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_199),
.B(n_204),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_201),
.Y(n_230)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_207),
.Y(n_224)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_144),
.B(n_14),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_132),
.A2(n_15),
.B1(n_45),
.B2(n_34),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_117),
.Y(n_207)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_116),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_128),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_210),
.A2(n_198),
.B1(n_201),
.B2(n_179),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_213),
.A2(n_222),
.B1(n_225),
.B2(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_216),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_155),
.B1(n_137),
.B2(n_152),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_163),
.B(n_157),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_232),
.B(n_177),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_194),
.A2(n_137),
.B1(n_129),
.B2(n_160),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_130),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_164),
.B(n_153),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_178),
.A2(n_160),
.B1(n_145),
.B2(n_159),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_213),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_246),
.B(n_258),
.Y(n_291)
);

INVx4_ASAP7_75t_SL g247 ( 
.A(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_247),
.Y(n_279)
);

NOR4xp25_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_168),
.C(n_176),
.D(n_183),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_248),
.A2(n_269),
.B(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_185),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_254),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_215),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_252),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_238),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_182),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_215),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_256),
.B(n_259),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g258 ( 
.A(n_211),
.B(n_176),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_225),
.B1(n_239),
.B2(n_216),
.Y(n_280)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_262),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_228),
.B1(n_218),
.B2(n_193),
.Y(n_293)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_267),
.B(n_271),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_235),
.B(n_183),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_270),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_198),
.B(n_39),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_214),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_165),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_272),
.Y(n_276)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_221),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_222),
.B1(n_230),
.B2(n_240),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_274),
.A2(n_278),
.B1(n_293),
.B2(n_298),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_275),
.A2(n_277),
.B(n_285),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_269),
.A2(n_230),
.B(n_217),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_232),
.B1(n_241),
.B2(n_220),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_265),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_220),
.B1(n_211),
.B2(n_242),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_282),
.A2(n_295),
.B1(n_270),
.B2(n_267),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_233),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_284),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_224),
.B(n_228),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_233),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_302),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_260),
.A2(n_218),
.B1(n_234),
.B2(n_207),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_258),
.A2(n_226),
.B(n_237),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_296),
.A2(n_248),
.B(n_273),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_252),
.A2(n_234),
.B1(n_226),
.B2(n_212),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_253),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_247),
.Y(n_320)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_196),
.C(n_171),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_303),
.B(n_274),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_280),
.A2(n_251),
.B1(n_256),
.B2(n_254),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_321),
.B1(n_284),
.B2(n_278),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_246),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_320),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_290),
.Y(n_313)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_313),
.Y(n_345)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_315),
.A2(n_324),
.B(n_285),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_259),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_288),
.C(n_302),
.Y(n_337)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_317),
.A2(n_327),
.B1(n_279),
.B2(n_128),
.Y(n_348)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_247),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_322),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_263),
.B1(n_186),
.B2(n_212),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_295),
.B1(n_293),
.B2(n_318),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_276),
.A2(n_257),
.B1(n_236),
.B2(n_187),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_261),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_326),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_261),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_279),
.A2(n_202),
.B1(n_173),
.B2(n_209),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_223),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_328),
.B(n_331),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_189),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_294),
.Y(n_333)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_333),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_330),
.A2(n_296),
.B(n_291),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_336),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_321),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_300),
.Y(n_341)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_342),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_348),
.B1(n_359),
.B2(n_318),
.Y(n_363)
);

XNOR2x1_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_277),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_301),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_351),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_284),
.Y(n_350)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_308),
.B(n_291),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_302),
.C(n_277),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_316),
.C(n_315),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_297),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_354),
.B(n_309),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_322),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_320),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_282),
.B(n_292),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_356),
.B(n_298),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_299),
.Y(n_357)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_313),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_362),
.Y(n_388)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_368),
.C(n_372),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_359),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_303),
.C(n_322),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_351),
.A2(n_323),
.B1(n_306),
.B2(n_324),
.Y(n_370)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_326),
.C(n_306),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_341),
.B1(n_339),
.B2(n_334),
.Y(n_374)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_347),
.A2(n_325),
.B1(n_331),
.B2(n_328),
.Y(n_376)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_376),
.Y(n_398)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_379),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_319),
.C(n_314),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_383),
.C(n_384),
.Y(n_407)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_381),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_347),
.A2(n_295),
.B1(n_293),
.B2(n_281),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_382),
.A2(n_342),
.B1(n_340),
.B2(n_355),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_332),
.B(n_281),
.C(n_166),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_166),
.C(n_169),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_334),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_385),
.B(n_375),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_376),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_378),
.A2(n_342),
.B1(n_345),
.B2(n_339),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_SL g417 ( 
.A(n_390),
.B(n_392),
.C(n_393),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_386),
.B(n_336),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_400),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_371),
.A2(n_350),
.B(n_345),
.C(n_340),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_373),
.A2(n_333),
.B1(n_357),
.B2(n_346),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_373),
.A2(n_335),
.B1(n_353),
.B2(n_338),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_395),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_377),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_408),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_365),
.B(n_335),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_372),
.B(n_353),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_405),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_317),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_360),
.Y(n_408)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_410),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_375),
.Y(n_411)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_406),
.B(n_366),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_419),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_371),
.Y(n_414)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_414),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_396),
.A2(n_369),
.B1(n_361),
.B2(n_364),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_415),
.A2(n_420),
.B1(n_423),
.B2(n_424),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_402),
.A2(n_361),
.B(n_364),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_418),
.A2(n_425),
.B1(n_428),
.B2(n_398),
.Y(n_431)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_396),
.A2(n_368),
.B1(n_380),
.B2(n_349),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_422),
.B(n_426),
.Y(n_446)
);

OAI321xp33_ASAP7_75t_L g423 ( 
.A1(n_399),
.A2(n_349),
.A3(n_358),
.B1(n_382),
.B2(n_360),
.C(n_383),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_388),
.A2(n_358),
.B1(n_384),
.B2(n_317),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_167),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_389),
.A2(n_203),
.B1(n_160),
.B2(n_159),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_407),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_398),
.B1(n_405),
.B2(n_394),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_425),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_429),
.B(n_442),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_394),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_430),
.B(n_434),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_436),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_408),
.Y(n_434)
);

AO21x1_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_395),
.B(n_391),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_407),
.C(n_400),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_SL g451 ( 
.A(n_437),
.B(n_439),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_421),
.B(n_401),
.C(n_145),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_133),
.C(n_22),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_443),
.C(n_444),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_411),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_133),
.C(n_22),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_410),
.C(n_417),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_437),
.B(n_414),
.C(n_427),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_454),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_34),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_440),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_441),
.A2(n_26),
.B1(n_15),
.B2(n_45),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_458),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_36),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_26),
.C(n_138),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_457),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_138),
.C(n_135),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_432),
.A2(n_138),
.B(n_135),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_436),
.B(n_13),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_459),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_446),
.A2(n_135),
.B(n_105),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_460),
.A2(n_128),
.B1(n_46),
.B2(n_36),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_433),
.B1(n_445),
.B2(n_443),
.Y(n_462)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_463),
.Y(n_481)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_469),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_468),
.B(n_472),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_10),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_461),
.A2(n_149),
.B1(n_10),
.B2(n_13),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_12),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_6),
.Y(n_472)
);

OAI21xp33_ASAP7_75t_L g473 ( 
.A1(n_449),
.A2(n_6),
.B(n_12),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_473),
.A2(n_450),
.B(n_447),
.Y(n_474)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_474),
.Y(n_485)
);

AOI322xp5_ASAP7_75t_L g476 ( 
.A1(n_466),
.A2(n_451),
.A3(n_457),
.B1(n_455),
.B2(n_156),
.C1(n_6),
.C2(n_10),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_479),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_462),
.A2(n_467),
.B(n_473),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_477),
.B(n_464),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_481),
.B(n_470),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_484),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_464),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_0),
.Y(n_489)
);

AOI322xp5_ASAP7_75t_L g488 ( 
.A1(n_485),
.A2(n_480),
.A3(n_478),
.B1(n_156),
.B2(n_12),
.C1(n_3),
.C2(n_2),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_488),
.B(n_483),
.Y(n_490)
);

OAI211xp5_ASAP7_75t_L g491 ( 
.A1(n_489),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_490),
.A2(n_491),
.B(n_487),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_492),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_493),
.A2(n_1),
.B(n_3),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_1),
.Y(n_495)
);


endmodule