module real_aes_7440_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g534 ( .A1(n_0), .A2(n_180), .B(n_535), .C(n_538), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_1), .B(n_485), .Y(n_539) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g124 ( .A(n_2), .Y(n_124) );
INVx1_ASAP7_75t_L g192 ( .A(n_3), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_4), .B(n_152), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_5), .A2(n_458), .B(n_479), .Y(n_478) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_6), .A2(n_172), .B(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_7), .A2(n_35), .B1(n_146), .B2(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_8), .B(n_172), .Y(n_181) );
AND2x6_ASAP7_75t_L g164 ( .A(n_9), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_10), .A2(n_164), .B(n_463), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_11), .B(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_11), .B(n_36), .Y(n_125) );
INVx1_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
INVx1_ASAP7_75t_L g185 ( .A(n_13), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_14), .B(n_150), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_15), .B(n_152), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_16), .B(n_138), .Y(n_256) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_17), .A2(n_137), .A3(n_163), .B1(n_172), .B2(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_18), .B(n_146), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_19), .B(n_138), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_20), .A2(n_50), .B1(n_146), .B2(n_201), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_21), .A2(n_78), .B1(n_146), .B2(n_150), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_22), .B(n_146), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_23), .A2(n_163), .B(n_463), .C(n_512), .Y(n_511) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_24), .A2(n_55), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_24), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_25), .A2(n_163), .B(n_463), .C(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_26), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_27), .B(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_28), .A2(n_458), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_29), .B(n_167), .Y(n_215) );
INVx2_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_31), .A2(n_461), .B(n_471), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_32), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_33), .B(n_167), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_34), .B(n_222), .Y(n_492) );
INVx1_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_37), .B(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_38), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_39), .B(n_152), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_40), .B(n_458), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_41), .A2(n_461), .B(n_465), .C(n_471), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_42), .B(n_146), .Y(n_175) );
INVx1_ASAP7_75t_L g536 ( .A(n_43), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_44), .A2(n_89), .B1(n_201), .B2(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g466 ( .A(n_45), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_46), .B(n_146), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_47), .B(n_146), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_48), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_49), .B(n_158), .Y(n_179) );
AOI22xp33_ASAP7_75t_SL g254 ( .A1(n_51), .A2(n_56), .B1(n_146), .B2(n_150), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_52), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_53), .B(n_146), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_54), .B(n_146), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_55), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_55), .A2(n_129), .B1(n_130), .B2(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_57), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g165 ( .A(n_58), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_59), .B(n_458), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_60), .B(n_485), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_61), .A2(n_158), .B(n_188), .C(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_62), .B(n_146), .Y(n_193) );
INVx1_ASAP7_75t_L g141 ( .A(n_63), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_65), .B(n_152), .Y(n_503) );
AO32x2_ASAP7_75t_L g236 ( .A1(n_66), .A2(n_163), .A3(n_172), .B1(n_237), .B2(n_241), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_67), .B(n_153), .Y(n_549) );
INVx1_ASAP7_75t_L g156 ( .A(n_68), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_69), .A2(n_101), .B1(n_112), .B2(n_756), .Y(n_100) );
INVx1_ASAP7_75t_L g210 ( .A(n_70), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_71), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_72), .B(n_468), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_73), .A2(n_463), .B(n_471), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_74), .B(n_150), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_75), .Y(n_480) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_77), .B(n_467), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_79), .A2(n_83), .B1(n_442), .B2(n_749), .C1(n_754), .C2(n_755), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_80), .B(n_201), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_81), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_82), .B(n_150), .Y(n_214) );
INVx1_ASAP7_75t_L g754 ( .A(n_83), .Y(n_754) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_85), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_86), .B(n_162), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_87), .B(n_150), .Y(n_176) );
INVx2_ASAP7_75t_L g108 ( .A(n_88), .Y(n_108) );
OR2x2_ASAP7_75t_L g121 ( .A(n_88), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g445 ( .A(n_88), .B(n_123), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_90), .A2(n_99), .B1(n_150), .B2(n_151), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_91), .B(n_458), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_92), .Y(n_502) );
INVxp67_ASAP7_75t_L g483 ( .A(n_93), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_94), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_95), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g524 ( .A(n_96), .Y(n_524) );
INVx1_ASAP7_75t_L g545 ( .A(n_97), .Y(n_545) );
AND2x2_ASAP7_75t_L g473 ( .A(n_98), .B(n_167), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx12_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g757 ( .A(n_104), .Y(n_757) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
OR2x2_ASAP7_75t_L g450 ( .A(n_108), .B(n_123), .Y(n_450) );
NOR2x2_ASAP7_75t_L g755 ( .A(n_108), .B(n_122), .Y(n_755) );
OA211x2_ASAP7_75t_L g112 ( .A1(n_109), .A2(n_113), .B(n_118), .C(n_438), .Y(n_112) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g440 ( .A(n_115), .Y(n_440) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_126), .B(n_434), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g437 ( .A(n_121), .Y(n_437) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_130), .Y(n_126) );
INVx1_ASAP7_75t_SL g447 ( .A(n_130), .Y(n_447) );
OR3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_362), .C(n_411), .Y(n_130) );
NAND5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_277), .C(n_305), .D(n_335), .E(n_349), .Y(n_131) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_195), .B1(n_227), .B2(n_232), .C(n_243), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_168), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_134), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g257 ( .A(n_135), .Y(n_257) );
AND2x2_ASAP7_75t_L g265 ( .A(n_135), .B(n_171), .Y(n_265) );
AND2x2_ASAP7_75t_L g288 ( .A(n_135), .B(n_170), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_135), .B(n_182), .Y(n_303) );
OR2x2_ASAP7_75t_L g312 ( .A(n_135), .B(n_250), .Y(n_312) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_135), .Y(n_315) );
AND2x2_ASAP7_75t_L g423 ( .A(n_135), .B(n_250), .Y(n_423) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_166), .Y(n_135) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_136), .A2(n_183), .B(n_194), .Y(n_182) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_137), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_139), .B(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_155), .B(n_163), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B(n_152), .Y(n_144) );
INVx3_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_146), .Y(n_526) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
BUFx3_ASAP7_75t_L g239 ( .A(n_147), .Y(n_239) );
AND2x6_ASAP7_75t_L g463 ( .A(n_147), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
INVx1_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx2_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_152), .A2(n_175), .B(n_176), .Y(n_174) );
INVx2_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
O2A1O1Ixp5_ASAP7_75t_SL g208 ( .A1(n_152), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_152), .B(n_483), .Y(n_482) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g237 ( .A1(n_153), .A2(n_162), .B1(n_238), .B2(n_240), .Y(n_237) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
INVx1_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
AND2x2_ASAP7_75t_L g459 ( .A(n_154), .B(n_159), .Y(n_459) );
INVx1_ASAP7_75t_L g464 ( .A(n_154), .Y(n_464) );
O2A1O1Ixp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_160), .C(n_161), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_157), .A2(n_180), .B(n_192), .C(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_157), .A2(n_513), .B(n_514), .Y(n_512) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_161), .A2(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_162), .A2(n_180), .B1(n_200), .B2(n_202), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_162), .A2(n_180), .B1(n_253), .B2(n_254), .Y(n_252) );
INVx4_ASAP7_75t_L g537 ( .A(n_162), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g276 ( .A(n_163), .B(n_251), .C(n_252), .Y(n_276) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_164), .A2(n_174), .B(n_177), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_164), .A2(n_184), .B(n_191), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_164), .A2(n_208), .B(n_212), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_164), .A2(n_218), .B(n_223), .Y(n_217) );
AND2x4_ASAP7_75t_L g458 ( .A(n_164), .B(n_459), .Y(n_458) );
INVx4_ASAP7_75t_SL g472 ( .A(n_164), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_164), .B(n_459), .Y(n_546) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_167), .A2(n_207), .B(n_215), .Y(n_206) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_167), .A2(n_217), .B(n_226), .Y(n_216) );
INVx2_ASAP7_75t_L g241 ( .A(n_167), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_167), .A2(n_457), .B(n_460), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_167), .A2(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g518 ( .A(n_167), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_168), .B(n_315), .Y(n_371) );
INVx2_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
OAI311xp33_ASAP7_75t_L g313 ( .A1(n_169), .A2(n_314), .A3(n_315), .B1(n_316), .C1(n_331), .Y(n_313) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_182), .Y(n_169) );
AND2x2_ASAP7_75t_L g274 ( .A(n_170), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g281 ( .A(n_170), .Y(n_281) );
AND2x2_ASAP7_75t_L g402 ( .A(n_170), .B(n_231), .Y(n_402) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_171), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g258 ( .A(n_171), .B(n_182), .Y(n_258) );
AND2x2_ASAP7_75t_L g310 ( .A(n_171), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g324 ( .A(n_171), .B(n_257), .Y(n_324) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_181), .Y(n_171) );
INVx4_ASAP7_75t_L g251 ( .A(n_172), .Y(n_251) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_172), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_172), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_177) );
INVx2_ASAP7_75t_L g231 ( .A(n_182), .Y(n_231) );
AND2x2_ASAP7_75t_L g273 ( .A(n_182), .B(n_257), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_188), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_186), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_186), .A2(n_549), .B(n_550), .Y(n_548) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_188), .A2(n_524), .B(n_525), .C(n_526), .Y(n_523) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_189), .A2(n_213), .B(n_214), .Y(n_212) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g468 ( .A(n_190), .Y(n_468) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_203), .Y(n_195) );
OR2x2_ASAP7_75t_L g368 ( .A(n_196), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_196), .B(n_374), .Y(n_385) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_197), .B(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
AND2x2_ASAP7_75t_L g309 ( .A(n_198), .B(n_236), .Y(n_309) );
AND2x2_ASAP7_75t_L g320 ( .A(n_198), .B(n_216), .Y(n_320) );
AND2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_203), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_203), .B(n_270), .Y(n_314) );
INVx2_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g301 ( .A(n_204), .B(n_260), .Y(n_301) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_216), .Y(n_204) );
INVx2_ASAP7_75t_L g234 ( .A(n_205), .Y(n_234) );
AND2x2_ASAP7_75t_L g328 ( .A(n_205), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
OR2x2_ASAP7_75t_L g345 ( .A(n_206), .B(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_206), .Y(n_408) );
AND2x2_ASAP7_75t_L g247 ( .A(n_216), .B(n_242), .Y(n_247) );
INVx1_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
AND2x2_ASAP7_75t_L g289 ( .A(n_216), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g330 ( .A(n_216), .Y(n_330) );
INVx1_ASAP7_75t_L g346 ( .A(n_216), .Y(n_346) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_216), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVxp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_229), .B(n_334), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_229), .A2(n_319), .B1(n_368), .B2(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_230), .A2(n_412), .B(n_414), .C(n_432), .Y(n_411) );
INVx2_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
AND2x2_ASAP7_75t_L g322 ( .A(n_231), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g333 ( .A(n_231), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_232), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AND2x2_ASAP7_75t_L g306 ( .A(n_233), .B(n_270), .Y(n_306) );
BUFx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g338 ( .A(n_234), .B(n_329), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_234), .B(n_271), .Y(n_357) );
AND2x4_ASAP7_75t_L g293 ( .A(n_235), .B(n_267), .Y(n_293) );
AND2x2_ASAP7_75t_L g431 ( .A(n_235), .B(n_407), .Y(n_431) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_242), .Y(n_235) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx1_ASAP7_75t_L g271 ( .A(n_236), .Y(n_271) );
INVx1_ASAP7_75t_L g370 ( .A(n_236), .Y(n_370) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_239), .Y(n_470) );
INVx2_ASAP7_75t_L g538 ( .A(n_239), .Y(n_538) );
INVx1_ASAP7_75t_L g515 ( .A(n_241), .Y(n_515) );
OR2x2_ASAP7_75t_L g261 ( .A(n_242), .B(n_246), .Y(n_261) );
AND2x2_ASAP7_75t_L g270 ( .A(n_242), .B(n_271), .Y(n_270) );
NOR2xp67_ASAP7_75t_L g290 ( .A(n_242), .B(n_291), .Y(n_290) );
OAI221xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_248), .B1(n_259), .B2(n_262), .C(n_266), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_245), .A2(n_267), .B(n_269), .C(n_272), .Y(n_266) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_246), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_246), .B(n_268), .Y(n_374) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_246), .Y(n_381) );
AND2x2_ASAP7_75t_L g299 ( .A(n_247), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g336 ( .A(n_247), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_258), .Y(n_248) );
INVx2_ASAP7_75t_L g327 ( .A(n_249), .Y(n_327) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_249), .A2(n_260), .B1(n_377), .B2(n_379), .C1(n_380), .C2(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g433 ( .A(n_249), .B(n_402), .Y(n_433) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_257), .Y(n_249) );
INVx1_ASAP7_75t_L g323 ( .A(n_250), .Y(n_323) );
AO21x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_255), .Y(n_250) );
INVx3_ASAP7_75t_L g485 ( .A(n_251), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_251), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_251), .A2(n_521), .B(n_528), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_251), .B(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_251), .A2(n_544), .B(n_551), .Y(n_543) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g275 ( .A(n_256), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g361 ( .A(n_258), .B(n_295), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g372 ( .A1(n_259), .A2(n_373), .B(n_375), .Y(n_372) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g300 ( .A(n_260), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_260), .B(n_267), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_260), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx3_ASAP7_75t_L g326 ( .A(n_264), .Y(n_326) );
OR2x2_ASAP7_75t_L g378 ( .A(n_264), .B(n_300), .Y(n_378) );
AND2x2_ASAP7_75t_L g294 ( .A(n_265), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g332 ( .A(n_265), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_265), .B(n_326), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_265), .B(n_322), .Y(n_348) );
AND2x2_ASAP7_75t_L g352 ( .A(n_265), .B(n_334), .Y(n_352) );
INVxp67_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_269), .A2(n_342), .B1(n_347), .B2(n_348), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_269), .B(n_374), .Y(n_404) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g390 ( .A(n_270), .B(n_381), .Y(n_390) );
AND2x2_ASAP7_75t_L g419 ( .A(n_270), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g424 ( .A(n_270), .B(n_374), .Y(n_424) );
INVx1_ASAP7_75t_L g337 ( .A(n_271), .Y(n_337) );
BUFx2_ASAP7_75t_L g343 ( .A(n_271), .Y(n_343) );
INVx1_ASAP7_75t_L g428 ( .A(n_272), .Y(n_428) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_273), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
NOR2x1_ASAP7_75t_L g280 ( .A(n_275), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g287 ( .A(n_275), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
INVx3_ASAP7_75t_L g334 ( .A(n_275), .Y(n_334) );
OR2x2_ASAP7_75t_L g400 ( .A(n_275), .B(n_401), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_282), .B(n_285), .C(n_297), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_278), .A2(n_415), .B1(n_422), .B2(n_424), .C(n_425), .Y(n_414) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_286), .B(n_292), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_288), .B(n_326), .Y(n_340) );
AND2x2_ASAP7_75t_L g382 ( .A(n_288), .B(n_322), .Y(n_382) );
INVx1_ASAP7_75t_SL g395 ( .A(n_289), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_289), .B(n_343), .Y(n_398) );
INVx1_ASAP7_75t_L g416 ( .A(n_290), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_294), .A2(n_384), .B1(n_386), .B2(n_390), .C(n_391), .Y(n_383) );
AND2x2_ASAP7_75t_L g410 ( .A(n_295), .B(n_402), .Y(n_410) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g394 ( .A(n_296), .Y(n_394) );
AOI21xp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_301), .B(n_302), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g365 ( .A(n_300), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
INVx1_ASAP7_75t_L g379 ( .A(n_302), .Y(n_379) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_310), .C(n_313), .Y(n_305) );
OAI31xp33_ASAP7_75t_L g432 ( .A1(n_306), .A2(n_344), .A3(n_431), .B(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g406 ( .A(n_309), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g427 ( .A(n_309), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_311), .B(n_326), .Y(n_354) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g429 ( .A(n_312), .B(n_326), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_321), .B1(n_325), .B2(n_328), .Y(n_316) );
NAND2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_320), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g359 ( .A(n_320), .B(n_343), .Y(n_359) );
AND2x2_ASAP7_75t_L g413 ( .A(n_320), .B(n_408), .Y(n_413) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
NOR2xp67_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OAI32xp33_ASAP7_75t_L g391 ( .A1(n_326), .A2(n_360), .A3(n_392), .B1(n_394), .B2(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_329), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g389 ( .A(n_333), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B(n_339), .C(n_341), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_337), .B(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_338), .A2(n_350), .B1(n_351), .B2(n_352), .C(n_353), .Y(n_349) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g350 ( .A(n_348), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_358), .B2(n_360), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND4xp25_ASAP7_75t_SL g415 ( .A(n_358), .B(n_416), .C(n_417), .D(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NAND4xp25_ASAP7_75t_SL g362 ( .A(n_363), .B(n_376), .C(n_383), .D(n_396), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B(n_371), .C(n_372), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g393 ( .A(n_369), .Y(n_393) );
INVx2_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
OR2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B(n_403), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g422 ( .A(n_402), .B(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_405), .B(n_409), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B1(n_429), .B2(n_430), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND3xp33_ASAP7_75t_SL g438 ( .A(n_434), .B(n_439), .C(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B1(n_448), .B2(n_451), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g750 ( .A(n_444), .Y(n_750) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g751 ( .A(n_446), .Y(n_751) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g752 ( .A(n_449), .Y(n_752) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx4_ASAP7_75t_L g753 ( .A(n_451), .Y(n_753) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR5x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_622), .C(n_700), .D(n_724), .E(n_741), .Y(n_452) );
OAI211xp5_ASAP7_75t_SL g453 ( .A1(n_454), .A2(n_494), .B(n_540), .C(n_599), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_474), .Y(n_454) );
AND2x2_ASAP7_75t_L g553 ( .A(n_455), .B(n_476), .Y(n_553) );
INVx5_ASAP7_75t_SL g581 ( .A(n_455), .Y(n_581) );
AND2x2_ASAP7_75t_L g617 ( .A(n_455), .B(n_602), .Y(n_617) );
OR2x2_ASAP7_75t_L g656 ( .A(n_455), .B(n_475), .Y(n_656) );
OR2x2_ASAP7_75t_L g687 ( .A(n_455), .B(n_578), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_455), .B(n_591), .Y(n_723) );
AND2x2_ASAP7_75t_L g735 ( .A(n_455), .B(n_578), .Y(n_735) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_473), .Y(n_455) );
BUFx2_ASAP7_75t_L g510 ( .A(n_458), .Y(n_510) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_462), .A2(n_472), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_462), .A2(n_472), .B(n_533), .C(n_534), .Y(n_532) );
INVx5_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_469), .C(n_470), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_467), .A2(n_470), .B(n_502), .C(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g734 ( .A(n_474), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g597 ( .A(n_475), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_476), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_476), .Y(n_590) );
INVx3_ASAP7_75t_L g605 ( .A(n_476), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_476), .B(n_486), .Y(n_629) );
OR2x2_ASAP7_75t_L g638 ( .A(n_476), .B(n_581), .Y(n_638) );
AND2x2_ASAP7_75t_L g642 ( .A(n_476), .B(n_602), .Y(n_642) );
AND2x2_ASAP7_75t_L g648 ( .A(n_476), .B(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_L g685 ( .A(n_476), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_476), .B(n_543), .Y(n_699) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_484), .Y(n_476) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_485), .A2(n_531), .B(n_539), .Y(n_530) );
OR2x2_ASAP7_75t_L g591 ( .A(n_486), .B(n_543), .Y(n_591) );
AND2x2_ASAP7_75t_L g602 ( .A(n_486), .B(n_578), .Y(n_602) );
AND2x2_ASAP7_75t_L g614 ( .A(n_486), .B(n_605), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_486), .B(n_543), .Y(n_637) );
INVx1_ASAP7_75t_SL g649 ( .A(n_486), .Y(n_649) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g542 ( .A(n_487), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_487), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
AND2x2_ASAP7_75t_L g562 ( .A(n_496), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_496), .B(n_519), .Y(n_566) );
AND2x2_ASAP7_75t_L g569 ( .A(n_496), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_496), .B(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g594 ( .A(n_496), .B(n_585), .Y(n_594) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_496), .Y(n_613) );
AND2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g644 ( .A(n_496), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g690 ( .A(n_496), .B(n_573), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_496), .B(n_596), .Y(n_717) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g587 ( .A(n_497), .Y(n_587) );
AND2x2_ASAP7_75t_L g653 ( .A(n_497), .B(n_585), .Y(n_653) );
AND2x2_ASAP7_75t_L g737 ( .A(n_497), .B(n_605), .Y(n_737) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_506), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_506), .Y(n_726) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_519), .Y(n_506) );
AND2x2_ASAP7_75t_L g556 ( .A(n_507), .B(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g565 ( .A(n_507), .B(n_563), .Y(n_565) );
INVx5_ASAP7_75t_L g573 ( .A(n_507), .Y(n_573) );
AND2x2_ASAP7_75t_L g596 ( .A(n_507), .B(n_530), .Y(n_596) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_507), .Y(n_633) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
AOI21xp5_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_511), .B(n_515), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g674 ( .A(n_519), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_519), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g707 ( .A(n_519), .B(n_573), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_519), .A2(n_630), .B(n_737), .C(n_738), .Y(n_736) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_530), .Y(n_519) );
BUFx2_ASAP7_75t_L g557 ( .A(n_520), .Y(n_557) );
INVx2_ASAP7_75t_L g561 ( .A(n_520), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
INVx2_ASAP7_75t_L g563 ( .A(n_530), .Y(n_563) );
AND2x2_ASAP7_75t_L g570 ( .A(n_530), .B(n_561), .Y(n_570) );
AND2x2_ASAP7_75t_L g661 ( .A(n_530), .B(n_573), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AOI211x1_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_554), .B(n_567), .C(n_592), .Y(n_540) );
INVx1_ASAP7_75t_L g658 ( .A(n_541), .Y(n_658) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_553), .Y(n_541) );
INVx5_ASAP7_75t_SL g578 ( .A(n_543), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_543), .B(n_648), .Y(n_647) );
AOI311xp33_ASAP7_75t_L g666 ( .A1(n_543), .A2(n_667), .A3(n_669), .B(n_670), .C(n_676), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_543), .A2(n_614), .B(n_702), .C(n_705), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B(n_547), .Y(n_544) );
INVxp67_ASAP7_75t_L g621 ( .A(n_553), .Y(n_621) );
NAND4xp25_ASAP7_75t_SL g554 ( .A(n_555), .B(n_558), .C(n_564), .D(n_566), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_555), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g612 ( .A(n_556), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_559), .B(n_565), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_559), .B(n_572), .Y(n_692) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_560), .B(n_573), .Y(n_710) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g585 ( .A(n_561), .Y(n_585) );
INVxp67_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
AND2x4_ASAP7_75t_L g572 ( .A(n_563), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g646 ( .A(n_563), .B(n_585), .Y(n_646) );
INVx1_ASAP7_75t_L g673 ( .A(n_563), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_563), .B(n_660), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_564), .B(n_634), .Y(n_654) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_565), .B(n_587), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_565), .B(n_634), .Y(n_733) );
INVx1_ASAP7_75t_L g744 ( .A(n_566), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_571), .B(n_574), .C(n_582), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g586 ( .A(n_570), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g624 ( .A(n_570), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g606 ( .A(n_571), .Y(n_606) );
AND2x2_ASAP7_75t_L g583 ( .A(n_572), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_572), .B(n_634), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_572), .B(n_653), .Y(n_677) );
OR2x2_ASAP7_75t_L g593 ( .A(n_573), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g625 ( .A(n_573), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_573), .B(n_585), .Y(n_640) );
AND2x2_ASAP7_75t_L g697 ( .A(n_573), .B(n_653), .Y(n_697) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_573), .Y(n_704) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_575), .A2(n_587), .B1(n_709), .B2(n_711), .C(n_714), .Y(n_708) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g598 ( .A(n_578), .B(n_581), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_578), .B(n_648), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_578), .B(n_605), .Y(n_713) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g698 ( .A(n_580), .B(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g712 ( .A(n_580), .B(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_581), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g609 ( .A(n_581), .B(n_602), .Y(n_609) );
AND2x2_ASAP7_75t_L g679 ( .A(n_581), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_581), .B(n_628), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_581), .B(n_729), .Y(n_728) );
OAI21xp5_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_586), .B(n_588), .Y(n_582) );
INVx2_ASAP7_75t_L g615 ( .A(n_583), .Y(n_615) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g635 ( .A(n_585), .Y(n_635) );
OR2x2_ASAP7_75t_L g639 ( .A(n_587), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g742 ( .A(n_587), .B(n_710), .Y(n_742) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AOI21xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_595), .B(n_597), .Y(n_592) );
INVx1_ASAP7_75t_L g746 ( .A(n_593), .Y(n_746) );
INVx2_ASAP7_75t_SL g660 ( .A(n_594), .Y(n_660) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_597), .A2(n_678), .B(n_742), .C(n_743), .Y(n_741) );
OAI322xp33_ASAP7_75t_SL g610 ( .A1(n_598), .A2(n_611), .A3(n_614), .B1(n_615), .B2(n_616), .C1(n_618), .C2(n_621), .Y(n_610) );
INVx2_ASAP7_75t_L g630 ( .A(n_598), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_606), .B1(n_607), .B2(n_609), .C(n_610), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp33_ASAP7_75t_SL g676 ( .A1(n_601), .A2(n_677), .B1(n_678), .B2(n_681), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_602), .B(n_605), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_602), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g675 ( .A(n_604), .B(n_637), .Y(n_675) );
INVx1_ASAP7_75t_L g665 ( .A(n_605), .Y(n_665) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_609), .A2(n_719), .B(n_721), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g643 ( .A1(n_611), .A2(n_644), .B(n_647), .Y(n_643) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR2xp67_ASAP7_75t_SL g672 ( .A(n_613), .B(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_613), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g729 ( .A(n_614), .Y(n_729) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_623), .B(n_650), .C(n_666), .D(n_682), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B(n_631), .C(n_643), .Y(n_623) );
INVx1_ASAP7_75t_L g715 ( .A(n_624), .Y(n_715) );
AND2x2_ASAP7_75t_L g663 ( .A(n_625), .B(n_646), .Y(n_663) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_630), .B(n_665), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_636), .B1(n_639), .B2(n_641), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_633), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g681 ( .A(n_634), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g695 ( .A1(n_634), .A2(n_673), .B(n_696), .C(n_698), .Y(n_695) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g680 ( .A(n_637), .Y(n_680) );
INVx1_ASAP7_75t_L g740 ( .A(n_638), .Y(n_740) );
NAND2xp33_ASAP7_75t_SL g730 ( .A(n_639), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g669 ( .A(n_648), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_654), .B(n_655), .C(n_657), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_662), .B2(n_664), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_660), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_665), .B(n_686), .Y(n_748) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI21xp33_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_674), .B(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_688), .B1(n_691), .B2(n_693), .C(n_695), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_698), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
NAND3xp33_ASAP7_75t_SL g700 ( .A(n_701), .B(n_708), .C(n_718), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
CKINVDCx16_ASAP7_75t_R g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI211xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_727), .C(n_736), .Y(n_724) );
INVx1_ASAP7_75t_L g745 ( .A(n_725), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B1(n_732), .B2(n_734), .Y(n_727) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_743) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22x1_ASAP7_75t_SL g749 ( .A1(n_750), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
endmodule