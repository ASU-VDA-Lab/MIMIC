module fake_jpeg_30497_n_441 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_441);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_52),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_54),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_34),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_70),
.Y(n_90)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_76),
.Y(n_130)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_98),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_56),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_26),
.B1(n_37),
.B2(n_29),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_112),
.A2(n_37),
.B1(n_30),
.B2(n_36),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_44),
.A2(n_21),
.B(n_22),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_60),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_44),
.B(n_38),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_59),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_71),
.B1(n_74),
.B2(n_78),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_138),
.A2(n_153),
.B1(n_161),
.B2(n_163),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_77),
.B1(n_72),
.B2(n_49),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_53),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_162),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_87),
.B(n_30),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_149),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_147),
.B(n_95),
.CI(n_50),
.CON(n_191),
.SN(n_191)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_31),
.B1(n_105),
.B2(n_109),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_93),
.C(n_88),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_97),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_22),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_101),
.A2(n_32),
.B1(n_56),
.B2(n_47),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_123),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_159),
.B(n_164),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_100),
.B(n_36),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_32),
.B1(n_47),
.B2(n_21),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_32),
.B1(n_21),
.B2(n_73),
.Y(n_164)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_90),
.B(n_32),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_168),
.Y(n_188)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_169),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_117),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_191),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_94),
.C(n_99),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_140),
.C(n_143),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_100),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_91),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_132),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_161),
.Y(n_203)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_148),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_200),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_138),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_202),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_138),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_205),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_190),
.B(n_149),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_188),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_209),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_210),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_157),
.B(n_150),
.C(n_137),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_171),
.B(n_180),
.C(n_196),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_192),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_134),
.B1(n_140),
.B2(n_126),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_171),
.B1(n_184),
.B2(n_191),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_179),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_142),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_220),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_135),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_175),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_198),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_200),
.B1(n_217),
.B2(n_198),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_210),
.B1(n_209),
.B2(n_203),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_237),
.B1(n_238),
.B2(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_243),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_169),
.B1(n_191),
.B2(n_197),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_168),
.B1(n_132),
.B2(n_165),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_250),
.B1(n_229),
.B2(n_230),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_202),
.B1(n_213),
.B2(n_201),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_245),
.A2(n_90),
.B1(n_107),
.B2(n_182),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_254),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_218),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_252),
.C(n_248),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_218),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_248),
.B(n_255),
.Y(n_299)
);

CKINVDCx10_ASAP7_75t_R g249 ( 
.A(n_233),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_232),
.A2(n_182),
.B1(n_208),
.B2(n_178),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_233),
.B1(n_236),
.B2(n_223),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_221),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_200),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_219),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_226),
.C(n_178),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_204),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_146),
.Y(n_296)
);

XOR2x1_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_234),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_265),
.B(n_223),
.Y(n_280)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_227),
.Y(n_264)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_228),
.A2(n_237),
.B(n_234),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_240),
.B(n_220),
.Y(n_266)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_189),
.B(n_14),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_214),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_268),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_206),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_199),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_236),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_270),
.A2(n_96),
.B1(n_102),
.B2(n_130),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_265),
.B(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_271),
.B(n_273),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_268),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_127),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_238),
.B1(n_242),
.B2(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_284),
.B1(n_286),
.B2(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_257),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_249),
.A2(n_226),
.B1(n_224),
.B2(n_197),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_264),
.B1(n_260),
.B2(n_253),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_291),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_196),
.C(n_181),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_289),
.C(n_292),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_224),
.B1(n_186),
.B2(n_177),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_187),
.B1(n_195),
.B2(n_194),
.Y(n_286)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_133),
.C(n_145),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_195),
.B1(n_194),
.B2(n_152),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_144),
.B1(n_166),
.B2(n_160),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_107),
.C(n_156),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_92),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_296),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_269),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_311),
.Y(n_348)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_312),
.B1(n_316),
.B2(n_320),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_272),
.B(n_253),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_322),
.Y(n_341)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_257),
.C(n_155),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_314),
.C(n_289),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_127),
.C(n_130),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_275),
.B(n_0),
.Y(n_318)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_318),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_294),
.A2(n_93),
.B1(n_88),
.B2(n_102),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_279),
.B(n_10),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_324),
.B(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_299),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_326),
.B(n_328),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_299),
.C(n_292),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_335),
.C(n_339),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_313),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_331),
.B(n_333),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_280),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_342),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_318),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_314),
.C(n_301),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_302),
.A2(n_287),
.B(n_285),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_336),
.A2(n_136),
.B(n_96),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_277),
.B1(n_291),
.B2(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_285),
.C(n_290),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_302),
.B(n_286),
.CI(n_287),
.CON(n_340),
.SN(n_340)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_304),
.A2(n_293),
.B1(n_166),
.B2(n_160),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_307),
.A2(n_293),
.B1(n_158),
.B2(n_154),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_343),
.A2(n_325),
.B1(n_324),
.B2(n_316),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_141),
.C(n_125),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_347),
.C(n_144),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_128),
.C(n_125),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_341),
.B(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_355),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_336),
.A2(n_303),
.B(n_315),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_363),
.B(n_115),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_306),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_369),
.B1(n_158),
.B2(n_128),
.Y(n_380)
);

BUFx12_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_12),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_358),
.B(n_328),
.Y(n_372)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_345),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_364),
.Y(n_382)
);

OA21x2_ASAP7_75t_SL g361 ( 
.A1(n_329),
.A2(n_335),
.B(n_326),
.Y(n_361)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_361),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_332),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_366),
.Y(n_379)
);

AO22x1_ASAP7_75t_L g363 ( 
.A1(n_340),
.A2(n_320),
.B1(n_312),
.B2(n_95),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_16),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_136),
.Y(n_366)
);

OAI22x1_ASAP7_75t_SL g369 ( 
.A1(n_337),
.A2(n_339),
.B1(n_350),
.B2(n_349),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_350),
.A2(n_327),
.B1(n_345),
.B2(n_330),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_0),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_118),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_380),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_347),
.C(n_343),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_373),
.B(n_376),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_353),
.A2(n_346),
.B(n_95),
.Y(n_374)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_353),
.A2(n_154),
.B(n_152),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_362),
.C(n_366),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_358),
.C(n_371),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_370),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_363),
.A2(n_83),
.B1(n_79),
.B2(n_62),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_383),
.A2(n_387),
.B1(n_354),
.B2(n_115),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_385),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_365),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_118),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_386),
.B(n_388),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_401),
.C(n_32),
.Y(n_409)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_400),
.Y(n_408)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_377),
.Y(n_396)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_396),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_357),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_398),
.B(n_399),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_378),
.C(n_375),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_357),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_61),
.C(n_48),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_379),
.C(n_386),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_402),
.B(n_409),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_387),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_0),
.Y(n_419)
);

OAI22xp33_ASAP7_75t_L g404 ( 
.A1(n_396),
.A2(n_383),
.B1(n_384),
.B2(n_10),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_412),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_397),
.A2(n_13),
.B(n_12),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_407),
.A2(n_1),
.B(n_3),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_21),
.C(n_27),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_413),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_13),
.C(n_11),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_391),
.A2(n_13),
.B1(n_11),
.B2(n_2),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_405),
.A2(n_392),
.B(n_394),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_415),
.A2(n_420),
.B(n_3),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_393),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_1),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_406),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_418),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_429)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_419),
.Y(n_427)
);

AOI21xp33_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_27),
.B(n_3),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_421),
.B(n_422),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_27),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g424 ( 
.A1(n_417),
.A2(n_404),
.B(n_402),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_426),
.B(n_414),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_410),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_428),
.B(n_429),
.Y(n_434)
);

OAI221xp5_ASAP7_75t_L g432 ( 
.A1(n_430),
.A2(n_419),
.B1(n_422),
.B2(n_6),
.C(n_7),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_432),
.Y(n_436)
);

AOI322xp5_ASAP7_75t_L g433 ( 
.A1(n_427),
.A2(n_21),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_9),
.C2(n_4),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_425),
.C(n_5),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_437),
.B(n_9),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_4),
.C(n_6),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_436),
.B(n_9),
.Y(n_439)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_439),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_9),
.Y(n_441)
);


endmodule