module fake_aes_458_n_28 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
NOR2xp33_ASAP7_75t_L g13 ( .A(n_6), .B(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_11), .B(n_4), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_0), .B(n_7), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_0), .B(n_1), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_17), .B(n_1), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_16), .B1(n_15), .B2(n_13), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
OAI21xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_19), .B(n_18), .Y(n_24) );
NOR4xp75_ASAP7_75t_L g25 ( .A(n_24), .B(n_2), .C(n_3), .D(n_13), .Y(n_25) );
OA22x2_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_2), .B1(n_5), .B2(n_9), .Y(n_26) );
OAI22xp5_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_18), .B1(n_10), .B2(n_12), .Y(n_27) );
OA21x2_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_18), .B(n_24), .Y(n_28) );
endmodule