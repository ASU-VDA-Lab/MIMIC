module fake_jpeg_16153_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_45),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_51),
.B1(n_60),
.B2(n_30),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_52),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_56),
.B1(n_19),
.B2(n_30),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_25),
.C(n_24),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_27),
.B1(n_18),
.B2(n_35),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_18),
.B1(n_31),
.B2(n_34),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_24),
.B1(n_25),
.B2(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_32),
.Y(n_58)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_21),
.B1(n_32),
.B2(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_45),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_21),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_22),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_69),
.A2(n_77),
.B1(n_83),
.B2(n_34),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_75),
.Y(n_102)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_36),
.B(n_38),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_82),
.B(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_21),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_17),
.B1(n_35),
.B2(n_34),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_38),
.B1(n_42),
.B2(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_54),
.B1(n_64),
.B2(n_45),
.Y(n_119)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_87),
.Y(n_113)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_52),
.A3(n_50),
.B1(n_58),
.B2(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_103),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_49),
.B1(n_51),
.B2(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_106),
.B1(n_114),
.B2(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_110),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_60),
.B1(n_62),
.B2(n_54),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_43),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_98),
.C(n_101),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_64),
.C(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_75),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_70),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_54),
.B1(n_53),
.B2(n_68),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_54),
.B1(n_53),
.B2(n_68),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_68),
.B(n_1),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_116),
.A2(n_72),
.B(n_31),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_86),
.B1(n_78),
.B2(n_96),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_120),
.B1(n_17),
.B2(n_111),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_70),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_71),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_126),
.B(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_85),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_128),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_125),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_74),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_119),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_98),
.A2(n_94),
.B(n_92),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_139),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_43),
.C(n_63),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_42),
.C(n_45),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_144),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_141),
.B1(n_153),
.B2(n_108),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_74),
.B1(n_78),
.B2(n_81),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_64),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_152),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_42),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_108),
.C(n_123),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_0),
.B(n_1),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_93),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_97),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_157),
.A2(n_160),
.B(n_164),
.Y(n_203)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_106),
.B1(n_116),
.B2(n_114),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g204 ( 
.A1(n_159),
.A2(n_140),
.B1(n_129),
.B2(n_150),
.Y(n_204)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_110),
.Y(n_160)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_113),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_170),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_169),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_186),
.Y(n_190)
);

OAI22x1_ASAP7_75t_SL g174 ( 
.A1(n_137),
.A2(n_25),
.B1(n_123),
.B2(n_29),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_178),
.B1(n_143),
.B2(n_142),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_117),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_176),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_117),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_146),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_182),
.B(n_183),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_137),
.B1(n_153),
.B2(n_134),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_133),
.C(n_139),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_10),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_147),
.B(n_10),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_123),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_3),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_109),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_172),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_191),
.B(n_198),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_131),
.B(n_128),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_206),
.B(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_134),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_194),
.C(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_147),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_136),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_199),
.A2(n_168),
.B1(n_185),
.B2(n_161),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_216),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_202),
.C(n_205),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_130),
.C(n_155),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_174),
.B1(n_184),
.B2(n_157),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_141),
.C(n_151),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_0),
.B(n_2),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_160),
.C(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_211),
.C(n_212),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_154),
.C(n_149),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_154),
.C(n_109),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_3),
.B(n_4),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_20),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_185),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_233),
.B1(n_215),
.B2(n_20),
.Y(n_257)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g220 ( 
.A(n_197),
.Y(n_220)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_222),
.B(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_186),
.C(n_182),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_231),
.Y(n_264)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_209),
.A2(n_204),
.B(n_180),
.C(n_158),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_192),
.B(n_199),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_203),
.A2(n_158),
.A3(n_156),
.B1(n_168),
.B2(n_179),
.C1(n_165),
.C2(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_177),
.B1(n_163),
.B2(n_161),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_163),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_210),
.B(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_203),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_183),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_196),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_201),
.B1(n_189),
.B2(n_194),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_193),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_226),
.C(n_243),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_246),
.C(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_227),
.C(n_241),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_232),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_234),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_252),
.C(n_223),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_189),
.C(n_211),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_254),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_210),
.B1(n_204),
.B2(n_206),
.Y(n_255)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_SL g259 ( 
.A(n_229),
.B(n_20),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_233),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_20),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_237),
.C(n_230),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_3),
.B(n_4),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_271),
.C(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_239),
.C(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_252),
.C(n_244),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_282),
.C(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_238),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_279),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_225),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_225),
.C(n_20),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_247),
.B1(n_254),
.B2(n_255),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_291),
.B1(n_290),
.B2(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_261),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_293),
.Y(n_298)
);

AOI22x1_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_253),
.B1(n_247),
.B2(n_257),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_264),
.B1(n_258),
.B2(n_265),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_R g293 ( 
.A(n_270),
.B(n_260),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_269),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_267),
.C(n_273),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_267),
.C(n_282),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_302),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_11),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_11),
.B(n_15),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_308),
.B(n_5),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_5),
.C(n_6),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_13),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_285),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_309),
.A3(n_292),
.B1(n_295),
.B2(n_283),
.C1(n_9),
.C2(n_13),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_288),
.B1(n_290),
.B2(n_293),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_9),
.C(n_14),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_299),
.C(n_304),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_9),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_302),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_311),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_16),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_322),
.C(n_324),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_323),
.B(n_325),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_314),
.B(n_6),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_312),
.C(n_325),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_318),
.C(n_328),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_326),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_7),
.B(n_327),
.Y(n_332)
);


endmodule