module fake_ariane_2803_n_1723 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1723);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1723;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_0),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_12),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_98),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_57),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_71),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_70),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_40),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_111),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_75),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_31),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_34),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_97),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_51),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_77),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_3),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_17),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_135),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_95),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_16),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_81),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_61),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_82),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_85),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_126),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_7),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_49),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

HB1xp67_ASAP7_75t_SL g192 ( 
.A(n_145),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_39),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_45),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_22),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_53),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_8),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_14),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_129),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_41),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_43),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_19),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_38),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_9),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_63),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_102),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_0),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_33),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_49),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_54),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_137),
.Y(n_216)
);

BUFx2_ASAP7_75t_SL g217 ( 
.A(n_108),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_30),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_93),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_34),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_64),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_106),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_90),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_60),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_40),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_36),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_29),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_31),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_5),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_88),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_44),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_148),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_3),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_22),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_86),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_55),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_117),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_73),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_136),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_103),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_153),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_27),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_58),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_11),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_96),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_14),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_69),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_125),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_79),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_41),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_94),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_118),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_62),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_147),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_35),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_87),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_23),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_65),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_51),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_140),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_76),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_123),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_107),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_134),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_45),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_24),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_42),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_149),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_83),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_151),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_19),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_50),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_48),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_48),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_110),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_113),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_42),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_124),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_74),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_91),
.Y(n_286)
);

BUFx2_ASAP7_75t_SL g287 ( 
.A(n_114),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_18),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_127),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_37),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_2),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_7),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_101),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_100),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_29),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_130),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_66),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_121),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_44),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_84),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_116),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_38),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_112),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_37),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_142),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_32),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_47),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_16),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_132),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_304),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_249),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_156),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_210),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_159),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_159),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_268),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_161),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_161),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_235),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_258),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_163),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_172),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_169),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_261),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_169),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_176),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_176),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_184),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_184),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_197),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_197),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_198),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_192),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_212),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_198),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_194),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_212),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_204),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_227),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_205),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_156),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_204),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_212),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_211),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_211),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_212),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_162),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_182),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_215),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_189),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_190),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_215),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_193),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_212),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_239),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_196),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_239),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_256),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_199),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_263),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_162),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_263),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_299),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_201),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_248),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_299),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_207),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_282),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_168),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_299),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_289),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_289),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_208),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_310),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_213),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_270),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

INVxp33_ASAP7_75t_SL g384 ( 
.A(n_311),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

NOR2x1_ASAP7_75t_L g386 ( 
.A(n_315),
.B(n_298),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_315),
.B(n_219),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_338),
.A2(n_369),
.B1(n_381),
.B2(n_295),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_316),
.B(n_219),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_321),
.A2(n_157),
.B1(n_179),
.B2(n_206),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_281),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_173),
.C(n_168),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_339),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_319),
.B(n_203),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_300),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_325),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_342),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_312),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_157),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_317),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_370),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_335),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_335),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_324),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_314),
.A2(n_220),
.B1(n_307),
.B2(n_292),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_328),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_329),
.B(n_247),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_330),
.B(n_331),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_330),
.B(n_331),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_332),
.B(n_203),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_314),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_341),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_333),
.B(n_179),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_334),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_352),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_334),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_340),
.Y(n_438)
);

BUFx8_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_346),
.B(n_300),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_380),
.B(n_247),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_347),
.B(n_186),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_347),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_351),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_387),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_358),
.C(n_355),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_397),
.B(n_322),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_407),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_407),
.Y(n_454)
);

BUFx6f_ASAP7_75t_SL g455 ( 
.A(n_392),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_427),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_322),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_395),
.B(n_368),
.C(n_362),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

AND3x4_ASAP7_75t_L g462 ( 
.A(n_392),
.B(n_252),
.C(n_214),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_401),
.B(n_326),
.Y(n_464)
);

OAI22x1_ASAP7_75t_L g465 ( 
.A1(n_395),
.A2(n_364),
.B1(n_343),
.B2(n_373),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_405),
.B(n_326),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_354),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

INVx8_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_392),
.B(n_313),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_392),
.B(n_371),
.Y(n_473)
);

AO21x2_ASAP7_75t_L g474 ( 
.A1(n_442),
.A2(n_357),
.B(n_354),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_429),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_206),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_411),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_415),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_389),
.A2(n_379),
.B1(n_353),
.B2(n_377),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_433),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_429),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_433),
.B(n_439),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_429),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_420),
.B(n_349),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_429),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_429),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_436),
.Y(n_489)
);

CKINVDCx6p67_ASAP7_75t_R g490 ( 
.A(n_427),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_436),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_444),
.A2(n_323),
.B1(n_228),
.B2(n_309),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_436),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_423),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_439),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_436),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_436),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_415),
.B(n_357),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_439),
.B(n_359),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_436),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_418),
.B(n_359),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_436),
.Y(n_503)
);

NAND3xp33_ASAP7_75t_L g504 ( 
.A(n_444),
.B(n_439),
.C(n_389),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_439),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_437),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_425),
.B(n_360),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_437),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_437),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_437),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_SL g514 ( 
.A(n_430),
.B(n_225),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_L g515 ( 
.A(n_437),
.B(n_299),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_447),
.Y(n_517)
);

BUFx6f_ASAP7_75t_SL g518 ( 
.A(n_412),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_447),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_418),
.B(n_360),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_447),
.B(n_247),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_447),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_447),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_447),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_442),
.A2(n_380),
.B1(n_378),
.B2(n_376),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_423),
.Y(n_526)
);

BUFx4f_ASAP7_75t_L g527 ( 
.A(n_447),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_413),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_403),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_425),
.B(n_361),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_425),
.B(n_389),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_425),
.B(n_361),
.Y(n_532)
);

BUFx8_ASAP7_75t_SL g533 ( 
.A(n_409),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_403),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_403),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_391),
.A2(n_280),
.B1(n_229),
.B2(n_230),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_403),
.B(n_247),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_424),
.B(n_365),
.C(n_363),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_409),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_383),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_387),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_403),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_408),
.B(n_247),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_408),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_384),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_408),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_404),
.B(n_363),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_388),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_408),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_384),
.Y(n_551)
);

NAND2xp33_ASAP7_75t_SL g552 ( 
.A(n_387),
.B(n_226),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_388),
.Y(n_553)
);

AO21x2_ASAP7_75t_L g554 ( 
.A1(n_432),
.A2(n_366),
.B(n_365),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_408),
.Y(n_555)
);

AOI21x1_ASAP7_75t_L g556 ( 
.A1(n_385),
.A2(n_372),
.B(n_366),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_388),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_425),
.B(n_372),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_393),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_424),
.B(n_416),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_393),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_421),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_406),
.B(n_375),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_393),
.Y(n_564)
);

AND3x2_ASAP7_75t_L g565 ( 
.A(n_412),
.B(n_175),
.C(n_173),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_417),
.Y(n_566)
);

BUFx6f_ASAP7_75t_SL g567 ( 
.A(n_412),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_404),
.B(n_375),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_406),
.B(n_376),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_385),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_421),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_406),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_398),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_406),
.B(n_378),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_421),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_412),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_398),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_421),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_421),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_412),
.B(n_232),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_431),
.B(n_214),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_394),
.Y(n_583)
);

INVx6_ASAP7_75t_L g584 ( 
.A(n_431),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_394),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_431),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_432),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_390),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_435),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_399),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_431),
.B(n_233),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_399),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_431),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_582),
.A2(n_400),
.B1(n_386),
.B2(n_435),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_531),
.B(n_402),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_L g596 ( 
.A(n_478),
.B(n_399),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_587),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_587),
.Y(n_598)
);

BUFx6f_ASAP7_75t_SL g599 ( 
.A(n_452),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_534),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_534),
.Y(n_601)
);

NOR2xp67_ASAP7_75t_L g602 ( 
.A(n_478),
.B(n_410),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_548),
.B(n_410),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_543),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_543),
.Y(n_605)
);

AO22x1_ASAP7_75t_L g606 ( 
.A1(n_462),
.A2(n_402),
.B1(n_426),
.B2(n_244),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_473),
.B(n_410),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_582),
.B(n_414),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_414),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_577),
.B(n_414),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_545),
.A2(n_446),
.B(n_445),
.C(n_441),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_545),
.A2(n_446),
.B(n_445),
.C(n_441),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_458),
.B(n_428),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_470),
.B(n_428),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_547),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_547),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_568),
.B(n_428),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_467),
.B(n_434),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_550),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_541),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_464),
.B(n_434),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_470),
.A2(n_446),
.B1(n_445),
.B2(n_441),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_550),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_467),
.B(n_434),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_468),
.B(n_438),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_468),
.B(n_438),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_470),
.B(n_586),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_480),
.B(n_438),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_466),
.B(n_440),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_542),
.B(n_402),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_455),
.A2(n_462),
.B1(n_470),
.B2(n_518),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_480),
.B(n_440),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_L g635 ( 
.A(n_459),
.B(n_440),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_450),
.B(n_400),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_527),
.A2(n_580),
.B(n_562),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_L g638 ( 
.A(n_449),
.B(n_386),
.C(n_246),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_560),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_586),
.B(n_267),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_472),
.B(n_426),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_593),
.B(n_426),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_593),
.B(n_390),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_593),
.B(n_498),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_580),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_541),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_472),
.B(n_390),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_472),
.B(n_390),
.Y(n_648)
);

OAI22xp33_ASAP7_75t_L g649 ( 
.A1(n_486),
.A2(n_252),
.B1(n_220),
.B2(n_272),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_474),
.B(n_390),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_495),
.B(n_298),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_560),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_455),
.A2(n_217),
.B1(n_287),
.B2(n_254),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_474),
.B(n_584),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_586),
.B(n_267),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_481),
.B(n_236),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_448),
.B(n_257),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_474),
.B(n_584),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_584),
.B(n_178),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_455),
.B(n_259),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_529),
.B(n_275),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_518),
.A2(n_217),
.B1(n_287),
.B2(n_253),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_528),
.B(n_158),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_457),
.B(n_391),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_566),
.Y(n_665)
);

NOR3xp33_ASAP7_75t_L g666 ( 
.A(n_546),
.B(n_200),
.C(n_272),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_584),
.B(n_178),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_566),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_529),
.B(n_275),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_529),
.B(n_195),
.Y(n_670)
);

AND2x6_ASAP7_75t_SL g671 ( 
.A(n_477),
.B(n_195),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_566),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_536),
.B(n_200),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_504),
.B(n_260),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_536),
.B(n_218),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_452),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_536),
.B(n_218),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_555),
.B(n_269),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_518),
.A2(n_188),
.B1(n_224),
.B2(n_223),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_555),
.B(n_262),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_573),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_555),
.B(n_269),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_572),
.B(n_292),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_572),
.B(n_307),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_572),
.B(n_271),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_549),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_576),
.B(n_160),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_482),
.B(n_280),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_576),
.B(n_164),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_576),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_579),
.B(n_581),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_579),
.B(n_276),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_579),
.B(n_277),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_494),
.B(n_278),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_459),
.B(n_165),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_486),
.A2(n_227),
.B1(n_245),
.B2(n_280),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_591),
.B(n_279),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_482),
.B(n_452),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_526),
.B(n_283),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_459),
.B(n_487),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_589),
.B(n_288),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_507),
.B(n_290),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_590),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_549),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_590),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_570),
.Y(n_706)
);

INVx8_ASAP7_75t_L g707 ( 
.A(n_567),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_459),
.B(n_166),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_459),
.B(n_167),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_553),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_477),
.B(n_394),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_482),
.B(n_291),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_487),
.B(n_496),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_553),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_530),
.B(n_302),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_557),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_532),
.B(n_306),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_558),
.B(n_308),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_495),
.B(n_394),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_487),
.B(n_170),
.Y(n_720)
);

NAND3xp33_ASAP7_75t_L g721 ( 
.A(n_460),
.B(n_486),
.C(n_528),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_486),
.B(n_174),
.C(n_171),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_557),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_573),
.B(n_227),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_487),
.B(n_496),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_487),
.B(n_177),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_525),
.A2(n_569),
.B(n_563),
.C(n_575),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_567),
.B(n_245),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_533),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_501),
.B(n_180),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_520),
.B(n_181),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_477),
.A2(n_245),
.B1(n_422),
.B2(n_443),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_574),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_546),
.B(n_1),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_552),
.B(n_297),
.C(n_251),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_492),
.A2(n_1),
.B(n_4),
.C(n_5),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_539),
.B(n_183),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_574),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_457),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_551),
.B(n_4),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_551),
.B(n_6),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_592),
.B(n_185),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_496),
.B(n_187),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_578),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_567),
.B(n_6),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_592),
.B(n_191),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_578),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_592),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_556),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_588),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_588),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_559),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_499),
.A2(n_443),
.B1(n_422),
.B2(n_396),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_496),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_496),
.B(n_505),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_505),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_559),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_561),
.Y(n_758)
);

AND2x4_ASAP7_75t_SL g759 ( 
.A(n_535),
.B(n_394),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_613),
.B(n_554),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_633),
.B(n_484),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_600),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_636),
.A2(n_465),
.B1(n_514),
.B2(n_537),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_729),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_707),
.B(n_465),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_636),
.A2(n_639),
.B1(n_652),
.B2(n_606),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_629),
.B(n_571),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_SL g768 ( 
.A(n_657),
.B(n_286),
.C(n_240),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_601),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_623),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_707),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_599),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_604),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_724),
.A2(n_554),
.B1(n_535),
.B2(n_490),
.Y(n_774)
);

INVx4_ASAP7_75t_L g775 ( 
.A(n_707),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_599),
.Y(n_776)
);

CKINVDCx6p67_ASAP7_75t_R g777 ( 
.A(n_676),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_698),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_605),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_739),
.B(n_664),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_613),
.B(n_554),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_621),
.B(n_500),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_596),
.B(n_535),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_595),
.A2(n_490),
.B1(n_561),
.B2(n_564),
.Y(n_784)
);

BUFx6f_ASAP7_75t_SL g785 ( 
.A(n_676),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_641),
.B(n_595),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_621),
.B(n_565),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_615),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_631),
.B(n_500),
.Y(n_789)
);

NOR2x2_ASAP7_75t_L g790 ( 
.A(n_711),
.B(n_540),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_722),
.B(n_540),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_616),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_631),
.B(n_500),
.Y(n_793)
);

BUFx5_ASAP7_75t_L g794 ( 
.A(n_619),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_595),
.B(n_510),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_644),
.A2(n_556),
.B1(n_519),
.B2(n_524),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_674),
.A2(n_564),
.B1(n_451),
.B2(n_469),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_681),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_SL g799 ( 
.A1(n_611),
.A2(n_502),
.B(n_453),
.C(n_454),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_681),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_603),
.B(n_617),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_665),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_754),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_629),
.B(n_571),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_754),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_624),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_632),
.B(n_510),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_711),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_734),
.Y(n_809)
);

AO22x1_ASAP7_75t_L g810 ( 
.A1(n_740),
.A2(n_571),
.B1(n_266),
.B2(n_294),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_602),
.B(n_510),
.Y(n_811)
);

INVx4_ASAP7_75t_L g812 ( 
.A(n_759),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_700),
.A2(n_527),
.B(n_454),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_626),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_668),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_721),
.B(n_519),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_645),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_672),
.B(n_651),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_741),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_642),
.B(n_453),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_607),
.A2(n_519),
.B(n_524),
.C(n_461),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_618),
.B(n_524),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_625),
.B(n_451),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_759),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_607),
.B(n_461),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_703),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_719),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_594),
.B(n_724),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_705),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_728),
.B(n_469),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_688),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_706),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_608),
.B(n_475),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_671),
.Y(n_834)
);

BUFx8_ASAP7_75t_L g835 ( 
.A(n_712),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_733),
.B(n_475),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_719),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_738),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_744),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_674),
.A2(n_503),
.B1(n_479),
.B2(n_485),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_728),
.B(n_476),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_747),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_666),
.B(n_538),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_749),
.A2(n_612),
.B(n_637),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_745),
.B(n_527),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_649),
.A2(n_456),
.B1(n_463),
.B2(n_471),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_597),
.Y(n_847)
);

INVx6_ASAP7_75t_L g848 ( 
.A(n_663),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_647),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_660),
.Y(n_850)
);

INVxp33_ASAP7_75t_SL g851 ( 
.A(n_679),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_680),
.B(n_693),
.Y(n_852)
);

AOI211xp5_ASAP7_75t_L g853 ( 
.A1(n_656),
.A2(n_544),
.B(n_538),
.C(n_515),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_648),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_660),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_745),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_654),
.A2(n_509),
.B1(n_479),
.B2(n_485),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_750),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_697),
.B(n_456),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_598),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_614),
.B(n_476),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_680),
.B(n_491),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_SL g863 ( 
.A(n_735),
.B(n_238),
.C(n_202),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_L g864 ( 
.A(n_691),
.B(n_544),
.C(n_471),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_691),
.A2(n_463),
.B1(n_483),
.B2(n_523),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_659),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_658),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_667),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_749),
.A2(n_489),
.B(n_483),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_690),
.B(n_491),
.Y(n_870)
);

BUFx8_ASAP7_75t_L g871 ( 
.A(n_751),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_627),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_702),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_693),
.A2(n_488),
.B1(n_489),
.B2(n_523),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_628),
.B(n_630),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_634),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_620),
.B(n_493),
.Y(n_877)
);

INVx5_ASAP7_75t_L g878 ( 
.A(n_646),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_646),
.B(n_493),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_686),
.B(n_503),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_715),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_686),
.B(n_506),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_697),
.B(n_488),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_704),
.B(n_710),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_696),
.A2(n_511),
.B1(n_509),
.B2(n_506),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_704),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_748),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_710),
.B(n_511),
.Y(n_888)
);

NAND2x1_ASAP7_75t_L g889 ( 
.A(n_752),
.B(n_497),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_757),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_662),
.B(n_583),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_614),
.A2(n_497),
.B1(n_502),
.B2(n_522),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_714),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_670),
.Y(n_894)
);

OR2x6_ASAP7_75t_L g895 ( 
.A(n_651),
.B(n_516),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_714),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_653),
.B(n_583),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_638),
.B(n_508),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_694),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_716),
.B(n_516),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_716),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_755),
.B(n_515),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_R g903 ( 
.A(n_635),
.B(n_508),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_727),
.B(n_512),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_673),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_756),
.B(n_512),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_675),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_723),
.Y(n_908)
);

AOI221xp5_ASAP7_75t_SL g909 ( 
.A1(n_677),
.A2(n_517),
.B1(n_513),
.B2(n_522),
.C(n_521),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_699),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_609),
.A2(n_513),
.B1(n_517),
.B2(n_585),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_723),
.B(n_583),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_758),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_758),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_678),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_640),
.A2(n_585),
.B1(n_583),
.B2(n_521),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_622),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_682),
.B(n_583),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_SL g919 ( 
.A1(n_732),
.A2(n_717),
.B1(n_718),
.B2(n_701),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_683),
.B(n_585),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_684),
.B(n_585),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_700),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_643),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_610),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_730),
.B(n_394),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_650),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_713),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_661),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_640),
.B(n_571),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_731),
.B(n_685),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_661),
.Y(n_931)
);

NOR2x1_ASAP7_75t_R g932 ( 
.A(n_687),
.B(n_209),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_669),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_692),
.B(n_585),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_655),
.A2(n_689),
.B1(n_687),
.B2(n_737),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_689),
.B(n_216),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_764),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_801),
.A2(n_852),
.B(n_782),
.Y(n_938)
);

OAI22x1_ASAP7_75t_L g939 ( 
.A1(n_763),
.A2(n_655),
.B1(n_695),
.B2(n_743),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_801),
.A2(n_736),
.B(n_669),
.C(n_746),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_899),
.B(n_742),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_782),
.A2(n_713),
.B(n_725),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_828),
.A2(n_725),
.B1(n_743),
.B2(n_726),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_910),
.B(n_786),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_780),
.B(n_695),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_789),
.A2(n_726),
.B(n_720),
.Y(n_946)
);

NOR3xp33_ASAP7_75t_SL g947 ( 
.A(n_802),
.B(n_815),
.C(n_783),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_762),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_769),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_771),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_771),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_786),
.B(n_708),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_793),
.A2(n_930),
.B(n_862),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_770),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_823),
.A2(n_720),
.B(n_709),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_772),
.B(n_709),
.C(n_708),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_823),
.A2(n_753),
.B(n_273),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_918),
.A2(n_265),
.B(n_222),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_918),
.A2(n_274),
.B(n_231),
.Y(n_959)
);

XOR2x2_ASAP7_75t_SL g960 ( 
.A(n_766),
.B(n_8),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_917),
.A2(n_284),
.B1(n_234),
.B2(n_237),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_856),
.B(n_867),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_851),
.B(n_285),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_894),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_SL g965 ( 
.A(n_776),
.B(n_221),
.C(n_241),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_807),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_795),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_859),
.A2(n_394),
.B(n_396),
.C(n_242),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_920),
.A2(n_296),
.B(n_250),
.Y(n_969)
);

HB1xp67_ASAP7_75t_L g970 ( 
.A(n_795),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_850),
.B(n_293),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_855),
.B(n_243),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_809),
.B(n_394),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_774),
.B(n_305),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_791),
.A2(n_303),
.B1(n_264),
.B2(n_301),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_775),
.B(n_396),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_844),
.A2(n_396),
.B(n_422),
.C(n_443),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_R g978 ( 
.A(n_777),
.B(n_255),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_771),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_808),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_883),
.A2(n_396),
.B(n_571),
.C(n_422),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_867),
.B(n_10),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_935),
.A2(n_396),
.B(n_443),
.C(n_422),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_907),
.A2(n_12),
.B(n_13),
.C(n_18),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_904),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_819),
.B(n_396),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_873),
.B(n_881),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_SL g988 ( 
.A1(n_934),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_936),
.A2(n_396),
.B(n_443),
.C(n_422),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_831),
.B(n_20),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_843),
.A2(n_919),
.B1(n_761),
.B2(n_787),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_915),
.A2(n_21),
.B(n_25),
.C(n_26),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_920),
.A2(n_68),
.B(n_155),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_796),
.A2(n_443),
.B(n_422),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_785),
.B(n_67),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_785),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_834),
.B(n_25),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_760),
.A2(n_443),
.B(n_422),
.C(n_28),
.Y(n_998)
);

INVx8_ASAP7_75t_L g999 ( 
.A(n_818),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_816),
.A2(n_443),
.B1(n_422),
.B2(n_28),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_917),
.B(n_26),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_760),
.A2(n_443),
.B1(n_30),
.B2(n_32),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_816),
.A2(n_443),
.B1(n_33),
.B2(n_35),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_905),
.B(n_27),
.Y(n_1004)
);

AOI22x1_ASAP7_75t_L g1005 ( 
.A1(n_923),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_866),
.B(n_46),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_849),
.B(n_52),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_781),
.A2(n_52),
.B(n_56),
.C(n_59),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_917),
.B(n_78),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_778),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_921),
.A2(n_80),
.B(n_92),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_812),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_921),
.A2(n_99),
.B(n_104),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_860),
.B(n_109),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_854),
.B(n_122),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_917),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_773),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_779),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_926),
.B(n_924),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_835),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_860),
.B(n_144),
.Y(n_1021)
);

NAND2x1_ASAP7_75t_L g1022 ( 
.A(n_812),
.B(n_150),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_790),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_781),
.A2(n_898),
.B(n_874),
.C(n_841),
.Y(n_1024)
);

AOI221xp5_ASAP7_75t_L g1025 ( 
.A1(n_826),
.A2(n_829),
.B1(n_814),
.B2(n_817),
.C(n_806),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_872),
.B(n_876),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_788),
.B(n_792),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_869),
.A2(n_844),
.B(n_820),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_922),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_868),
.B(n_784),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_832),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_835),
.A2(n_818),
.B1(n_765),
.B2(n_845),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_904),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_838),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_839),
.B(n_842),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_858),
.B(n_847),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_847),
.B(n_875),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_830),
.A2(n_933),
.B(n_928),
.C(n_931),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_860),
.B(n_848),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_848),
.B(n_800),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_818),
.B(n_800),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_871),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_864),
.A2(n_865),
.B(n_768),
.C(n_869),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_890),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_SL g1045 ( 
.A(n_796),
.B(n_821),
.C(n_887),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_871),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_798),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_R g1048 ( 
.A(n_778),
.B(n_824),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_SL g1049 ( 
.A1(n_803),
.A2(n_805),
.B(n_813),
.C(n_822),
.Y(n_1049)
);

AO22x1_ASAP7_75t_L g1050 ( 
.A1(n_811),
.A2(n_878),
.B1(n_908),
.B2(n_861),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_822),
.A2(n_875),
.B(n_911),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_863),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_824),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_798),
.A2(n_911),
.B1(n_904),
.B2(n_906),
.Y(n_1054)
);

NAND2x1p5_ASAP7_75t_L g1055 ( 
.A(n_878),
.B(n_908),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_895),
.B(n_811),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_912),
.A2(n_825),
.B(n_799),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_794),
.B(n_906),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_833),
.B(n_794),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_833),
.B(n_794),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_846),
.A2(n_805),
.B1(n_803),
.B2(n_892),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_794),
.B(n_884),
.Y(n_1062)
);

BUFx8_ASAP7_75t_SL g1063 ( 
.A(n_922),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_886),
.B(n_893),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_794),
.B(n_922),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_870),
.A2(n_927),
.B1(n_878),
.B2(n_908),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_896),
.B(n_914),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_901),
.A2(n_913),
.B1(n_929),
.B2(n_861),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_932),
.B(n_927),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_870),
.A2(n_927),
.B1(n_908),
.B2(n_878),
.Y(n_1070)
);

AOI211x1_ASAP7_75t_L g1071 ( 
.A1(n_990),
.A2(n_810),
.B(n_836),
.C(n_891),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_1057),
.A2(n_877),
.B(n_880),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_948),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_SL g1074 ( 
.A1(n_991),
.A2(n_836),
.B(n_912),
.Y(n_1074)
);

NAND2x1p5_ASAP7_75t_L g1075 ( 
.A(n_1012),
.B(n_827),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_971),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_938),
.B(n_884),
.Y(n_1077)
);

NOR2x1_ASAP7_75t_SL g1078 ( 
.A(n_1012),
.B(n_895),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1028),
.A2(n_925),
.B(n_900),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1037),
.B(n_877),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_963),
.B(n_837),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1012),
.Y(n_1082)
);

INVx5_ASAP7_75t_L g1083 ( 
.A(n_999),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_972),
.B(n_837),
.Y(n_1084)
);

AOI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_964),
.A2(n_853),
.B1(n_909),
.B2(n_885),
.C(n_897),
.Y(n_1085)
);

AOI221x1_ASAP7_75t_L g1086 ( 
.A1(n_939),
.A2(n_888),
.B1(n_900),
.B2(n_882),
.C(n_880),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_994),
.A2(n_888),
.B(n_882),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1024),
.A2(n_916),
.B(n_840),
.C(n_797),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_953),
.A2(n_879),
.B(n_889),
.Y(n_1089)
);

OAI22x1_ASAP7_75t_L g1090 ( 
.A1(n_1032),
.A2(n_929),
.B1(n_804),
.B2(n_767),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1051),
.A2(n_879),
.B(n_895),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1002),
.A2(n_857),
.B1(n_804),
.B2(n_767),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_942),
.A2(n_909),
.B(n_903),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_940),
.A2(n_902),
.B(n_1043),
.C(n_945),
.Y(n_1094)
);

NAND2x1_ASAP7_75t_L g1095 ( 
.A(n_1047),
.B(n_1053),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_962),
.B(n_987),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_964),
.A2(n_992),
.B(n_984),
.C(n_941),
.Y(n_1097)
);

NAND2xp33_ASAP7_75t_L g1098 ( 
.A(n_1012),
.B(n_1047),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_940),
.A2(n_992),
.B(n_984),
.C(n_956),
.Y(n_1099)
);

AO32x2_ASAP7_75t_L g1100 ( 
.A1(n_1054),
.A2(n_943),
.A3(n_1061),
.B1(n_1070),
.B2(n_1066),
.Y(n_1100)
);

BUFx4_ASAP7_75t_SL g1101 ( 
.A(n_1010),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1045),
.A2(n_955),
.B(n_977),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1069),
.A2(n_974),
.B1(n_967),
.B2(n_975),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1026),
.B(n_1019),
.Y(n_1104)
);

AO21x2_ASAP7_75t_L g1105 ( 
.A1(n_946),
.A2(n_1060),
.B(n_1059),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_977),
.A2(n_1062),
.B(n_1065),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_966),
.B(n_1027),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_980),
.B(n_1023),
.Y(n_1108)
);

CKINVDCx11_ASAP7_75t_R g1109 ( 
.A(n_1020),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_966),
.B(n_1025),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1049),
.A2(n_1058),
.B(n_1015),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1056),
.Y(n_1112)
);

AO22x2_ASAP7_75t_L g1113 ( 
.A1(n_960),
.A2(n_1030),
.B1(n_1001),
.B2(n_1044),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_949),
.B(n_1017),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1018),
.B(n_1064),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_980),
.B(n_970),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1067),
.B(n_1035),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_956),
.A2(n_1007),
.B(n_982),
.C(n_1003),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1056),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1036),
.B(n_1031),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_SL g1121 ( 
.A(n_1052),
.B(n_978),
.C(n_997),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_968),
.A2(n_1009),
.B(n_1050),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_970),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_SL g1124 ( 
.A1(n_988),
.A2(n_1022),
.B(n_1008),
.C(n_998),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_967),
.B(n_1041),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1063),
.Y(n_1126)
);

NOR2x1_ASAP7_75t_SL g1127 ( 
.A(n_1029),
.B(n_1053),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1038),
.A2(n_957),
.A3(n_983),
.B(n_981),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_993),
.A2(n_1013),
.B(n_1011),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1055),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1048),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1034),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1055),
.A2(n_976),
.B(n_1016),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1068),
.A2(n_952),
.B(n_985),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_958),
.A2(n_969),
.B(n_959),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_1046),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1002),
.A2(n_1045),
.B1(n_1004),
.B2(n_1005),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_989),
.A2(n_985),
.B(n_1033),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_937),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1033),
.A2(n_1014),
.B(n_1021),
.Y(n_1140)
);

AO21x2_ASAP7_75t_L g1141 ( 
.A1(n_1006),
.A2(n_961),
.B(n_973),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_950),
.B(n_951),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_986),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1040),
.A2(n_1029),
.B(n_999),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_SL g1145 ( 
.A1(n_1000),
.A2(n_1039),
.B(n_947),
.C(n_965),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_999),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_950),
.A2(n_951),
.B(n_979),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_950),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_996),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_947),
.A2(n_950),
.B(n_951),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1042),
.B(n_965),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_951),
.A2(n_979),
.B(n_995),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_979),
.B(n_774),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_979),
.A2(n_1057),
.B(n_994),
.Y(n_1154)
);

NAND3x1_ASAP7_75t_L g1155 ( 
.A(n_1032),
.B(n_763),
.C(n_1069),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_954),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_938),
.B(n_991),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_939),
.A2(n_1024),
.A3(n_760),
.B(n_781),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_937),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_938),
.A2(n_852),
.B(n_1028),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_L g1161 ( 
.A(n_991),
.B(n_397),
.C(n_763),
.Y(n_1161)
);

AO32x2_ASAP7_75t_L g1162 ( 
.A1(n_1054),
.A2(n_943),
.A3(n_796),
.B1(n_420),
.B2(n_1061),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_948),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_991),
.A2(n_801),
.B1(n_763),
.B2(n_852),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_991),
.A2(n_763),
.B(n_636),
.C(n_859),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_937),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_938),
.A2(n_852),
.B(n_1028),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1057),
.A2(n_994),
.B(n_942),
.Y(n_1168)
);

AND2x2_ASAP7_75t_SL g1169 ( 
.A(n_1002),
.B(n_582),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1057),
.A2(n_994),
.B(n_942),
.Y(n_1170)
);

CKINVDCx11_ASAP7_75t_R g1171 ( 
.A(n_1020),
.Y(n_1171)
);

BUFx10_ASAP7_75t_L g1172 ( 
.A(n_996),
.Y(n_1172)
);

AO21x1_ASAP7_75t_L g1173 ( 
.A1(n_938),
.A2(n_852),
.B(n_974),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_938),
.B(n_991),
.Y(n_1174)
);

AO32x2_ASAP7_75t_L g1175 ( 
.A1(n_1054),
.A2(n_943),
.A3(n_796),
.B1(n_420),
.B2(n_1061),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1024),
.A2(n_801),
.B(n_505),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_938),
.B(n_991),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_954),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1057),
.A2(n_994),
.B(n_942),
.Y(n_1179)
);

INVx6_ASAP7_75t_L g1180 ( 
.A(n_1020),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_991),
.A2(n_763),
.B(n_636),
.C(n_859),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_991),
.A2(n_851),
.B1(n_780),
.B2(n_528),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1028),
.A2(n_938),
.B(n_1051),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_938),
.A2(n_852),
.B(n_1028),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_938),
.B(n_991),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_948),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1057),
.A2(n_994),
.B(n_942),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_938),
.B(n_991),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_939),
.A2(n_1024),
.A3(n_760),
.B(n_781),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_991),
.A2(n_801),
.B1(n_763),
.B2(n_852),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_938),
.B(n_991),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_938),
.A2(n_852),
.B(n_1028),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_R g1193 ( 
.A(n_1010),
.B(n_478),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_944),
.B(n_780),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_944),
.B(n_780),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1057),
.A2(n_994),
.B(n_942),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1057),
.A2(n_994),
.B(n_942),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1056),
.B(n_786),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_938),
.A2(n_852),
.B(n_1028),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_938),
.B(n_991),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1086),
.A2(n_1183),
.B(n_1199),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1169),
.A2(n_1161),
.B1(n_1113),
.B2(n_1164),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1183),
.A2(n_1199),
.B(n_1170),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1083),
.B(n_1112),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1165),
.A2(n_1181),
.B(n_1190),
.C(n_1164),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1139),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1190),
.A2(n_1094),
.B(n_1137),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1137),
.A2(n_1182),
.B(n_1099),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1114),
.Y(n_1209)
);

INVx8_ASAP7_75t_L g1210 ( 
.A(n_1198),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_L g1211 ( 
.A1(n_1097),
.A2(n_1113),
.B1(n_1118),
.B2(n_1200),
.C(n_1191),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1160),
.A2(n_1184),
.B(n_1167),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1180),
.Y(n_1213)
);

AOI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1157),
.A2(n_1200),
.B1(n_1174),
.B2(n_1177),
.C(n_1191),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1114),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1104),
.B(n_1117),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1073),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1105),
.Y(n_1218)
);

NOR3xp33_ASAP7_75t_L g1219 ( 
.A(n_1157),
.B(n_1174),
.C(n_1177),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1168),
.A2(n_1187),
.B(n_1179),
.Y(n_1220)
);

BUFx8_ASAP7_75t_L g1221 ( 
.A(n_1076),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1105),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1132),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1193),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1163),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1185),
.A2(n_1188),
.B(n_1192),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_SL g1227 ( 
.A1(n_1185),
.A2(n_1188),
.B1(n_1110),
.B2(n_1151),
.C(n_1107),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1154),
.A2(n_1129),
.B(n_1079),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1180),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1102),
.A2(n_1091),
.B(n_1072),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1110),
.A2(n_1103),
.B1(n_1155),
.B2(n_1107),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1158),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1186),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1176),
.A2(n_1088),
.B(n_1085),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1123),
.Y(n_1235)
);

AOI221x1_ASAP7_75t_L g1236 ( 
.A1(n_1140),
.A2(n_1138),
.B1(n_1111),
.B2(n_1102),
.C(n_1122),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1129),
.A2(n_1089),
.B(n_1087),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1106),
.A2(n_1111),
.B(n_1093),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1077),
.A2(n_1133),
.B(n_1138),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1158),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1085),
.A2(n_1077),
.B(n_1084),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1121),
.A2(n_1096),
.B1(n_1081),
.B2(n_1108),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1083),
.B(n_1152),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1135),
.A2(n_1074),
.B(n_1092),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1115),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1131),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1173),
.A2(n_1134),
.B(n_1153),
.Y(n_1247)
);

INVx4_ASAP7_75t_L g1248 ( 
.A(n_1166),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1083),
.B(n_1119),
.Y(n_1249)
);

INVx5_ASAP7_75t_SL g1250 ( 
.A(n_1198),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1150),
.A2(n_1080),
.B(n_1147),
.Y(n_1251)
);

AO21x2_ASAP7_75t_L g1252 ( 
.A1(n_1141),
.A2(n_1124),
.B(n_1120),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1159),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1104),
.B(n_1117),
.Y(n_1254)
);

NAND2x1p5_ASAP7_75t_L g1255 ( 
.A(n_1083),
.B(n_1152),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1120),
.A2(n_1130),
.B(n_1075),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1090),
.A2(n_1143),
.B(n_1095),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1098),
.A2(n_1141),
.B(n_1127),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1082),
.A2(n_1144),
.B(n_1148),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1145),
.A2(n_1071),
.B1(n_1178),
.B2(n_1156),
.C(n_1162),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1166),
.B(n_1125),
.C(n_1126),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1142),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1112),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1162),
.A2(n_1175),
.B(n_1189),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1078),
.A2(n_1175),
.B(n_1162),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1175),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1128),
.A2(n_1119),
.B(n_1189),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1158),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1189),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1149),
.A2(n_1146),
.B(n_1100),
.C(n_1101),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1172),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1128),
.B(n_1136),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1172),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1100),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1100),
.B(n_1109),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1128),
.A2(n_1181),
.B(n_1165),
.C(n_1161),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1171),
.A2(n_1170),
.B(n_1168),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1166),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1114),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1116),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1161),
.A2(n_1182),
.B1(n_1169),
.B2(n_851),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1114),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1104),
.B(n_1194),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1161),
.A2(n_1181),
.B(n_1165),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1086),
.A2(n_1183),
.B(n_1199),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_1157),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1114),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1161),
.A2(n_1182),
.B1(n_1169),
.B2(n_851),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1168),
.A2(n_1197),
.B(n_1196),
.Y(n_1289)
);

CKINVDCx8_ASAP7_75t_R g1290 ( 
.A(n_1136),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1114),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_1157),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1105),
.Y(n_1293)
);

AND2x6_ASAP7_75t_L g1294 ( 
.A(n_1157),
.B(n_1174),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1114),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1193),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1161),
.A2(n_1181),
.B(n_1165),
.Y(n_1297)
);

XOR2xp5_ASAP7_75t_L g1298 ( 
.A(n_1136),
.B(n_540),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1161),
.B(n_1181),
.C(n_1165),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1165),
.A2(n_1181),
.B(n_1190),
.C(n_1164),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_1139),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1168),
.A2(n_1197),
.B(n_1196),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1194),
.B(n_1195),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1180),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1168),
.A2(n_1197),
.B(n_1196),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1168),
.A2(n_1197),
.B(n_1196),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1114),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1139),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1105),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1083),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1116),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1161),
.A2(n_1182),
.B1(n_1181),
.B2(n_1165),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1114),
.Y(n_1313)
);

BUFx4f_ASAP7_75t_SL g1314 ( 
.A(n_1172),
.Y(n_1314)
);

OAI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1161),
.A2(n_1182),
.B1(n_1190),
.B2(n_1164),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1161),
.A2(n_1182),
.B1(n_1190),
.B2(n_1164),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1168),
.A2(n_1197),
.B(n_1196),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1104),
.B(n_1194),
.Y(n_1318)
);

INVx3_ASAP7_75t_SL g1319 ( 
.A(n_1136),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1083),
.B(n_1112),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1168),
.A2(n_1197),
.B(n_1196),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1086),
.A2(n_939),
.A3(n_1024),
.B(n_1173),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1168),
.A2(n_1197),
.B(n_1196),
.Y(n_1323)
);

INVx3_ASAP7_75t_SL g1324 ( 
.A(n_1136),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1205),
.A2(n_1300),
.B(n_1207),
.C(n_1208),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1283),
.B(n_1318),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1217),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1290),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1315),
.A2(n_1316),
.B1(n_1288),
.B2(n_1281),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1216),
.B(n_1254),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1253),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1303),
.B(n_1245),
.Y(n_1332)
);

O2A1O1Ixp5_ASAP7_75t_L g1333 ( 
.A1(n_1315),
.A2(n_1316),
.B(n_1284),
.C(n_1297),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1209),
.B(n_1215),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1299),
.A2(n_1202),
.B1(n_1312),
.B2(n_1211),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1202),
.A2(n_1276),
.B1(n_1231),
.B2(n_1234),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_SL g1337 ( 
.A1(n_1226),
.A2(n_1212),
.B(n_1273),
.C(n_1219),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1279),
.B(n_1282),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_SL g1339 ( 
.A1(n_1270),
.A2(n_1275),
.B(n_1241),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1219),
.A2(n_1275),
.B(n_1272),
.C(n_1214),
.Y(n_1340)
);

O2A1O1Ixp5_ASAP7_75t_L g1341 ( 
.A1(n_1286),
.A2(n_1292),
.B(n_1258),
.C(n_1257),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1265),
.A2(n_1227),
.B(n_1260),
.C(n_1244),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1240),
.A2(n_1222),
.B(n_1218),
.C(n_1274),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1206),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1301),
.A2(n_1308),
.B1(n_1242),
.B2(n_1235),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1236),
.A2(n_1237),
.B(n_1228),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_L g1347 ( 
.A(n_1261),
.B(n_1248),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1246),
.A2(n_1224),
.B1(n_1296),
.B2(n_1248),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1287),
.B(n_1291),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1295),
.B(n_1307),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1223),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1224),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1262),
.B(n_1263),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1204),
.A2(n_1249),
.B(n_1320),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1237),
.A2(n_1228),
.B(n_1238),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1313),
.B(n_1294),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1225),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1266),
.A2(n_1247),
.B(n_1239),
.C(n_1269),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1296),
.A2(n_1278),
.B1(n_1229),
.B2(n_1304),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1213),
.A2(n_1271),
.B(n_1273),
.C(n_1233),
.Y(n_1360)
);

AOI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1293),
.A2(n_1309),
.B(n_1268),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_SL g1362 ( 
.A(n_1221),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1232),
.A2(n_1269),
.B(n_1268),
.C(n_1309),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1247),
.A2(n_1239),
.B(n_1232),
.C(n_1267),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1250),
.B(n_1256),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1238),
.A2(n_1305),
.B(n_1289),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1294),
.B(n_1264),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1250),
.B(n_1256),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1278),
.A2(n_1314),
.B1(n_1298),
.B2(n_1264),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1264),
.B(n_1252),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1319),
.A2(n_1324),
.B(n_1252),
.C(n_1201),
.Y(n_1371)
);

AND2x2_ASAP7_75t_SL g1372 ( 
.A(n_1201),
.B(n_1285),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1230),
.A2(n_1201),
.B(n_1285),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1319),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1221),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1310),
.A2(n_1255),
.B(n_1243),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1221),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1267),
.A2(n_1240),
.B(n_1210),
.C(n_1294),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1277),
.A2(n_1314),
.B(n_1203),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1324),
.A2(n_1210),
.B1(n_1310),
.B2(n_1203),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1310),
.A2(n_1243),
.B(n_1255),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1222),
.A2(n_1322),
.B(n_1251),
.C(n_1259),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1322),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1322),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1220),
.B(n_1323),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1302),
.B(n_1305),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1302),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1306),
.A2(n_1317),
.B(n_1321),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1317),
.B(n_1321),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1323),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1280),
.B(n_1311),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1315),
.A2(n_1161),
.B1(n_1182),
.B2(n_1316),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1283),
.B(n_1318),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1280),
.B(n_1311),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_1261),
.B(n_1248),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1280),
.B(n_1311),
.Y(n_1396)
);

NOR2xp67_ASAP7_75t_R g1397 ( 
.A(n_1248),
.B(n_1180),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1315),
.A2(n_1161),
.B(n_1316),
.C(n_1181),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1283),
.B(n_1318),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1236),
.A2(n_1212),
.B(n_1237),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1205),
.A2(n_1181),
.B(n_1165),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1207),
.A2(n_1300),
.B(n_1205),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1205),
.A2(n_1181),
.B(n_1165),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_1207),
.A2(n_1316),
.B(n_1315),
.C(n_1297),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1280),
.B(n_1311),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1293),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1217),
.Y(n_1407)
);

CKINVDCx16_ASAP7_75t_R g1408 ( 
.A(n_1298),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1327),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1372),
.B(n_1367),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1406),
.B(n_1383),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1351),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1406),
.B(n_1383),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1384),
.B(n_1356),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1385),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1373),
.A2(n_1364),
.B(n_1358),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1384),
.B(n_1346),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1357),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1407),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1370),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_SL g1422 ( 
.A(n_1362),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1334),
.B(n_1338),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1400),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1346),
.B(n_1400),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1344),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1349),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1387),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1350),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1386),
.B(n_1394),
.Y(n_1430)
);

AO21x2_ASAP7_75t_L g1431 ( 
.A1(n_1364),
.A2(n_1358),
.B(n_1342),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1343),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1342),
.A2(n_1382),
.B(n_1336),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1404),
.A2(n_1333),
.B(n_1398),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1343),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1405),
.B(n_1390),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1388),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1376),
.B(n_1381),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1363),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1401),
.A2(n_1403),
.B(n_1404),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1402),
.B(n_1325),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1389),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1332),
.B(n_1378),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1325),
.A2(n_1335),
.B(n_1392),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1388),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1341),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1329),
.A2(n_1345),
.B1(n_1408),
.B2(n_1326),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1378),
.B(n_1369),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1379),
.A2(n_1361),
.B(n_1355),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1333),
.A2(n_1362),
.B1(n_1339),
.B2(n_1340),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1330),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1354),
.B(n_1371),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1366),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1366),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1437),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1442),
.B(n_1337),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1415),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1410),
.B(n_1355),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1441),
.B(n_1440),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1442),
.Y(n_1460)
);

NAND4xp25_ASAP7_75t_L g1461 ( 
.A(n_1444),
.B(n_1337),
.C(n_1348),
.D(n_1360),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1452),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1437),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1441),
.A2(n_1434),
.B1(n_1447),
.B2(n_1440),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1449),
.A2(n_1379),
.B(n_1361),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1411),
.B(n_1355),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1428),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1428),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1410),
.B(n_1353),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1434),
.B(n_1331),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1409),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1415),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1414),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_1445),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1422),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1411),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1446),
.B(n_1399),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1411),
.B(n_1393),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1413),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1413),
.B(n_1380),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1415),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1467),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1464),
.A2(n_1433),
.B1(n_1448),
.B2(n_1431),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1465),
.A2(n_1449),
.B(n_1435),
.Y(n_1484)
);

OAI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1464),
.A2(n_1447),
.B1(n_1450),
.B2(n_1448),
.C(n_1439),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1469),
.B(n_1430),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1459),
.A2(n_1448),
.B1(n_1450),
.B2(n_1452),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1460),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1477),
.B(n_1427),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1462),
.A2(n_1433),
.B1(n_1431),
.B2(n_1452),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1463),
.Y(n_1491)
);

OAI33xp33_ASAP7_75t_L g1492 ( 
.A1(n_1459),
.A2(n_1439),
.A3(n_1423),
.B1(n_1418),
.B2(n_1427),
.B3(n_1429),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1467),
.Y(n_1493)
);

NAND4xp25_ASAP7_75t_L g1494 ( 
.A(n_1461),
.B(n_1456),
.C(n_1470),
.D(n_1425),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1470),
.A2(n_1433),
.B1(n_1431),
.B2(n_1451),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1460),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1469),
.B(n_1430),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1467),
.Y(n_1498)
);

AOI31xp33_ASAP7_75t_L g1499 ( 
.A1(n_1475),
.A2(n_1446),
.A3(n_1443),
.B(n_1359),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1476),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1456),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1456),
.B(n_1424),
.C(n_1417),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1468),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1461),
.A2(n_1433),
.B1(n_1431),
.B2(n_1451),
.Y(n_1504)
);

AOI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1477),
.A2(n_1417),
.B1(n_1432),
.B2(n_1443),
.C(n_1424),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1480),
.A2(n_1452),
.B1(n_1443),
.B2(n_1418),
.Y(n_1506)
);

OAI221xp5_ASAP7_75t_L g1507 ( 
.A1(n_1461),
.A2(n_1452),
.B1(n_1432),
.B2(n_1414),
.C(n_1421),
.Y(n_1507)
);

AOI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1455),
.A2(n_1454),
.B(n_1453),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1478),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_1477),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1476),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1473),
.B(n_1429),
.Y(n_1512)
);

AOI33xp33_ASAP7_75t_L g1513 ( 
.A1(n_1458),
.A2(n_1417),
.A3(n_1412),
.B1(n_1419),
.B2(n_1420),
.B3(n_1436),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1462),
.B(n_1438),
.Y(n_1514)
);

AO21x2_ASAP7_75t_L g1515 ( 
.A1(n_1474),
.A2(n_1435),
.B(n_1416),
.Y(n_1515)
);

NOR4xp25_ASAP7_75t_SL g1516 ( 
.A(n_1475),
.B(n_1481),
.C(n_1457),
.D(n_1472),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1479),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1499),
.B(n_1457),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1502),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1508),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1508),
.Y(n_1521)
);

INVx5_ASAP7_75t_L g1522 ( 
.A(n_1514),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1515),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1482),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1486),
.B(n_1458),
.Y(n_1525)
);

INVx4_ASAP7_75t_SL g1526 ( 
.A(n_1514),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1491),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1493),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1515),
.A2(n_1435),
.B(n_1416),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1501),
.B(n_1473),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1510),
.B(n_1479),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1509),
.B(n_1458),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1486),
.B(n_1497),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1497),
.B(n_1458),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1496),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1498),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1498),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

NOR2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1494),
.B(n_1377),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1500),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1515),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1488),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1484),
.Y(n_1545)
);

OAI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1494),
.A2(n_1480),
.B(n_1466),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1515),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1509),
.B(n_1471),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1511),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1519),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1530),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1534),
.B(n_1516),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1524),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_1516),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1530),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1542),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1524),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1519),
.A2(n_1485),
.B1(n_1483),
.B2(n_1504),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1546),
.B(n_1505),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1489),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1518),
.B(n_1488),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1546),
.B(n_1505),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1527),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1517),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1525),
.B(n_1535),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1527),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1531),
.B(n_1489),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1536),
.B(n_1499),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1529),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1542),
.A2(n_1487),
.B(n_1502),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1529),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1536),
.B(n_1512),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1549),
.B(n_1512),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1532),
.B(n_1478),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1525),
.B(n_1469),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1507),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1544),
.B(n_1526),
.Y(n_1579)
);

NAND4xp25_ASAP7_75t_L g1580 ( 
.A(n_1544),
.B(n_1485),
.C(n_1507),
.D(n_1487),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1530),
.Y(n_1581)
);

CKINVDCx16_ASAP7_75t_R g1582 ( 
.A(n_1544),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1537),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1525),
.B(n_1469),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1532),
.B(n_1478),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1549),
.B(n_1478),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1544),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1541),
.B(n_1506),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1579),
.B(n_1514),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1579),
.Y(n_1590)
);

O2A1O1Ixp33_ASAP7_75t_SL g1591 ( 
.A1(n_1561),
.A2(n_1375),
.B(n_1533),
.C(n_1528),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1576),
.B(n_1533),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1576),
.B(n_1548),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1535),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1553),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1560),
.B(n_1506),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1550),
.B(n_1558),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1550),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1564),
.B(n_1537),
.Y(n_1601)
);

NOR2x1p5_ASAP7_75t_SL g1602 ( 
.A(n_1559),
.B(n_1520),
.Y(n_1602)
);

NAND2x1_ASAP7_75t_L g1603 ( 
.A(n_1579),
.B(n_1528),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1579),
.B(n_1522),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1538),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1582),
.B(n_1538),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1559),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1585),
.B(n_1418),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1567),
.B(n_1577),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1565),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1587),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1587),
.B(n_1555),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1555),
.B(n_1539),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1565),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1569),
.B(n_1539),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1568),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1495),
.C(n_1490),
.D(n_1426),
.Y(n_1617)
);

AND4x1_ASAP7_75t_L g1618 ( 
.A(n_1578),
.B(n_1492),
.C(n_1422),
.D(n_1397),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1567),
.B(n_1526),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1426),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.B(n_1540),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1580),
.A2(n_1530),
.B1(n_1520),
.B2(n_1521),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1540),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1622),
.B(n_1562),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1604),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1618),
.B(n_1578),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1609),
.B(n_1572),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

NAND2x1_ASAP7_75t_SL g1630 ( 
.A(n_1611),
.B(n_1563),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1622),
.B(n_1580),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1601),
.B(n_1574),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1598),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1612),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1590),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1619),
.B(n_1563),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1594),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1619),
.B(n_1584),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1621),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1597),
.A2(n_1551),
.B(n_1556),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1623),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1604),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1596),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1607),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1610),
.B(n_1575),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1614),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1620),
.B(n_1584),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_1568),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1629),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1627),
.A2(n_1595),
.B(n_1617),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1636),
.B(n_1566),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1629),
.Y(n_1652)
);

AOI322xp5_ASAP7_75t_L g1653 ( 
.A1(n_1631),
.A2(n_1613),
.A3(n_1617),
.B1(n_1520),
.B2(n_1521),
.C1(n_1554),
.C2(n_1552),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1629),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1631),
.A2(n_1589),
.B1(n_1588),
.B2(n_1552),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1637),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1636),
.B(n_1566),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1635),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1637),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1624),
.A2(n_1589),
.B1(n_1554),
.B2(n_1521),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1639),
.B(n_1602),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1624),
.A2(n_1589),
.B1(n_1557),
.B2(n_1581),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1615),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1643),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1643),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1632),
.A2(n_1522),
.B1(n_1608),
.B2(n_1592),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1632),
.A2(n_1520),
.B1(n_1521),
.B2(n_1591),
.C(n_1606),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1649),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1658),
.B(n_1634),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1651),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1652),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1657),
.B(n_1634),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1654),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1663),
.B(n_1639),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1661),
.B(n_1635),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1663),
.B(n_1641),
.Y(n_1676)
);

NOR2x1_ASAP7_75t_L g1677 ( 
.A(n_1661),
.B(n_1626),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1678)
);

AOI221xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1660),
.B1(n_1662),
.B2(n_1655),
.C(n_1667),
.Y(n_1679)
);

AOI211xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1669),
.A2(n_1633),
.B(n_1666),
.C(n_1626),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1677),
.A2(n_1653),
.B1(n_1630),
.B2(n_1676),
.C(n_1674),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1671),
.A2(n_1630),
.B(n_1628),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1675),
.Y(n_1684)
);

OAI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1671),
.A2(n_1633),
.B(n_1664),
.C(n_1659),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1668),
.A2(n_1665),
.B(n_1656),
.C(n_1628),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1672),
.B(n_1673),
.Y(n_1687)
);

OAI21xp33_ASAP7_75t_L g1688 ( 
.A1(n_1678),
.A2(n_1638),
.B(n_1645),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1677),
.A2(n_1648),
.B(n_1642),
.Y(n_1689)
);

OAI21xp33_ASAP7_75t_L g1690 ( 
.A1(n_1683),
.A2(n_1645),
.B(n_1638),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1682),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1689),
.A2(n_1648),
.B(n_1625),
.Y(n_1692)
);

OAI21xp33_ASAP7_75t_L g1693 ( 
.A1(n_1688),
.A2(n_1625),
.B(n_1642),
.Y(n_1693)
);

AOI22x1_ASAP7_75t_L g1694 ( 
.A1(n_1684),
.A2(n_1646),
.B1(n_1644),
.B2(n_1642),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1691),
.B(n_1687),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1690),
.B(n_1681),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1692),
.B(n_1680),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1694),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1693),
.B(n_1679),
.C(n_1685),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1691),
.B(n_1625),
.Y(n_1700)
);

INVx5_ASAP7_75t_L g1701 ( 
.A(n_1700),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_L g1702 ( 
.A(n_1699),
.B(n_1686),
.C(n_1646),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1697),
.Y(n_1703)
);

OAI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1696),
.A2(n_1644),
.B(n_1603),
.C(n_1605),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1695),
.A2(n_1698),
.B(n_1640),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1703),
.Y(n_1706)
);

NAND3x1_ASAP7_75t_L g1707 ( 
.A(n_1705),
.B(n_1701),
.C(n_1702),
.Y(n_1707)
);

AOI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1704),
.A2(n_1640),
.B1(n_1647),
.B2(n_1599),
.Y(n_1708)
);

NOR4xp75_ASAP7_75t_SL g1709 ( 
.A(n_1707),
.B(n_1374),
.C(n_1328),
.D(n_1352),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1709),
.A2(n_1706),
.B1(n_1708),
.B2(n_1593),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1710),
.B(n_1640),
.Y(n_1711)
);

OAI321xp33_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1556),
.A3(n_1557),
.B1(n_1551),
.B2(n_1581),
.C(n_1640),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1647),
.B1(n_1571),
.B2(n_1583),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1713),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1713),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1715),
.A2(n_1714),
.B1(n_1583),
.B2(n_1571),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1714),
.B(n_1523),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1717),
.A2(n_1543),
.B(n_1523),
.Y(n_1718)
);

NOR2xp33_ASAP7_75t_L g1719 ( 
.A(n_1716),
.B(n_1573),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1719),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1718),
.A2(n_1545),
.B1(n_1523),
.B2(n_1547),
.Y(n_1721)
);

AOI31xp33_ASAP7_75t_L g1722 ( 
.A1(n_1720),
.A2(n_1523),
.A3(n_1543),
.B(n_1547),
.Y(n_1722)
);

AOI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1721),
.B(n_1347),
.C(n_1395),
.Y(n_1723)
);


endmodule