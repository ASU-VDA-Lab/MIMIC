module fake_ariane_1079_n_2605 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_363, n_720, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_711, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_718, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_712, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_2605);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_363;
input n_720;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_711;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_2605;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_1442;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_931;
wire n_1491;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2312;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_2599;
wire n_727;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_2508;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_862;
wire n_1700;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_876;
wire n_791;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_1118;
wire n_943;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_2158;
wire n_2578;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_911;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_907;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_918;
wire n_1968;
wire n_1885;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_1781;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx2_ASAP7_75t_L g721 ( 
.A(n_129),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_119),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_616),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_375),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_600),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_495),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_631),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_633),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_606),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_674),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_422),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_465),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_196),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_461),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_650),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_651),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_190),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_713),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_162),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_182),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_653),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_187),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_449),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_111),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_593),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_706),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_676),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_46),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_531),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_398),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_618),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_198),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_459),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_672),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_664),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_408),
.Y(n_756)
);

BUFx10_ASAP7_75t_L g757 ( 
.A(n_426),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_442),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_678),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_393),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_645),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_592),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_605),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_708),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_197),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_215),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_416),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_639),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_527),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_153),
.Y(n_770)
);

BUFx10_ASAP7_75t_L g771 ( 
.A(n_451),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_689),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_714),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_528),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_590),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_686),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_654),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_636),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_173),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_701),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_499),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_166),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_458),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_684),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_611),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_709),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_372),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_634),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_640),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_628),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_637),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_42),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_707),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_586),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_644),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_283),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_136),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_312),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_619),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_643),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_705),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_572),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_550),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_33),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_660),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_670),
.Y(n_806)
);

CKINVDCx16_ASAP7_75t_R g807 ( 
.A(n_323),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_681),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_350),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_698),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_588),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_659),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_688),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_677),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_685),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_694),
.Y(n_816)
);

CKINVDCx14_ASAP7_75t_R g817 ( 
.A(n_683),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_695),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_635),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_601),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_594),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_90),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_191),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_646),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_317),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_582),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_668),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_219),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_236),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_487),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_427),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_621),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_129),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_655),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_680),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_679),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_454),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_388),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_692),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_703),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_284),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_394),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_613),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_642),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_265),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_319),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_669),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_506),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_622),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_675),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_124),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_23),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_663),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_700),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_718),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_411),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_157),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_406),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_720),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_38),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_526),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_693),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_130),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_610),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_137),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_321),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_143),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_596),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_30),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_59),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_35),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_597),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_110),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_240),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_711),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_303),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_589),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_22),
.Y(n_878)
);

BUFx10_ASAP7_75t_L g879 ( 
.A(n_666),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_627),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_712),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_629),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_334),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_61),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_607),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_608),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_276),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_37),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_432),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_715),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_61),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_60),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_435),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_323),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_702),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_623),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_599),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_265),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_28),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_345),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_437),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_206),
.Y(n_902)
);

CKINVDCx14_ASAP7_75t_R g903 ( 
.A(n_301),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_551),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_368),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_407),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_162),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_595),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_94),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_603),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_612),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_348),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_222),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_444),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_691),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_346),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_70),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_682),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_462),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_620),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_485),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_217),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_638),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_615),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_405),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_187),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_24),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_626),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_716),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_617),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_699),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_8),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_302),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_68),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_614),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_647),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_107),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_77),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_662),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_445),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_34),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_648),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_226),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_652),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_609),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_510),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_658),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_558),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_132),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_667),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_71),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_571),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_624),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_7),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_28),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_385),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_313),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_665),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_697),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_717),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_591),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_127),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_299),
.Y(n_963)
);

BUFx2_ASAP7_75t_SL g964 ( 
.A(n_630),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_354),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_95),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_224),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_247),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_333),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_3),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_413),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_656),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_704),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_149),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_401),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_587),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_259),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_476),
.Y(n_978)
);

BUFx10_ASAP7_75t_L g979 ( 
.A(n_305),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_111),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_436),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_673),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_118),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_470),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_210),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_48),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_439),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_625),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_274),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_671),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_35),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_657),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_132),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_632),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_330),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_309),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_254),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_409),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_710),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_378),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_602),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_580),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_260),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_690),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_641),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_223),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_649),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_687),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_502),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_310),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_696),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_477),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_604),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_598),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_493),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_62),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_51),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_661),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_118),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_37),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_752),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_807),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_903),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_731),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_779),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_745),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_760),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_878),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_793),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_803),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_792),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_796),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_804),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_825),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_805),
.Y(n_1035)
);

INVxp67_ASAP7_75t_SL g1036 ( 
.A(n_995),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_995),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_842),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_897),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_829),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_833),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_841),
.Y(n_1042)
);

INVxp67_ASAP7_75t_SL g1043 ( 
.A(n_995),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_852),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_894),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_863),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_870),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_905),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_871),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_874),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_888),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_892),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_947),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_L g1054 ( 
.A(n_1022),
.B(n_722),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1036),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_1024),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1037),
.Y(n_1057)
);

HB1xp67_ASAP7_75t_L g1058 ( 
.A(n_1053),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1043),
.B(n_758),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1028),
.A2(n_977),
.B1(n_969),
.B2(n_740),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1045),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1021),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1025),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1031),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1028),
.B(n_817),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1032),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_1033),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_1040),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1041),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_1042),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1044),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_1046),
.Y(n_1072)
);

AND2x6_ASAP7_75t_L g1073 ( 
.A(n_1047),
.B(n_747),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1023),
.A2(n_744),
.B1(n_899),
.B2(n_765),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1049),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_1030),
.Y(n_1076)
);

NOR2x1_ASAP7_75t_L g1077 ( 
.A(n_1050),
.B(n_854),
.Y(n_1077)
);

AND2x2_ASAP7_75t_R g1078 ( 
.A(n_1035),
.B(n_937),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1051),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1052),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1034),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1034),
.B(n_844),
.Y(n_1082)
);

INVxp33_ASAP7_75t_SL g1083 ( 
.A(n_1038),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_1039),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1048),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1062),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_1056),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1065),
.A2(n_876),
.B1(n_748),
.B2(n_851),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1061),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1081),
.B(n_767),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1055),
.B(n_965),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_1058),
.B(n_968),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_1076),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_1082),
.B(n_737),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1064),
.A2(n_917),
.B1(n_721),
.B2(n_958),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1057),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1059),
.B(n_761),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1071),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1079),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1080),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1067),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1067),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1068),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1068),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1069),
.B(n_739),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1063),
.B(n_1066),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1075),
.Y(n_1107)
);

INVxp67_ASAP7_75t_SL g1108 ( 
.A(n_1069),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1070),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1070),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1072),
.B(n_802),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1072),
.B(n_1026),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_1084),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1077),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_1073),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1073),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1073),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_1085),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1054),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1083),
.B(n_816),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1060),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1074),
.B(n_946),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_1078),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1064),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1061),
.Y(n_1125)
);

CKINVDCx6p67_ASAP7_75t_R g1126 ( 
.A(n_1058),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1064),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1065),
.B(n_742),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1064),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1081),
.B(n_1027),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1065),
.B(n_766),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1093),
.B(n_1029),
.Y(n_1132)
);

CKINVDCx6p67_ASAP7_75t_R g1133 ( 
.A(n_1113),
.Y(n_1133)
);

OR2x6_ASAP7_75t_L g1134 ( 
.A(n_1112),
.B(n_938),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1090),
.B(n_1008),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1097),
.B(n_886),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1118),
.B(n_982),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1089),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1086),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1119),
.A2(n_782),
.B1(n_797),
.B2(n_770),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1086),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1107),
.B(n_923),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1098),
.B(n_1002),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1118),
.B(n_1120),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1124),
.B(n_1127),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1118),
.B(n_1016),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_1130),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_1111),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1087),
.B(n_1019),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1099),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1125),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1129),
.B(n_798),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1096),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1100),
.B(n_1106),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1109),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1126),
.B(n_1020),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1122),
.A2(n_867),
.B1(n_955),
.B2(n_949),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1110),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1108),
.B(n_809),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1092),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1092),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1131),
.B(n_823),
.C(n_822),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1095),
.B(n_733),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1101),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1102),
.Y(n_1165)
);

BUFx2_ASAP7_75t_R g1166 ( 
.A(n_1123),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1088),
.B(n_828),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1094),
.A2(n_902),
.B(n_909),
.C(n_898),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1103),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1128),
.B(n_1114),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1104),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1117),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1091),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1105),
.B(n_1010),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1116),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1115),
.B(n_951),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1115),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1123),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1121),
.B(n_845),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1089),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1119),
.B(n_846),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1089),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1086),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1089),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1090),
.B(n_857),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1119),
.B(n_860),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1119),
.B(n_865),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1089),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1089),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1119),
.B(n_866),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1119),
.B(n_869),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_1093),
.B(n_954),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1090),
.B(n_873),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1122),
.A2(n_963),
.B1(n_967),
.B2(n_962),
.C(n_957),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1090),
.B(n_883),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1093),
.B(n_980),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1093),
.B(n_970),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1090),
.B(n_884),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1118),
.B(n_887),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1112),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1093),
.B(n_733),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1097),
.A2(n_900),
.B1(n_907),
.B2(n_891),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1090),
.A2(n_784),
.B1(n_872),
.B2(n_750),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1086),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1090),
.B(n_912),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1090),
.B(n_913),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1090),
.A2(n_1007),
.B1(n_964),
.B2(n_734),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1090),
.B(n_916),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1089),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1090),
.B(n_922),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1090),
.B(n_926),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1090),
.B(n_927),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1086),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1089),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1119),
.B(n_932),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1090),
.B(n_933),
.Y(n_1216)
);

OAI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1097),
.A2(n_941),
.B1(n_943),
.B2(n_934),
.Y(n_1217)
);

OAI221xp5_ASAP7_75t_L g1218 ( 
.A1(n_1088),
.A2(n_983),
.B1(n_993),
.B2(n_989),
.C(n_974),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1118),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1089),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1086),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1119),
.B(n_1003),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1089),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1119),
.B(n_1006),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1122),
.A2(n_771),
.B1(n_879),
.B2(n_757),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1090),
.B(n_966),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1090),
.B(n_985),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1093),
.B(n_979),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1119),
.B(n_986),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1119),
.B(n_991),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1118),
.B(n_997),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1118),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1119),
.B(n_979),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1147),
.B(n_757),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1138),
.Y(n_1235)
);

NOR2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1133),
.B(n_1132),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1156),
.Y(n_1237)
);

AND2x6_ASAP7_75t_L g1238 ( 
.A(n_1139),
.B(n_728),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1141),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1134),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1173),
.B(n_996),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1178),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1183),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1135),
.B(n_1017),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1204),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1213),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1136),
.B(n_751),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1160),
.B(n_1161),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1178),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1221),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1134),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1166),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1179),
.B(n_999),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1145),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1201),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1148),
.B(n_1185),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1151),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1150),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_L g1259 ( 
.A(n_1193),
.B(n_772),
.C(n_762),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1200),
.B(n_773),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1163),
.A2(n_879),
.B1(n_771),
.B2(n_994),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1192),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1181),
.A2(n_780),
.B(n_781),
.C(n_774),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1228),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1178),
.B(n_783),
.Y(n_1265)
);

AND2x2_ASAP7_75t_SL g1266 ( 
.A(n_1225),
.B(n_724),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1218),
.A2(n_800),
.B1(n_801),
.B2(n_791),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1219),
.B(n_723),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1196),
.B(n_725),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1153),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1169),
.Y(n_1271)
);

NOR2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1197),
.B(n_810),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1195),
.B(n_832),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1198),
.B(n_839),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1232),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1180),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1205),
.B(n_847),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1206),
.A2(n_861),
.B(n_868),
.C(n_856),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1182),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1184),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1137),
.B(n_877),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1208),
.A2(n_906),
.B1(n_908),
.B2(n_895),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1157),
.B(n_0),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1210),
.B(n_919),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1188),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1189),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1209),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1214),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1211),
.B(n_921),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1186),
.B(n_726),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1194),
.A2(n_935),
.B1(n_936),
.B2(n_928),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1212),
.B(n_1216),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1220),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1176),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1223),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1159),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1233),
.B(n_1226),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1227),
.B(n_952),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1176),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1167),
.A2(n_972),
.B1(n_975),
.B2(n_971),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1155),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1187),
.B(n_730),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1158),
.B(n_727),
.Y(n_1303)
);

AND2x2_ASAP7_75t_SL g1304 ( 
.A(n_1207),
.B(n_729),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1144),
.B(n_732),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1190),
.A2(n_914),
.B1(n_945),
.B2(n_840),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1191),
.B(n_735),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1172),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_SL g1309 ( 
.A(n_1203),
.B(n_1222),
.C(n_1215),
.Y(n_1309)
);

NOR2x1_ASAP7_75t_R g1310 ( 
.A(n_1149),
.B(n_1146),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1154),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1224),
.B(n_736),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1164),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1229),
.B(n_738),
.Y(n_1314)
);

NAND2xp33_ASAP7_75t_L g1315 ( 
.A(n_1162),
.B(n_741),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1170),
.A2(n_746),
.B(n_743),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1142),
.B(n_0),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1165),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1230),
.B(n_749),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1140),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1175),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1143),
.B(n_753),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1171),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1152),
.B(n_1),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1199),
.B(n_1009),
.Y(n_1325)
);

NOR3xp33_ASAP7_75t_SL g1326 ( 
.A(n_1202),
.B(n_755),
.C(n_754),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1177),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1217),
.B(n_756),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1168),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1231),
.B(n_759),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1174),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1173),
.B(n_763),
.Y(n_1332)
);

AND2x2_ASAP7_75t_SL g1333 ( 
.A(n_1132),
.B(n_747),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1132),
.B(n_1),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_1179),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1139),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1173),
.B(n_764),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1147),
.B(n_768),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1147),
.B(n_775),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1138),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1132),
.Y(n_1341)
);

NOR3xp33_ASAP7_75t_SL g1342 ( 
.A(n_1149),
.B(n_777),
.C(n_776),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1138),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1147),
.B(n_778),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1138),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1133),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1138),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1173),
.B(n_785),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1147),
.B(n_786),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1139),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1147),
.B(n_2),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1139),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1133),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1173),
.B(n_787),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1132),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1173),
.B(n_788),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1147),
.B(n_789),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1139),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1139),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1147),
.B(n_790),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1133),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_1132),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1133),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1133),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1173),
.B(n_794),
.Y(n_1365)
);

BUFx6f_ASAP7_75t_L g1366 ( 
.A(n_1133),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1173),
.B(n_795),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1139),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1173),
.B(n_799),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1139),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1173),
.B(n_806),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1147),
.B(n_808),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_R g1373 ( 
.A(n_1133),
.B(n_811),
.Y(n_1373)
);

NAND3xp33_ASAP7_75t_SL g1374 ( 
.A(n_1147),
.B(n_814),
.C(n_813),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1138),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1138),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1173),
.B(n_812),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1173),
.B(n_815),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1133),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1179),
.A2(n_769),
.B1(n_890),
.B2(n_747),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1139),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1133),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1173),
.B(n_818),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1163),
.A2(n_819),
.B1(n_821),
.B2(n_820),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_L g1385 ( 
.A1(n_1181),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1335),
.B(n_1012),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1269),
.B(n_1013),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1353),
.Y(n_1388)
);

OAI21xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1298),
.A2(n_12),
.B(n_4),
.Y(n_1389)
);

NAND3xp33_ASAP7_75t_SL g1390 ( 
.A(n_1320),
.B(n_849),
.C(n_831),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1256),
.B(n_824),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1311),
.B(n_5),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1292),
.A2(n_987),
.B(n_981),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1353),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1239),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1297),
.B(n_5),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1254),
.B(n_6),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1296),
.B(n_988),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1361),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1361),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1290),
.A2(n_992),
.B(n_990),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1255),
.B(n_998),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1362),
.B(n_826),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1355),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1363),
.B(n_6),
.Y(n_1405)
);

INVx3_ASAP7_75t_SL g1406 ( 
.A(n_1364),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1294),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1301),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1366),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1366),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1307),
.A2(n_1004),
.B1(n_862),
.B2(n_918),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_SL g1412 ( 
.A1(n_1384),
.A2(n_864),
.B1(n_893),
.B2(n_838),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1247),
.A2(n_890),
.B(n_769),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1262),
.B(n_1272),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1258),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1243),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1319),
.A2(n_830),
.B(n_827),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1302),
.A2(n_1001),
.B1(n_959),
.B2(n_882),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1235),
.Y(n_1419)
);

NAND2xp33_ASAP7_75t_L g1420 ( 
.A(n_1326),
.B(n_834),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1245),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1257),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1246),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1328),
.B(n_973),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1264),
.B(n_835),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1379),
.Y(n_1426)
);

NAND3xp33_ASAP7_75t_SL g1427 ( 
.A(n_1253),
.B(n_1372),
.C(n_1360),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1309),
.B(n_836),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1263),
.A2(n_896),
.B(n_925),
.C(n_858),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1382),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1333),
.B(n_7),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1312),
.A2(n_1015),
.B(n_1014),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1236),
.B(n_1346),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1276),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1341),
.B(n_8),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1299),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1250),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1314),
.A2(n_843),
.B(n_837),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1273),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1334),
.B(n_9),
.Y(n_1440)
);

NAND2x1p5_ASAP7_75t_L g1441 ( 
.A(n_1242),
.B(n_769),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_R g1442 ( 
.A(n_1252),
.B(n_1237),
.Y(n_1442)
);

CKINVDCx6p67_ASAP7_75t_R g1443 ( 
.A(n_1251),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1279),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1280),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1274),
.A2(n_1284),
.B(n_1277),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1282),
.B(n_850),
.C(n_848),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1240),
.B(n_10),
.Y(n_1448)
);

CKINVDCx10_ASAP7_75t_R g1449 ( 
.A(n_1248),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_R g1450 ( 
.A(n_1374),
.B(n_853),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1278),
.A2(n_911),
.B(n_940),
.C(n_880),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1304),
.B(n_855),
.Y(n_1452)
);

INVx5_ASAP7_75t_L g1453 ( 
.A(n_1248),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1242),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1266),
.B(n_859),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1244),
.B(n_11),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1249),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1289),
.A2(n_1018),
.B(n_1011),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1313),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1249),
.B(n_890),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1313),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1271),
.B(n_12),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1241),
.B(n_13),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1317),
.A2(n_961),
.B(n_904),
.C(n_881),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_R g1465 ( 
.A(n_1331),
.B(n_875),
.Y(n_1465)
);

NOR3xp33_ASAP7_75t_SL g1466 ( 
.A(n_1338),
.B(n_889),
.C(n_885),
.Y(n_1466)
);

NAND3xp33_ASAP7_75t_SL g1467 ( 
.A(n_1351),
.B(n_953),
.C(n_929),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_R g1468 ( 
.A(n_1275),
.B(n_901),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_R g1469 ( 
.A(n_1238),
.B(n_910),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1340),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1318),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1339),
.B(n_978),
.Y(n_1472)
);

CKINVDCx8_ASAP7_75t_R g1473 ( 
.A(n_1238),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1283),
.A2(n_984),
.B1(n_939),
.B2(n_920),
.Y(n_1474)
);

AND2x6_ASAP7_75t_L g1475 ( 
.A(n_1336),
.B(n_939),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_R g1476 ( 
.A(n_1238),
.B(n_915),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1322),
.A2(n_1005),
.B(n_930),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1332),
.A2(n_931),
.B(n_924),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1350),
.B(n_1381),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1324),
.A2(n_956),
.B(n_942),
.C(n_948),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1281),
.A2(n_939),
.B1(n_984),
.B2(n_950),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1352),
.B(n_13),
.Y(n_1482)
);

NOR3xp33_ASAP7_75t_SL g1483 ( 
.A(n_1344),
.B(n_960),
.C(n_944),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1358),
.A2(n_356),
.B(n_355),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1260),
.B(n_1265),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1373),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1343),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1345),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1337),
.A2(n_1000),
.B(n_976),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1303),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1234),
.A2(n_1306),
.B(n_1354),
.C(n_1348),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1356),
.A2(n_984),
.B(n_358),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1359),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1493)
);

A2O1A1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1259),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1261),
.B(n_17),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1347),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1365),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1325),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1375),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1367),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1407),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1413),
.A2(n_1385),
.B(n_1370),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1388),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1404),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1485),
.B(n_1414),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1440),
.B(n_1291),
.Y(n_1506)
);

AOI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1446),
.A2(n_1330),
.B(n_1268),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1415),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1490),
.B(n_1368),
.Y(n_1509)
);

AOI221x1_ASAP7_75t_L g1510 ( 
.A1(n_1427),
.A2(n_1305),
.B1(n_1321),
.B2(n_1371),
.C(n_1369),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1436),
.B(n_1377),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1490),
.B(n_1471),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1479),
.B(n_1267),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1395),
.Y(n_1514)
);

AO32x2_ASAP7_75t_L g1515 ( 
.A1(n_1493),
.A2(n_1300),
.A3(n_1329),
.B1(n_1342),
.B2(n_1310),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1452),
.B(n_1378),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1484),
.A2(n_1327),
.B(n_1308),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1459),
.B(n_1453),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1492),
.A2(n_1323),
.B(n_1285),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1482),
.A2(n_1380),
.B(n_1286),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1441),
.A2(n_1491),
.B(n_1421),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1416),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1408),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1423),
.A2(n_1287),
.B(n_1270),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1428),
.A2(n_1383),
.B(n_1357),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1425),
.Y(n_1526)
);

AOI221x1_ASAP7_75t_L g1527 ( 
.A1(n_1494),
.A2(n_1295),
.B1(n_1293),
.B2(n_1288),
.C(n_1316),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1389),
.A2(n_1315),
.B1(n_1349),
.B2(n_1376),
.C(n_22),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1426),
.B(n_20),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1396),
.B(n_1455),
.Y(n_1530)
);

NOR2xp67_ASAP7_75t_L g1531 ( 
.A(n_1453),
.B(n_357),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1498),
.B(n_21),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1394),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1437),
.A2(n_360),
.B(n_359),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1397),
.A2(n_362),
.B(n_361),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1419),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1433),
.B(n_363),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_SL g1538 ( 
.A1(n_1392),
.A2(n_24),
.B(n_23),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1442),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1391),
.A2(n_365),
.B(n_364),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1461),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1422),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1456),
.A2(n_367),
.B(n_366),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1463),
.B(n_21),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1393),
.A2(n_370),
.B(n_369),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1430),
.Y(n_1546)
);

AOI31xp67_ASAP7_75t_L g1547 ( 
.A1(n_1424),
.A2(n_373),
.A3(n_374),
.B(n_371),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1448),
.B(n_25),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1461),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1497),
.A2(n_377),
.B(n_376),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1434),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1400),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1388),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1480),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1409),
.B(n_379),
.Y(n_1555)
);

NAND2xp33_ASAP7_75t_L g1556 ( 
.A(n_1466),
.B(n_26),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1431),
.A2(n_30),
.B(n_31),
.C(n_29),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1500),
.A2(n_381),
.B(n_380),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1468),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1411),
.A2(n_27),
.B(n_29),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1462),
.B(n_31),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1449),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1399),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1429),
.A2(n_383),
.B(n_382),
.Y(n_1564)
);

AO31x2_ASAP7_75t_L g1565 ( 
.A1(n_1451),
.A2(n_386),
.A3(n_387),
.B(n_384),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1403),
.B(n_32),
.Y(n_1566)
);

NOR2xp67_ASAP7_75t_L g1567 ( 
.A(n_1457),
.B(n_1390),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1444),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1439),
.A2(n_390),
.B(n_389),
.Y(n_1569)
);

NOR2xp67_ASAP7_75t_L g1570 ( 
.A(n_1387),
.B(n_391),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1399),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1445),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1470),
.A2(n_395),
.B(n_392),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1464),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1495),
.B(n_36),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1406),
.Y(n_1576)
);

NOR2x1_ASAP7_75t_L g1577 ( 
.A(n_1486),
.B(n_396),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1432),
.A2(n_399),
.B(n_397),
.Y(n_1578)
);

NOR2xp67_ASAP7_75t_SL g1579 ( 
.A(n_1473),
.B(n_1410),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1488),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1496),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1410),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1438),
.A2(n_402),
.B(n_400),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1454),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1499),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1472),
.A2(n_404),
.B(n_403),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1487),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1458),
.A2(n_412),
.B(n_410),
.Y(n_1588)
);

INVx5_ASAP7_75t_L g1589 ( 
.A(n_1460),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1460),
.A2(n_415),
.B(n_414),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1477),
.A2(n_418),
.B(n_417),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1465),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1478),
.A2(n_420),
.B(n_419),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1489),
.A2(n_423),
.B(n_421),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_SL g1595 ( 
.A1(n_1386),
.A2(n_39),
.B(n_36),
.C(n_38),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1454),
.B(n_39),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1418),
.A2(n_40),
.B(n_41),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1487),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1412),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1401),
.A2(n_425),
.B(n_424),
.Y(n_1600)
);

AOI221x1_ASAP7_75t_L g1601 ( 
.A1(n_1467),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.C(n_46),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1469),
.B(n_43),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1476),
.B(n_44),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1443),
.Y(n_1604)
);

AO31x2_ASAP7_75t_L g1605 ( 
.A1(n_1417),
.A2(n_429),
.A3(n_430),
.B(n_428),
.Y(n_1605)
);

AO31x2_ASAP7_75t_L g1606 ( 
.A1(n_1475),
.A2(n_433),
.A3(n_434),
.B(n_431),
.Y(n_1606)
);

INVxp33_ASAP7_75t_L g1607 ( 
.A(n_1405),
.Y(n_1607)
);

BUFx2_ASAP7_75t_R g1608 ( 
.A(n_1398),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1447),
.A2(n_45),
.B(n_47),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_SL g1610 ( 
.A(n_1475),
.B(n_1435),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1475),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1474),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1420),
.A2(n_440),
.B(n_438),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1483),
.B(n_1481),
.Y(n_1614)
);

A2O1A1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1402),
.A2(n_51),
.B(n_52),
.C(n_50),
.Y(n_1615)
);

AO31x2_ASAP7_75t_L g1616 ( 
.A1(n_1450),
.A2(n_443),
.A3(n_446),
.B(n_441),
.Y(n_1616)
);

AO31x2_ASAP7_75t_L g1617 ( 
.A1(n_1446),
.A2(n_448),
.A3(n_450),
.B(n_447),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1485),
.B(n_49),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1427),
.A2(n_53),
.B(n_54),
.C(n_52),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1484),
.A2(n_453),
.B(n_452),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1484),
.A2(n_456),
.B(n_455),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1446),
.A2(n_460),
.B(n_457),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1446),
.A2(n_464),
.B(n_463),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1427),
.A2(n_50),
.B(n_53),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1415),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1446),
.B(n_54),
.Y(n_1626)
);

NAND3x1_ASAP7_75t_L g1627 ( 
.A(n_1431),
.B(n_55),
.C(n_56),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1508),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1625),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1504),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1562),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1523),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1580),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1530),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1536),
.Y(n_1635)
);

AO21x2_ASAP7_75t_L g1636 ( 
.A1(n_1507),
.A2(n_467),
.B(n_466),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1521),
.A2(n_469),
.B(n_468),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1506),
.B(n_57),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1542),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1526),
.B(n_58),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1571),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1510),
.A2(n_58),
.B(n_59),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1505),
.B(n_60),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1512),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1517),
.A2(n_472),
.B(n_471),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1514),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1501),
.Y(n_1647)
);

INVx6_ASAP7_75t_L g1648 ( 
.A(n_1571),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1626),
.A2(n_62),
.B(n_63),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1527),
.A2(n_474),
.B(n_473),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1519),
.A2(n_478),
.B(n_475),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1561),
.B(n_63),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1529),
.A2(n_1516),
.B1(n_1566),
.B2(n_1599),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1620),
.A2(n_480),
.B(n_479),
.Y(n_1654)
);

AO21x2_ASAP7_75t_L g1655 ( 
.A1(n_1525),
.A2(n_482),
.B(n_481),
.Y(n_1655)
);

OAI21x1_ASAP7_75t_L g1656 ( 
.A1(n_1621),
.A2(n_1543),
.B(n_1622),
.Y(n_1656)
);

CKINVDCx14_ASAP7_75t_R g1657 ( 
.A(n_1546),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1560),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1522),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1582),
.Y(n_1660)
);

OR2x6_ASAP7_75t_L g1661 ( 
.A(n_1559),
.B(n_483),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_SL g1662 ( 
.A1(n_1624),
.A2(n_64),
.B(n_65),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1551),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1582),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1623),
.A2(n_1535),
.B(n_1534),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1597),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1511),
.B(n_67),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1568),
.Y(n_1668)
);

OAI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1619),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.C(n_72),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1572),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1548),
.B(n_69),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1544),
.A2(n_1575),
.B1(n_1557),
.B2(n_1513),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1541),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1581),
.Y(n_1674)
);

OA21x2_ASAP7_75t_L g1675 ( 
.A1(n_1550),
.A2(n_1558),
.B(n_1569),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1614),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1589),
.B(n_73),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1573),
.A2(n_486),
.B(n_484),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1509),
.Y(n_1679)
);

INVx2_ASAP7_75t_SL g1680 ( 
.A(n_1503),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1585),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1600),
.A2(n_489),
.B(n_488),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1589),
.B(n_74),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1604),
.B(n_490),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1524),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1518),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1587),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1598),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1617),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1617),
.Y(n_1690)
);

CKINVDCx11_ASAP7_75t_R g1691 ( 
.A(n_1604),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1593),
.A2(n_492),
.B(n_491),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1618),
.B(n_75),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1556),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1538),
.Y(n_1695)
);

OA21x2_ASAP7_75t_L g1696 ( 
.A1(n_1528),
.A2(n_496),
.B(n_494),
.Y(n_1696)
);

NOR2xp67_ASAP7_75t_L g1697 ( 
.A(n_1533),
.B(n_497),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1539),
.B(n_76),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1601),
.B(n_78),
.C(n_79),
.Y(n_1699)
);

NAND2x1p5_ASAP7_75t_L g1700 ( 
.A(n_1579),
.B(n_498),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1596),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1607),
.B(n_78),
.Y(n_1702)
);

CKINVDCx11_ASAP7_75t_R g1703 ( 
.A(n_1592),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1549),
.Y(n_1704)
);

AOI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1502),
.A2(n_501),
.B(n_500),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1563),
.B(n_1553),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1635),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1647),
.B(n_1532),
.Y(n_1708)
);

BUFx12f_ASAP7_75t_L g1709 ( 
.A(n_1691),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1650),
.A2(n_1675),
.B(n_1665),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1638),
.B(n_1515),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1630),
.B(n_1627),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1646),
.B(n_1584),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1659),
.Y(n_1714)
);

O2A1O1Ixp33_ASAP7_75t_L g1715 ( 
.A1(n_1672),
.A2(n_1554),
.B(n_1574),
.C(n_1602),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1653),
.A2(n_1658),
.B1(n_1666),
.B2(n_1694),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1669),
.A2(n_1609),
.B1(n_1615),
.B2(n_1603),
.Y(n_1717)
);

CKINVDCx20_ASAP7_75t_R g1718 ( 
.A(n_1631),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1643),
.B(n_1515),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1628),
.B(n_1576),
.Y(n_1720)
);

AOI21x1_ASAP7_75t_SL g1721 ( 
.A1(n_1698),
.A2(n_1537),
.B(n_1555),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1634),
.A2(n_1612),
.B1(n_1608),
.B2(n_1567),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1699),
.A2(n_1613),
.B(n_1610),
.C(n_1570),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1629),
.B(n_1552),
.Y(n_1724)
);

OA22x2_ASAP7_75t_L g1725 ( 
.A1(n_1661),
.A2(n_1577),
.B1(n_1595),
.B2(n_1616),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1663),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1674),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1639),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1668),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1644),
.B(n_1531),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1701),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_SL g1732 ( 
.A1(n_1640),
.A2(n_1695),
.B(n_1649),
.C(n_1657),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1667),
.B(n_1616),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1673),
.B(n_1611),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1652),
.B(n_1671),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1703),
.Y(n_1736)
);

AOI211xp5_ASAP7_75t_L g1737 ( 
.A1(n_1676),
.A2(n_1540),
.B(n_1586),
.C(n_1591),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1688),
.B(n_1606),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1670),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1662),
.A2(n_1578),
.B(n_1545),
.C(n_1594),
.Y(n_1740)
);

AOI31xp33_ASAP7_75t_L g1741 ( 
.A1(n_1700),
.A2(n_1590),
.A3(n_1588),
.B(n_1611),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1693),
.B(n_79),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1704),
.B(n_80),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1679),
.B(n_80),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1681),
.B(n_1606),
.Y(n_1745)
);

O2A1O1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1677),
.A2(n_1564),
.B(n_1583),
.C(n_1520),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1632),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1633),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1687),
.B(n_81),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1650),
.A2(n_1547),
.B(n_1565),
.Y(n_1750)
);

AOI21x1_ASAP7_75t_SL g1751 ( 
.A1(n_1706),
.A2(n_1565),
.B(n_81),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1685),
.Y(n_1752)
);

BUFx6f_ASAP7_75t_L g1753 ( 
.A(n_1686),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1753),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1720),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1731),
.B(n_1680),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1736),
.B(n_1648),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1714),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1711),
.A2(n_1689),
.B1(n_1690),
.B2(n_1642),
.Y(n_1759)
);

OAI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1750),
.A2(n_1710),
.B(n_1746),
.Y(n_1760)
);

AND2x6_ASAP7_75t_L g1761 ( 
.A(n_1719),
.B(n_1683),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1734),
.B(n_1686),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1709),
.B(n_1661),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1726),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1735),
.B(n_1702),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1739),
.B(n_1660),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1708),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1707),
.Y(n_1768)
);

AO31x2_ASAP7_75t_L g1769 ( 
.A1(n_1717),
.A2(n_1637),
.A3(n_1636),
.B(n_1705),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1712),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1727),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1728),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1713),
.B(n_1664),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1729),
.Y(n_1774)
);

AO21x2_ASAP7_75t_L g1775 ( 
.A1(n_1733),
.A2(n_1655),
.B(n_1656),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1724),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1716),
.A2(n_1715),
.B1(n_1732),
.B2(n_1722),
.C(n_1723),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1752),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1747),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1738),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1753),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1745),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1748),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1730),
.B(n_1684),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1749),
.Y(n_1785)
);

INVxp67_ASAP7_75t_SL g1786 ( 
.A(n_1725),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1744),
.Y(n_1787)
);

AO21x2_ASAP7_75t_L g1788 ( 
.A1(n_1741),
.A2(n_1740),
.B(n_1651),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1743),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1718),
.B(n_1648),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1742),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1737),
.B(n_1641),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1751),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1721),
.B(n_1684),
.Y(n_1794)
);

BUFx2_ASAP7_75t_SL g1795 ( 
.A(n_1718),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1731),
.B(n_1696),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1731),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1707),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1715),
.A2(n_1696),
.B(n_1697),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1731),
.B(n_1637),
.Y(n_1800)
);

OR2x6_ASAP7_75t_L g1801 ( 
.A(n_1709),
.B(n_1645),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1709),
.Y(n_1802)
);

INVx4_ASAP7_75t_L g1803 ( 
.A(n_1709),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1758),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1795),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1783),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_L g1807 ( 
.A(n_1777),
.B(n_1675),
.C(n_1605),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1767),
.B(n_1605),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1763),
.A2(n_1692),
.B1(n_1654),
.B2(n_1682),
.Y(n_1809)
);

INVxp33_ASAP7_75t_L g1810 ( 
.A(n_1790),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1764),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1776),
.B(n_1678),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1771),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1755),
.B(n_82),
.Y(n_1814)
);

INVx3_ASAP7_75t_L g1815 ( 
.A(n_1754),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1770),
.B(n_82),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1765),
.B(n_83),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1797),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1778),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1772),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1774),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1768),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1791),
.B(n_83),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1800),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1798),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1779),
.Y(n_1826)
);

OAI322xp33_ASAP7_75t_L g1827 ( 
.A1(n_1786),
.A2(n_89),
.A3(n_88),
.B1(n_86),
.B2(n_84),
.C1(n_85),
.C2(n_87),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1787),
.B(n_84),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1756),
.Y(n_1829)
);

INVx5_ASAP7_75t_SL g1830 ( 
.A(n_1763),
.Y(n_1830)
);

INVxp67_ASAP7_75t_L g1831 ( 
.A(n_1785),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1773),
.B(n_85),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1802),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1782),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1789),
.B(n_86),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1780),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1754),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1796),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1784),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1789),
.B(n_87),
.Y(n_1840)
);

INVx8_ASAP7_75t_L g1841 ( 
.A(n_1781),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1792),
.B(n_88),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1766),
.B(n_89),
.Y(n_1843)
);

AOI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1759),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1760),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1775),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1793),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1803),
.B(n_91),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1761),
.B(n_92),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1761),
.B(n_93),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1761),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1762),
.B(n_94),
.Y(n_1852)
);

AOI222xp33_ASAP7_75t_L g1853 ( 
.A1(n_1799),
.A2(n_97),
.B1(n_99),
.B2(n_95),
.C1(n_96),
.C2(n_98),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1769),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1788),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1794),
.Y(n_1856)
);

INVx4_ASAP7_75t_L g1857 ( 
.A(n_1801),
.Y(n_1857)
);

AND2x4_ASAP7_75t_SL g1858 ( 
.A(n_1757),
.B(n_96),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1801),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1769),
.B(n_97),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1776),
.B(n_98),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1758),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1776),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1797),
.B(n_99),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1776),
.B(n_100),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1776),
.B(n_100),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1783),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1758),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1776),
.B(n_101),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1758),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1758),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1758),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1756),
.Y(n_1873)
);

NOR2x1_ASAP7_75t_SL g1874 ( 
.A(n_1763),
.B(n_101),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1783),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1776),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1863),
.Y(n_1877)
);

OAI31xp33_ASAP7_75t_L g1878 ( 
.A1(n_1860),
.A2(n_104),
.A3(n_102),
.B(n_103),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1863),
.B(n_102),
.Y(n_1879)
);

AO21x2_ASAP7_75t_L g1880 ( 
.A1(n_1855),
.A2(n_103),
.B(n_104),
.Y(n_1880)
);

AOI22xp33_ASAP7_75t_L g1881 ( 
.A1(n_1853),
.A2(n_1807),
.B1(n_1844),
.B2(n_1856),
.Y(n_1881)
);

OA21x2_ASAP7_75t_L g1882 ( 
.A1(n_1838),
.A2(n_105),
.B(n_106),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1827),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.C(n_108),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1847),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1876),
.B(n_108),
.Y(n_1885)
);

BUFx4f_ASAP7_75t_SL g1886 ( 
.A(n_1833),
.Y(n_1886)
);

AOI221x1_ASAP7_75t_SL g1887 ( 
.A1(n_1848),
.A2(n_112),
.B1(n_109),
.B2(n_110),
.C(n_113),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1806),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1867),
.Y(n_1889)
);

OAI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1849),
.A2(n_113),
.B1(n_109),
.B2(n_112),
.Y(n_1890)
);

AO21x2_ASAP7_75t_L g1891 ( 
.A1(n_1846),
.A2(n_114),
.B(n_115),
.Y(n_1891)
);

OAI33xp33_ASAP7_75t_L g1892 ( 
.A1(n_1831),
.A2(n_116),
.A3(n_119),
.B1(n_114),
.B2(n_115),
.B3(n_117),
.Y(n_1892)
);

OAI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1850),
.A2(n_120),
.B1(n_116),
.B2(n_117),
.C(n_121),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1857),
.B(n_120),
.Y(n_1894)
);

OR2x6_ASAP7_75t_L g1895 ( 
.A(n_1841),
.B(n_121),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1804),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1811),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1813),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1875),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1829),
.B(n_122),
.Y(n_1900)
);

OAI211xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1864),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_1901)
);

OAI211xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1842),
.A2(n_126),
.B(n_123),
.C(n_125),
.Y(n_1902)
);

AOI31xp33_ASAP7_75t_L g1903 ( 
.A1(n_1810),
.A2(n_127),
.A3(n_125),
.B(n_126),
.Y(n_1903)
);

OAI211xp5_ASAP7_75t_L g1904 ( 
.A1(n_1824),
.A2(n_131),
.B(n_128),
.C(n_130),
.Y(n_1904)
);

OA21x2_ASAP7_75t_L g1905 ( 
.A1(n_1845),
.A2(n_128),
.B(n_131),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1819),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1862),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1859),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_1908)
);

AOI31xp33_ASAP7_75t_L g1909 ( 
.A1(n_1805),
.A2(n_135),
.A3(n_133),
.B(n_134),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1822),
.Y(n_1910)
);

NOR4xp25_ASAP7_75t_SL g1911 ( 
.A(n_1824),
.B(n_1851),
.C(n_1836),
.D(n_1818),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1834),
.B(n_1873),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1808),
.B(n_136),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1868),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1830),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1825),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1812),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1870),
.Y(n_1918)
);

OAI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1832),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.C(n_143),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1839),
.B(n_141),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1826),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1871),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1872),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1854),
.A2(n_145),
.B1(n_142),
.B2(n_144),
.C(n_146),
.Y(n_1924)
);

OAI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1861),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1830),
.B(n_147),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1820),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1814),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1821),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1828),
.A2(n_151),
.B1(n_148),
.B2(n_150),
.C(n_152),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1865),
.B(n_150),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1841),
.Y(n_1932)
);

AO21x2_ASAP7_75t_L g1933 ( 
.A1(n_1816),
.A2(n_1874),
.B(n_1840),
.Y(n_1933)
);

OAI332xp33_ASAP7_75t_L g1934 ( 
.A1(n_1852),
.A2(n_156),
.A3(n_155),
.B1(n_153),
.B2(n_157),
.B3(n_151),
.C1(n_152),
.C2(n_154),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1866),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1869),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1835),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1823),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1817),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1809),
.A2(n_1848),
.B1(n_1843),
.B2(n_1858),
.Y(n_1940)
);

NAND4xp75_ASAP7_75t_L g1941 ( 
.A(n_1815),
.B(n_160),
.C(n_158),
.D(n_159),
.Y(n_1941)
);

INVx4_ASAP7_75t_L g1942 ( 
.A(n_1837),
.Y(n_1942)
);

OA21x2_ASAP7_75t_L g1943 ( 
.A1(n_1838),
.A2(n_158),
.B(n_159),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1860),
.A2(n_163),
.B1(n_160),
.B2(n_161),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1853),
.A2(n_161),
.B(n_163),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1804),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1804),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1804),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1804),
.Y(n_1949)
);

OAI31xp33_ASAP7_75t_SL g1950 ( 
.A1(n_1861),
.A2(n_166),
.A3(n_164),
.B(n_165),
.Y(n_1950)
);

INVxp67_ASAP7_75t_L g1951 ( 
.A(n_1863),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1838),
.B(n_164),
.Y(n_1952)
);

AO21x2_ASAP7_75t_L g1953 ( 
.A1(n_1855),
.A2(n_165),
.B(n_167),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1804),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1827),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.C(n_170),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1804),
.Y(n_1956)
);

NOR2x1_ASAP7_75t_L g1957 ( 
.A(n_1863),
.B(n_168),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1804),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_R g1959 ( 
.A(n_1833),
.B(n_169),
.Y(n_1959)
);

INVx3_ASAP7_75t_L g1960 ( 
.A(n_1830),
.Y(n_1960)
);

OAI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1853),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_1961)
);

AOI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1860),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1863),
.B(n_174),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1849),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_1964)
);

AOI211xp5_ASAP7_75t_L g1965 ( 
.A1(n_1827),
.A2(n_183),
.B(n_192),
.C(n_175),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1863),
.B(n_176),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1804),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1863),
.B(n_177),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1884),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1929),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1888),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1933),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1914),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1936),
.B(n_177),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1877),
.B(n_178),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1886),
.Y(n_1976)
);

OR2x2_ASAP7_75t_L g1977 ( 
.A(n_1912),
.B(n_1913),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_178),
.Y(n_1978)
);

AOI21xp33_ASAP7_75t_L g1979 ( 
.A1(n_1950),
.A2(n_179),
.B(n_180),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1896),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1889),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1957),
.A2(n_179),
.B(n_180),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1897),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1898),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1899),
.Y(n_1985)
);

BUFx2_ASAP7_75t_L g1986 ( 
.A(n_1951),
.Y(n_1986)
);

NAND3xp33_ASAP7_75t_SL g1987 ( 
.A(n_1911),
.B(n_181),
.C(n_182),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1906),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1959),
.Y(n_1989)
);

OAI21x1_ASAP7_75t_L g1990 ( 
.A1(n_1952),
.A2(n_181),
.B(n_183),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1879),
.B(n_184),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1907),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1960),
.B(n_184),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1910),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1895),
.Y(n_1995)
);

BUFx2_ASAP7_75t_L g1996 ( 
.A(n_1894),
.Y(n_1996)
);

NAND2x1_ASAP7_75t_L g1997 ( 
.A(n_1963),
.B(n_185),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1916),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1926),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1966),
.B(n_185),
.Y(n_2000)
);

OA21x2_ASAP7_75t_L g2001 ( 
.A1(n_1927),
.A2(n_186),
.B(n_188),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1918),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1921),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1922),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1935),
.B(n_186),
.Y(n_2005)
);

OR2x6_ASAP7_75t_L g2006 ( 
.A(n_1895),
.B(n_188),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1923),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1946),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1932),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1968),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1938),
.B(n_189),
.Y(n_2011)
);

OAI21x1_ASAP7_75t_L g2012 ( 
.A1(n_1940),
.A2(n_1958),
.B(n_1956),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1885),
.Y(n_2013)
);

INVx8_ASAP7_75t_L g2014 ( 
.A(n_1920),
.Y(n_2014)
);

OA21x2_ASAP7_75t_L g2015 ( 
.A1(n_1947),
.A2(n_189),
.B(n_190),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1948),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1949),
.B(n_1954),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1967),
.Y(n_2018)
);

OAI21x1_ASAP7_75t_L g2019 ( 
.A1(n_1882),
.A2(n_191),
.B(n_192),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1882),
.B(n_193),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1943),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1943),
.B(n_193),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1903),
.B(n_194),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1905),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1880),
.B(n_194),
.Y(n_2025)
);

INVx4_ASAP7_75t_L g2026 ( 
.A(n_1900),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1953),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1905),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1939),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_1881),
.B(n_1931),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1917),
.B(n_195),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1891),
.Y(n_2032)
);

OAI21x1_ASAP7_75t_L g2033 ( 
.A1(n_1964),
.A2(n_195),
.B(n_196),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1937),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1944),
.A2(n_197),
.B(n_198),
.Y(n_2035)
);

INVx1_ASAP7_75t_SL g2036 ( 
.A(n_1941),
.Y(n_2036)
);

OR2x6_ASAP7_75t_L g2037 ( 
.A(n_1945),
.B(n_1904),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1928),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1890),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_1915),
.Y(n_2040)
);

INVx4_ASAP7_75t_SL g2041 ( 
.A(n_1909),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1962),
.B(n_199),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1919),
.Y(n_2043)
);

OA21x2_ASAP7_75t_L g2044 ( 
.A1(n_1930),
.A2(n_199),
.B(n_200),
.Y(n_2044)
);

BUFx2_ASAP7_75t_L g2045 ( 
.A(n_1883),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1893),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1924),
.Y(n_2047)
);

INVx4_ASAP7_75t_SL g2048 ( 
.A(n_1887),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1878),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1901),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1902),
.Y(n_2051)
);

OA21x2_ASAP7_75t_L g2052 ( 
.A1(n_1925),
.A2(n_200),
.B(n_201),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1961),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1965),
.Y(n_2054)
);

OAI21x1_ASAP7_75t_L g2055 ( 
.A1(n_1908),
.A2(n_201),
.B(n_202),
.Y(n_2055)
);

OR2x6_ASAP7_75t_L g2056 ( 
.A(n_1934),
.B(n_202),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1892),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1955),
.Y(n_2058)
);

INVx4_ASAP7_75t_SL g2059 ( 
.A(n_1886),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1914),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1914),
.Y(n_2061)
);

BUFx2_ASAP7_75t_L g2062 ( 
.A(n_1933),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1914),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1884),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1884),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1914),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1914),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_1877),
.B(n_203),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1914),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1884),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1960),
.B(n_203),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1886),
.B(n_204),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1914),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1914),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1884),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1960),
.B(n_204),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1884),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1973),
.B(n_205),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1977),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2029),
.B(n_205),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2013),
.B(n_206),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2060),
.B(n_207),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2001),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1976),
.B(n_207),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2008),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2012),
.B(n_208),
.Y(n_2086)
);

OAI322xp33_ASAP7_75t_L g2087 ( 
.A1(n_2054),
.A2(n_213),
.A3(n_212),
.B1(n_210),
.B2(n_208),
.C1(n_209),
.C2(n_211),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2017),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2061),
.B(n_209),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2015),
.Y(n_2090)
);

OR2x2_ASAP7_75t_L g2091 ( 
.A(n_2063),
.B(n_211),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1996),
.B(n_212),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1980),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2028),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1986),
.B(n_213),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2066),
.B(n_214),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2026),
.B(n_214),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_1999),
.B(n_215),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2009),
.B(n_216),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_1989),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1983),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2010),
.B(n_216),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2032),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2067),
.B(n_217),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2069),
.B(n_218),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_2007),
.Y(n_2106)
);

NAND3xp33_ASAP7_75t_L g2107 ( 
.A(n_2045),
.B(n_218),
.C(n_219),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_1972),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2073),
.B(n_220),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2074),
.B(n_220),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_2024),
.B(n_221),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2062),
.B(n_221),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1974),
.B(n_222),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_2016),
.B(n_223),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2018),
.B(n_2021),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2039),
.B(n_224),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1975),
.B(n_225),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_2059),
.B(n_225),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2059),
.B(n_226),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1984),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1988),
.B(n_227),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1992),
.B(n_227),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2002),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2004),
.B(n_2011),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2020),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1995),
.B(n_228),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2022),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2027),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_2014),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1978),
.B(n_228),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1969),
.Y(n_2131)
);

OR2x2_ASAP7_75t_L g2132 ( 
.A(n_1970),
.B(n_229),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2064),
.B(n_229),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2065),
.Y(n_2134)
);

AOI31xp33_ASAP7_75t_L g2135 ( 
.A1(n_1979),
.A2(n_1987),
.A3(n_2023),
.B(n_1982),
.Y(n_2135)
);

NOR2x1_ASAP7_75t_L g2136 ( 
.A(n_2006),
.B(n_230),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2046),
.B(n_230),
.Y(n_2137)
);

OAI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_2057),
.A2(n_2043),
.B1(n_2058),
.B2(n_2047),
.C(n_2037),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2070),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_1995),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2075),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2077),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1971),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2068),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_2014),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_2005),
.B(n_231),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2050),
.B(n_231),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1981),
.Y(n_2148)
);

INVx1_ASAP7_75t_SL g2149 ( 
.A(n_2041),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_1990),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2030),
.B(n_232),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2034),
.B(n_232),
.Y(n_2152)
);

INVx1_ASAP7_75t_SL g2153 ( 
.A(n_2041),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_2036),
.B(n_233),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2051),
.B(n_233),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2076),
.B(n_234),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2040),
.B(n_234),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2025),
.B(n_235),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2019),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2038),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2053),
.B(n_235),
.Y(n_2161)
);

BUFx2_ASAP7_75t_L g2162 ( 
.A(n_2006),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1985),
.Y(n_2163)
);

INVx2_ASAP7_75t_SL g2164 ( 
.A(n_1997),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_R g2165 ( 
.A(n_2072),
.B(n_236),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1994),
.Y(n_2166)
);

INVx1_ASAP7_75t_SL g2167 ( 
.A(n_1991),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1998),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_2049),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2000),
.B(n_237),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_2033),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2003),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1993),
.B(n_237),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2052),
.Y(n_2174)
);

INVx2_ASAP7_75t_SL g2175 ( 
.A(n_2071),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2048),
.B(n_238),
.Y(n_2176)
);

NAND3xp33_ASAP7_75t_L g2177 ( 
.A(n_2037),
.B(n_238),
.C(n_239),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2048),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2031),
.B(n_239),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2044),
.B(n_240),
.Y(n_2180)
);

OR2x2_ASAP7_75t_L g2181 ( 
.A(n_2056),
.B(n_241),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2042),
.B(n_241),
.Y(n_2182)
);

OR2x2_ASAP7_75t_L g2183 ( 
.A(n_2056),
.B(n_242),
.Y(n_2183)
);

AOI22xp33_ASAP7_75t_L g2184 ( 
.A1(n_2035),
.A2(n_2055),
.B1(n_244),
.B2(n_242),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2013),
.B(n_243),
.Y(n_2185)
);

INVx2_ASAP7_75t_SL g2186 ( 
.A(n_2014),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1977),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_2008),
.Y(n_2188)
);

NAND3xp33_ASAP7_75t_L g2189 ( 
.A(n_2045),
.B(n_243),
.C(n_244),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1973),
.B(n_245),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1973),
.B(n_245),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1973),
.B(n_246),
.Y(n_2192)
);

CKINVDCx16_ASAP7_75t_R g2193 ( 
.A(n_1976),
.Y(n_2193)
);

BUFx2_ASAP7_75t_L g2194 ( 
.A(n_1996),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_1999),
.B(n_246),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2008),
.Y(n_2196)
);

OA21x2_ASAP7_75t_L g2197 ( 
.A1(n_1972),
.A2(n_247),
.B(n_248),
.Y(n_2197)
);

NAND3xp33_ASAP7_75t_L g2198 ( 
.A(n_2045),
.B(n_248),
.C(n_249),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2008),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2013),
.B(n_249),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2008),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1973),
.B(n_250),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2013),
.B(n_250),
.Y(n_2203)
);

CKINVDCx16_ASAP7_75t_R g2204 ( 
.A(n_1976),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2008),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_2013),
.B(n_251),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2008),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2013),
.B(n_251),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2008),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2029),
.B(n_252),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1973),
.B(n_252),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2008),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2008),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1977),
.Y(n_2214)
);

AND2x4_ASAP7_75t_L g2215 ( 
.A(n_1999),
.B(n_253),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2008),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1973),
.B(n_253),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2013),
.B(n_254),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2013),
.B(n_255),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2008),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1973),
.B(n_255),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_1999),
.B(n_256),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2013),
.B(n_256),
.Y(n_2223)
);

AOI33xp33_ASAP7_75t_L g2224 ( 
.A1(n_2058),
.A2(n_259),
.A3(n_261),
.B1(n_257),
.B2(n_258),
.B3(n_260),
.Y(n_2224)
);

INVxp67_ASAP7_75t_L g2225 ( 
.A(n_2045),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_1976),
.B(n_257),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2008),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2013),
.B(n_258),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1973),
.B(n_261),
.Y(n_2229)
);

INVx2_ASAP7_75t_SL g2230 ( 
.A(n_2014),
.Y(n_2230)
);

NOR2x1_ASAP7_75t_L g2231 ( 
.A(n_1987),
.B(n_262),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2008),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2013),
.B(n_262),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2013),
.B(n_263),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2013),
.B(n_263),
.Y(n_2235)
);

OR2x2_ASAP7_75t_L g2236 ( 
.A(n_2029),
.B(n_264),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2008),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1977),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2008),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2008),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1977),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1977),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2029),
.B(n_264),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2167),
.B(n_266),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2162),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2093),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2101),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2145),
.B(n_266),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2162),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2194),
.B(n_267),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2129),
.B(n_2186),
.Y(n_2251)
);

INVxp67_ASAP7_75t_SL g2252 ( 
.A(n_2225),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2120),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2112),
.B(n_267),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2123),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2230),
.B(n_268),
.Y(n_2256)
);

NOR3x1_ASAP7_75t_L g2257 ( 
.A(n_2178),
.B(n_2177),
.C(n_2181),
.Y(n_2257)
);

NAND2xp33_ASAP7_75t_SL g2258 ( 
.A(n_2164),
.B(n_268),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2124),
.B(n_269),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2100),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2144),
.B(n_269),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2083),
.B(n_270),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2081),
.B(n_270),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2185),
.B(n_271),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2171),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2200),
.B(n_271),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2079),
.B(n_272),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2188),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2203),
.B(n_272),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2140),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2193),
.B(n_273),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2187),
.B(n_273),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_2204),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2212),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2125),
.Y(n_2275)
);

NOR2x1_ASAP7_75t_L g2276 ( 
.A(n_2136),
.B(n_274),
.Y(n_2276)
);

AND2x4_ASAP7_75t_L g2277 ( 
.A(n_2092),
.B(n_275),
.Y(n_2277)
);

O2A1O1Ixp33_ASAP7_75t_SL g2278 ( 
.A1(n_2183),
.A2(n_277),
.B(n_275),
.C(n_276),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2132),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2090),
.B(n_277),
.Y(n_2280)
);

AOI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2231),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2127),
.Y(n_2282)
);

OR2x2_ASAP7_75t_L g2283 ( 
.A(n_2214),
.B(n_278),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2106),
.Y(n_2284)
);

AND2x4_ASAP7_75t_L g2285 ( 
.A(n_2097),
.B(n_2098),
.Y(n_2285)
);

AOI22xp33_ASAP7_75t_L g2286 ( 
.A1(n_2174),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2133),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2159),
.B(n_281),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2111),
.Y(n_2289)
);

OR2x2_ASAP7_75t_L g2290 ( 
.A(n_2238),
.B(n_282),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2206),
.B(n_282),
.Y(n_2291)
);

INVx2_ASAP7_75t_SL g2292 ( 
.A(n_2118),
.Y(n_2292)
);

INVx1_ASAP7_75t_SL g2293 ( 
.A(n_2149),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2150),
.B(n_2088),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2085),
.Y(n_2295)
);

OAI22xp33_ASAP7_75t_L g2296 ( 
.A1(n_2135),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2196),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2199),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2208),
.B(n_285),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_2241),
.B(n_286),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2201),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2205),
.Y(n_2302)
);

INVx2_ASAP7_75t_SL g2303 ( 
.A(n_2119),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2207),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2209),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2213),
.Y(n_2306)
);

INVxp67_ASAP7_75t_SL g2307 ( 
.A(n_2197),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2114),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2216),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2220),
.Y(n_2310)
);

NOR2x1_ASAP7_75t_L g2311 ( 
.A(n_2176),
.B(n_286),
.Y(n_2311)
);

OR2x2_ASAP7_75t_L g2312 ( 
.A(n_2242),
.B(n_287),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2218),
.B(n_287),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2227),
.B(n_288),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2197),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2115),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2219),
.B(n_288),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2232),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2237),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2239),
.B(n_289),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2153),
.B(n_289),
.Y(n_2321)
);

OR2x2_ASAP7_75t_L g2322 ( 
.A(n_2240),
.B(n_290),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2116),
.B(n_290),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2223),
.B(n_291),
.Y(n_2324)
);

NAND2x1_ASAP7_75t_L g2325 ( 
.A(n_2108),
.B(n_291),
.Y(n_2325)
);

HB1xp67_ASAP7_75t_L g2326 ( 
.A(n_2161),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2103),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2094),
.Y(n_2328)
);

AOI222xp33_ASAP7_75t_L g2329 ( 
.A1(n_2169),
.A2(n_294),
.B1(n_296),
.B2(n_292),
.C1(n_293),
.C2(n_295),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_SL g2330 ( 
.A(n_2084),
.B(n_2226),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2228),
.B(n_292),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2086),
.Y(n_2332)
);

INVx1_ASAP7_75t_SL g2333 ( 
.A(n_2165),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2233),
.B(n_2234),
.Y(n_2334)
);

AND2x4_ASAP7_75t_L g2335 ( 
.A(n_2095),
.B(n_293),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2080),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2160),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2235),
.B(n_294),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2175),
.B(n_295),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2210),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2195),
.B(n_296),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2146),
.B(n_297),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2151),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2180),
.B(n_297),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2236),
.Y(n_2345)
);

HB1xp67_ASAP7_75t_L g2346 ( 
.A(n_2108),
.Y(n_2346)
);

NOR2x1_ASAP7_75t_L g2347 ( 
.A(n_2243),
.B(n_298),
.Y(n_2347)
);

INVxp67_ASAP7_75t_SL g2348 ( 
.A(n_2152),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2102),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2138),
.A2(n_298),
.B(n_299),
.Y(n_2350)
);

OAI21xp33_ASAP7_75t_L g2351 ( 
.A1(n_2224),
.A2(n_300),
.B(n_301),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2157),
.B(n_300),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2121),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2215),
.Y(n_2354)
);

OR2x2_ASAP7_75t_L g2355 ( 
.A(n_2078),
.B(n_302),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2122),
.Y(n_2356)
);

OAI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2107),
.A2(n_303),
.B(n_304),
.Y(n_2357)
);

INVx3_ASAP7_75t_L g2358 ( 
.A(n_2222),
.Y(n_2358)
);

INVx2_ASAP7_75t_SL g2359 ( 
.A(n_2099),
.Y(n_2359)
);

INVxp67_ASAP7_75t_L g2360 ( 
.A(n_2089),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2117),
.B(n_304),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2130),
.B(n_305),
.Y(n_2362)
);

INVx2_ASAP7_75t_SL g2363 ( 
.A(n_2156),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2105),
.B(n_306),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2109),
.B(n_306),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2082),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2245),
.Y(n_2367)
);

INVxp67_ASAP7_75t_L g2368 ( 
.A(n_2330),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_2249),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2307),
.B(n_2147),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2258),
.Y(n_2371)
);

HB1xp67_ASAP7_75t_L g2372 ( 
.A(n_2260),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2275),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2282),
.Y(n_2374)
);

AOI22xp33_ASAP7_75t_L g2375 ( 
.A1(n_2351),
.A2(n_2128),
.B1(n_2134),
.B2(n_2131),
.Y(n_2375)
);

INVx1_ASAP7_75t_SL g2376 ( 
.A(n_2333),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_2273),
.B(n_2113),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_2292),
.B(n_2173),
.Y(n_2378)
);

OR2x2_ASAP7_75t_L g2379 ( 
.A(n_2252),
.B(n_2289),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2293),
.B(n_2190),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2334),
.B(n_2191),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2336),
.B(n_2192),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2326),
.Y(n_2383)
);

AOI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_2315),
.A2(n_2139),
.B1(n_2142),
.B2(n_2141),
.Y(n_2384)
);

AND2x4_ASAP7_75t_SL g2385 ( 
.A(n_2285),
.B(n_2170),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2303),
.B(n_2359),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2358),
.B(n_2202),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2363),
.B(n_2211),
.Y(n_2388)
);

INVx1_ASAP7_75t_SL g2389 ( 
.A(n_2362),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2251),
.B(n_2217),
.Y(n_2390)
);

OR2x2_ASAP7_75t_L g2391 ( 
.A(n_2340),
.B(n_2345),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2276),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2270),
.B(n_2221),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2246),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2325),
.Y(n_2395)
);

INVx2_ASAP7_75t_SL g2396 ( 
.A(n_2335),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2349),
.B(n_2229),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_2346),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2335),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2247),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2271),
.B(n_2091),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_2332),
.B(n_2354),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2267),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2253),
.Y(n_2404)
);

OR2x2_ASAP7_75t_L g2405 ( 
.A(n_2366),
.B(n_2096),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2272),
.Y(n_2406)
);

INVx1_ASAP7_75t_SL g2407 ( 
.A(n_2361),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2255),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2250),
.B(n_2104),
.Y(n_2409)
);

NOR2x1_ASAP7_75t_L g2410 ( 
.A(n_2262),
.B(n_2110),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_2353),
.B(n_2158),
.Y(n_2411)
);

NOR2xp33_ASAP7_75t_L g2412 ( 
.A(n_2360),
.B(n_2155),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2244),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2248),
.B(n_2179),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2327),
.Y(n_2415)
);

OAI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2280),
.A2(n_2189),
.B1(n_2198),
.B2(n_2137),
.Y(n_2416)
);

AOI22xp33_ASAP7_75t_L g2417 ( 
.A1(n_2343),
.A2(n_2143),
.B1(n_2163),
.B2(n_2148),
.Y(n_2417)
);

OR2x2_ASAP7_75t_L g2418 ( 
.A(n_2356),
.B(n_2166),
.Y(n_2418)
);

OAI22xp5_ASAP7_75t_L g2419 ( 
.A1(n_2288),
.A2(n_2154),
.B1(n_2182),
.B2(n_2184),
.Y(n_2419)
);

AOI21xp5_ASAP7_75t_L g2420 ( 
.A1(n_2296),
.A2(n_2350),
.B(n_2278),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2295),
.Y(n_2421)
);

OR2x2_ASAP7_75t_L g2422 ( 
.A(n_2268),
.B(n_2274),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2348),
.B(n_2126),
.Y(n_2423)
);

INVx1_ASAP7_75t_SL g2424 ( 
.A(n_2263),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2259),
.B(n_2168),
.Y(n_2425)
);

INVx1_ASAP7_75t_SL g2426 ( 
.A(n_2264),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2398),
.Y(n_2427)
);

NOR2xp33_ASAP7_75t_R g2428 ( 
.A(n_2376),
.B(n_2256),
.Y(n_2428)
);

NOR2x1_ASAP7_75t_L g2429 ( 
.A(n_2379),
.B(n_2314),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2372),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2424),
.B(n_2347),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2367),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2420),
.A2(n_2311),
.B(n_2344),
.Y(n_2433)
);

INVx1_ASAP7_75t_SL g2434 ( 
.A(n_2385),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2426),
.B(n_2261),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2377),
.B(n_2257),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2371),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2369),
.Y(n_2438)
);

INVxp67_ASAP7_75t_L g2439 ( 
.A(n_2377),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2389),
.B(n_2284),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2407),
.B(n_2281),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2381),
.B(n_2297),
.Y(n_2442)
);

OAI211xp5_ASAP7_75t_SL g2443 ( 
.A1(n_2375),
.A2(n_2370),
.B(n_2392),
.C(n_2383),
.Y(n_2443)
);

OAI21xp33_ASAP7_75t_L g2444 ( 
.A1(n_2402),
.A2(n_2294),
.B(n_2265),
.Y(n_2444)
);

OAI22xp5_ASAP7_75t_SL g2445 ( 
.A1(n_2368),
.A2(n_2321),
.B1(n_2339),
.B2(n_2331),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2419),
.A2(n_2308),
.B1(n_2287),
.B2(n_2279),
.Y(n_2446)
);

INVx1_ASAP7_75t_SL g2447 ( 
.A(n_2414),
.Y(n_2447)
);

AOI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2416),
.A2(n_2328),
.B1(n_2316),
.B2(n_2357),
.Y(n_2448)
);

OAI31xp33_ASAP7_75t_L g2449 ( 
.A1(n_2412),
.A2(n_2283),
.A3(n_2300),
.B(n_2290),
.Y(n_2449)
);

AOI22xp33_ASAP7_75t_L g2450 ( 
.A1(n_2403),
.A2(n_2337),
.B1(n_2172),
.B2(n_2312),
.Y(n_2450)
);

OAI322xp33_ASAP7_75t_L g2451 ( 
.A1(n_2422),
.A2(n_2302),
.A3(n_2301),
.B1(n_2304),
.B2(n_2306),
.C1(n_2305),
.C2(n_2298),
.Y(n_2451)
);

OAI22xp5_ASAP7_75t_L g2452 ( 
.A1(n_2401),
.A2(n_2286),
.B1(n_2322),
.B2(n_2320),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2399),
.Y(n_2453)
);

OAI32xp33_ASAP7_75t_L g2454 ( 
.A1(n_2395),
.A2(n_2254),
.A3(n_2323),
.B1(n_2355),
.B2(n_2338),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2390),
.B(n_2309),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_2378),
.B(n_2277),
.Y(n_2456)
);

AOI21xp33_ASAP7_75t_L g2457 ( 
.A1(n_2391),
.A2(n_2318),
.B(n_2310),
.Y(n_2457)
);

AOI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_2410),
.A2(n_2329),
.B1(n_2266),
.B2(n_2291),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2447),
.Y(n_2459)
);

INVx1_ASAP7_75t_SL g2460 ( 
.A(n_2428),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2442),
.B(n_2409),
.Y(n_2461)
);

NOR3xp33_ASAP7_75t_SL g2462 ( 
.A(n_2443),
.B(n_2387),
.C(n_2374),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2434),
.B(n_2396),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2439),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2430),
.B(n_2405),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2432),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2436),
.B(n_2456),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2455),
.B(n_2386),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2438),
.Y(n_2469)
);

BUFx2_ASAP7_75t_L g2470 ( 
.A(n_2429),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2427),
.Y(n_2471)
);

INVx1_ASAP7_75t_SL g2472 ( 
.A(n_2437),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2440),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_SL g2474 ( 
.A(n_2433),
.B(n_2386),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_2445),
.B(n_2454),
.Y(n_2475)
);

NAND2x1p5_ASAP7_75t_L g2476 ( 
.A(n_2453),
.B(n_2269),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_L g2477 ( 
.A(n_2435),
.B(n_2380),
.Y(n_2477)
);

INVx1_ASAP7_75t_SL g2478 ( 
.A(n_2431),
.Y(n_2478)
);

AOI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2470),
.A2(n_2452),
.B(n_2451),
.Y(n_2479)
);

OAI221xp5_ASAP7_75t_L g2480 ( 
.A1(n_2462),
.A2(n_2458),
.B1(n_2384),
.B2(n_2448),
.C(n_2441),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_SL g2481 ( 
.A(n_2472),
.B(n_2444),
.C(n_2423),
.Y(n_2481)
);

AOI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2478),
.A2(n_2413),
.B1(n_2425),
.B2(n_2406),
.Y(n_2482)
);

AOI222xp33_ASAP7_75t_L g2483 ( 
.A1(n_2475),
.A2(n_2450),
.B1(n_2415),
.B2(n_2373),
.C1(n_2421),
.C2(n_2417),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2460),
.B(n_2411),
.Y(n_2484)
);

AOI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_2474),
.A2(n_2457),
.B(n_2324),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2477),
.A2(n_2393),
.B1(n_2446),
.B2(n_2397),
.Y(n_2486)
);

AOI222xp33_ASAP7_75t_L g2487 ( 
.A1(n_2473),
.A2(n_2404),
.B1(n_2394),
.B2(n_2408),
.C1(n_2400),
.C2(n_2319),
.Y(n_2487)
);

O2A1O1Ixp33_ASAP7_75t_L g2488 ( 
.A1(n_2464),
.A2(n_2352),
.B(n_2365),
.C(n_2364),
.Y(n_2488)
);

XOR2xp5_ASAP7_75t_L g2489 ( 
.A(n_2486),
.B(n_2476),
.Y(n_2489)
);

OAI211xp5_ASAP7_75t_SL g2490 ( 
.A1(n_2479),
.A2(n_2459),
.B(n_2471),
.C(n_2469),
.Y(n_2490)
);

AOI221xp5_ASAP7_75t_L g2491 ( 
.A1(n_2480),
.A2(n_2466),
.B1(n_2461),
.B2(n_2465),
.C(n_2463),
.Y(n_2491)
);

AOI221xp5_ASAP7_75t_L g2492 ( 
.A1(n_2481),
.A2(n_2485),
.B1(n_2488),
.B2(n_2482),
.C(n_2484),
.Y(n_2492)
);

OR2x2_ASAP7_75t_L g2493 ( 
.A(n_2487),
.B(n_2382),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2483),
.A2(n_2468),
.B(n_2467),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2484),
.Y(n_2495)
);

OAI21xp5_ASAP7_75t_L g2496 ( 
.A1(n_2479),
.A2(n_2388),
.B(n_2418),
.Y(n_2496)
);

XNOR2xp5_ASAP7_75t_L g2497 ( 
.A(n_2486),
.B(n_2342),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2495),
.B(n_2449),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2493),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2494),
.B(n_2299),
.Y(n_2500)
);

XOR2x2_ASAP7_75t_L g2501 ( 
.A(n_2497),
.B(n_2313),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2496),
.B(n_2317),
.Y(n_2502)
);

OR2x2_ASAP7_75t_L g2503 ( 
.A(n_2489),
.B(n_2342),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_SL g2504 ( 
.A(n_2492),
.B(n_2087),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2490),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2491),
.B(n_2341),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_SL g2507 ( 
.A(n_2492),
.B(n_307),
.Y(n_2507)
);

NAND2xp33_ASAP7_75t_SL g2508 ( 
.A(n_2495),
.B(n_307),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2495),
.B(n_308),
.Y(n_2509)
);

AND2x4_ASAP7_75t_L g2510 ( 
.A(n_2495),
.B(n_308),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2495),
.B(n_309),
.Y(n_2511)
);

NOR3xp33_ASAP7_75t_L g2512 ( 
.A(n_2492),
.B(n_310),
.C(n_311),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2495),
.B(n_311),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2502),
.B(n_312),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2509),
.Y(n_2515)
);

AOI221xp5_ASAP7_75t_L g2516 ( 
.A1(n_2505),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.C(n_316),
.Y(n_2516)
);

OAI22x1_ASAP7_75t_L g2517 ( 
.A1(n_2499),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2517)
);

OAI221xp5_ASAP7_75t_L g2518 ( 
.A1(n_2504),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.C(n_320),
.Y(n_2518)
);

O2A1O1Ixp33_ASAP7_75t_L g2519 ( 
.A1(n_2507),
.A2(n_321),
.B(n_318),
.C(n_320),
.Y(n_2519)
);

A2O1A1Ixp33_ASAP7_75t_L g2520 ( 
.A1(n_2500),
.A2(n_325),
.B(n_322),
.C(n_324),
.Y(n_2520)
);

NOR3xp33_ASAP7_75t_L g2521 ( 
.A(n_2508),
.B(n_2498),
.C(n_2511),
.Y(n_2521)
);

AOI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_2501),
.A2(n_322),
.B(n_324),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2513),
.B(n_325),
.Y(n_2523)
);

XNOR2x1_ASAP7_75t_L g2524 ( 
.A(n_2503),
.B(n_326),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2514),
.B(n_2512),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_SL g2526 ( 
.A(n_2518),
.B(n_2510),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2517),
.Y(n_2527)
);

AOI221xp5_ASAP7_75t_L g2528 ( 
.A1(n_2521),
.A2(n_2506),
.B1(n_328),
.B2(n_326),
.C(n_327),
.Y(n_2528)
);

OAI21xp5_ASAP7_75t_L g2529 ( 
.A1(n_2522),
.A2(n_327),
.B(n_328),
.Y(n_2529)
);

AND2x2_ASAP7_75t_SL g2530 ( 
.A(n_2515),
.B(n_329),
.Y(n_2530)
);

CKINVDCx20_ASAP7_75t_R g2531 ( 
.A(n_2523),
.Y(n_2531)
);

INVxp67_ASAP7_75t_SL g2532 ( 
.A(n_2527),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2529),
.B(n_2520),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_2528),
.B(n_2516),
.Y(n_2534)
);

INVx3_ASAP7_75t_L g2535 ( 
.A(n_2530),
.Y(n_2535)
);

AND2x4_ASAP7_75t_L g2536 ( 
.A(n_2525),
.B(n_2524),
.Y(n_2536)
);

AOI322xp5_ASAP7_75t_L g2537 ( 
.A1(n_2532),
.A2(n_2531),
.A3(n_2526),
.B1(n_2519),
.B2(n_331),
.C1(n_334),
.C2(n_333),
.Y(n_2537)
);

AOI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_2535),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_2538)
);

XNOR2xp5_ASAP7_75t_L g2539 ( 
.A(n_2536),
.B(n_332),
.Y(n_2539)
);

AOI221xp5_ASAP7_75t_L g2540 ( 
.A1(n_2533),
.A2(n_2534),
.B1(n_336),
.B2(n_332),
.C(n_335),
.Y(n_2540)
);

OAI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2532),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_2541)
);

BUFx2_ASAP7_75t_L g2542 ( 
.A(n_2539),
.Y(n_2542)
);

NAND2xp33_ASAP7_75t_L g2543 ( 
.A(n_2538),
.B(n_337),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2541),
.Y(n_2544)
);

OAI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2540),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_2545)
);

BUFx2_ASAP7_75t_L g2546 ( 
.A(n_2537),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_SL g2547 ( 
.A1(n_2537),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_2547)
);

XNOR2xp5_ASAP7_75t_L g2548 ( 
.A(n_2539),
.B(n_341),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2539),
.Y(n_2549)
);

NOR2x1_ASAP7_75t_L g2550 ( 
.A(n_2541),
.B(n_341),
.Y(n_2550)
);

AO22x2_ASAP7_75t_L g2551 ( 
.A1(n_2539),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2539),
.Y(n_2552)
);

AOI21xp33_ASAP7_75t_L g2553 ( 
.A1(n_2539),
.A2(n_342),
.B(n_343),
.Y(n_2553)
);

OAI221xp5_ASAP7_75t_SL g2554 ( 
.A1(n_2537),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.C(n_347),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2539),
.B(n_347),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2541),
.A2(n_348),
.B(n_349),
.Y(n_2556)
);

OAI22x1_ASAP7_75t_L g2557 ( 
.A1(n_2548),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2543),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_2558)
);

AO22x2_ASAP7_75t_L g2559 ( 
.A1(n_2549),
.A2(n_352),
.B1(n_353),
.B2(n_503),
.Y(n_2559)
);

OAI22x1_ASAP7_75t_L g2560 ( 
.A1(n_2550),
.A2(n_507),
.B1(n_504),
.B2(n_505),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2551),
.B(n_508),
.Y(n_2561)
);

OAI22xp5_ASAP7_75t_SL g2562 ( 
.A1(n_2547),
.A2(n_512),
.B1(n_509),
.B2(n_511),
.Y(n_2562)
);

OAI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2556),
.A2(n_513),
.B(n_514),
.Y(n_2563)
);

AO22x2_ASAP7_75t_L g2564 ( 
.A1(n_2552),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_2564)
);

AOI22xp5_ASAP7_75t_L g2565 ( 
.A1(n_2546),
.A2(n_520),
.B1(n_518),
.B2(n_519),
.Y(n_2565)
);

AOI22xp33_ASAP7_75t_L g2566 ( 
.A1(n_2542),
.A2(n_523),
.B1(n_521),
.B2(n_522),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2551),
.Y(n_2567)
);

OAI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2555),
.A2(n_524),
.B(n_525),
.Y(n_2568)
);

AOI22x1_ASAP7_75t_L g2569 ( 
.A1(n_2544),
.A2(n_532),
.B1(n_529),
.B2(n_530),
.Y(n_2569)
);

AOI211xp5_ASAP7_75t_L g2570 ( 
.A1(n_2554),
.A2(n_2545),
.B(n_2553),
.C(n_535),
.Y(n_2570)
);

XNOR2x1_ASAP7_75t_L g2571 ( 
.A(n_2548),
.B(n_533),
.Y(n_2571)
);

XNOR2x1_ASAP7_75t_L g2572 ( 
.A(n_2548),
.B(n_534),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2567),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_2573)
);

HB1xp67_ASAP7_75t_L g2574 ( 
.A(n_2557),
.Y(n_2574)
);

OAI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2558),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2561),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2570),
.B(n_542),
.Y(n_2577)
);

AOI22x1_ASAP7_75t_L g2578 ( 
.A1(n_2560),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_2578)
);

OAI22x1_ASAP7_75t_L g2579 ( 
.A1(n_2569),
.A2(n_548),
.B1(n_546),
.B2(n_547),
.Y(n_2579)
);

OAI22x1_ASAP7_75t_SL g2580 ( 
.A1(n_2572),
.A2(n_2571),
.B1(n_2562),
.B2(n_2559),
.Y(n_2580)
);

OAI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2563),
.A2(n_549),
.B(n_552),
.Y(n_2581)
);

OAI21xp33_ASAP7_75t_L g2582 ( 
.A1(n_2565),
.A2(n_553),
.B(n_554),
.Y(n_2582)
);

XNOR2x1_ASAP7_75t_L g2583 ( 
.A(n_2559),
.B(n_555),
.Y(n_2583)
);

INVx8_ASAP7_75t_L g2584 ( 
.A(n_2568),
.Y(n_2584)
);

XOR2xp5_ASAP7_75t_L g2585 ( 
.A(n_2564),
.B(n_556),
.Y(n_2585)
);

OAI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_2566),
.A2(n_560),
.B1(n_557),
.B2(n_559),
.Y(n_2586)
);

OAI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2564),
.A2(n_719),
.B1(n_563),
.B2(n_561),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2583),
.Y(n_2588)
);

OR3x1_ASAP7_75t_L g2589 ( 
.A(n_2576),
.B(n_562),
.C(n_564),
.Y(n_2589)
);

AOI221xp5_ASAP7_75t_L g2590 ( 
.A1(n_2574),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.C(n_568),
.Y(n_2590)
);

AOI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2580),
.A2(n_573),
.B1(n_569),
.B2(n_570),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2585),
.Y(n_2592)
);

AOI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2577),
.A2(n_574),
.B(n_575),
.Y(n_2593)
);

AOI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2582),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_2594)
);

BUFx2_ASAP7_75t_L g2595 ( 
.A(n_2581),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2584),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_2596),
.A2(n_2584),
.B1(n_2578),
.B2(n_2579),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2588),
.A2(n_2575),
.B(n_2587),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2592),
.B(n_2573),
.Y(n_2599)
);

AOI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2593),
.A2(n_2586),
.B(n_579),
.Y(n_2600)
);

OR2x2_ASAP7_75t_L g2601 ( 
.A(n_2597),
.B(n_2599),
.Y(n_2601)
);

OR2x6_ASAP7_75t_L g2602 ( 
.A(n_2598),
.B(n_2595),
.Y(n_2602)
);

AO221x2_ASAP7_75t_L g2603 ( 
.A1(n_2601),
.A2(n_2589),
.B1(n_2600),
.B2(n_2591),
.C(n_2590),
.Y(n_2603)
);

OAI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_2603),
.A2(n_2602),
.B1(n_2594),
.B2(n_584),
.Y(n_2604)
);

AOI211xp5_ASAP7_75t_L g2605 ( 
.A1(n_2604),
.A2(n_585),
.B(n_581),
.C(n_583),
.Y(n_2605)
);


endmodule