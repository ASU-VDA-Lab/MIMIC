module fake_jpeg_7413_n_177 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_15),
.B1(n_25),
.B2(n_18),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_56),
.B1(n_38),
.B2(n_19),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_55),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_29),
.B1(n_18),
.B2(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_54),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_25),
.B1(n_29),
.B2(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_31),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_71),
.B1(n_16),
.B2(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_65),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_30),
.C(n_38),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.C(n_66),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_30),
.C(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_42),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_17),
.B(n_24),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_70),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_49),
.B1(n_28),
.B2(n_26),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_77),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_47),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_63),
.B1(n_59),
.B2(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_53),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_70),
.B1(n_60),
.B2(n_61),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_61),
.B1(n_48),
.B2(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_40),
.B1(n_55),
.B2(n_50),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_95),
.B1(n_100),
.B2(n_84),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_39),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_97),
.C(n_80),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_39),
.B(n_41),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_104),
.B(n_90),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_61),
.C(n_39),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_21),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_105),
.B(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_16),
.B1(n_39),
.B2(n_20),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_39),
.B(n_68),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_74),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_116),
.C(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_111),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_117),
.B(n_119),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_103),
.B1(n_99),
.B2(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_123),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_122),
.Y(n_124)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_128),
.B1(n_106),
.B2(n_104),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_136),
.C(n_117),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_76),
.B1(n_96),
.B2(n_75),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_109),
.C(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_112),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_140),
.C(n_145),
.Y(n_149)
);

OA21x2_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_99),
.B(n_100),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_76),
.B1(n_78),
.B2(n_4),
.Y(n_142)
);

XOR2x2_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_2),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_127),
.B1(n_4),
.B2(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_78),
.B1(n_13),
.B2(n_12),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_144),
.A2(n_135),
.B1(n_134),
.B2(n_132),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_10),
.C(n_3),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_2),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_125),
.C(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_153),
.B(n_10),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_125),
.B(n_126),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_145),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_162),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_140),
.C(n_138),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_147),
.C(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_166),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_150),
.B1(n_155),
.B2(n_151),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_170),
.B1(n_8),
.B2(n_3),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_156),
.B1(n_160),
.B2(n_153),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_159),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_164),
.B(n_5),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_174),
.B(n_171),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_169),
.C(n_5),
.Y(n_176)
);

HAxp5_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_8),
.CON(n_177),
.SN(n_177)
);


endmodule