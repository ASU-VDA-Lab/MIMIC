module real_jpeg_30771_n_11 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_107, n_6, n_104, n_106, n_110, n_112, n_7, n_3, n_5, n_4, n_105, n_109, n_1, n_113, n_103, n_11);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_107;
input n_6;
input n_104;
input n_106;
input n_110;
input n_112;
input n_7;
input n_3;
input n_5;
input n_4;
input n_105;
input n_109;
input n_1;
input n_113;
input n_103;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_0),
.B(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_1),
.B(n_89),
.Y(n_88)
);

HAxp5_ASAP7_75t_SL g93 ( 
.A(n_1),
.B(n_94),
.CON(n_93),
.SN(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_3),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_5),
.B(n_10),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_51),
.C(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_7),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_8),
.B(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_9),
.B(n_58),
.Y(n_57)
);

OAI31xp33_ASAP7_75t_L g50 ( 
.A1(n_10),
.A2(n_51),
.A3(n_56),
.B(n_60),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_21),
.Y(n_11)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_103),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_97),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_36),
.B(n_95),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_35),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_88),
.B(n_93),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_46),
.B(n_86),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_45),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_78),
.C(n_79),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_71),
.B(n_77),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_49)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_107),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_109),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_93),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_104),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_105),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_106),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_108),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_110),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_111),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_112),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_113),
.Y(n_90)
);


endmodule