module fake_jpeg_939_n_542 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_542);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_49),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_24),
.B(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_50),
.B(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_56),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_57),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_61),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_16),
.B(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_65),
.B(n_72),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_66),
.Y(n_155)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g156 ( 
.A(n_71),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_16),
.B(n_12),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

CKINVDCx9p33_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_16),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_80),
.B(n_16),
.Y(n_140)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_35),
.B(n_0),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_33),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_99),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_100),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

BUFx4f_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_118),
.B(n_140),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_26),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_123),
.B(n_162),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_26),
.B1(n_48),
.B2(n_22),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_135),
.A2(n_137),
.B1(n_154),
.B2(n_166),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_26),
.B1(n_48),
.B2(n_22),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_59),
.B(n_16),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_38),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_21),
.B1(n_38),
.B2(n_32),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_66),
.B(n_47),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_163),
.Y(n_209)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_69),
.A2(n_45),
.B1(n_44),
.B2(n_43),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_66),
.B(n_19),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_73),
.Y(n_201)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_104),
.B1(n_96),
.B2(n_92),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_172),
.A2(n_176),
.B1(n_208),
.B2(n_214),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_23),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_173),
.B(n_197),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_116),
.A2(n_82),
.B1(n_63),
.B2(n_95),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_178),
.B1(n_187),
.B2(n_195),
.Y(n_235)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_125),
.A2(n_85),
.B1(n_91),
.B2(n_41),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_138),
.B1(n_114),
.B2(n_78),
.Y(n_178)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_188),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_137),
.B1(n_135),
.B2(n_108),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_190),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_114),
.A2(n_84),
.B1(n_64),
.B2(n_89),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_113),
.B(n_32),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_152),
.B(n_32),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_200),
.B(n_201),
.Y(n_246)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_107),
.B(n_71),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_117),
.C(n_165),
.Y(n_231)
);

AO22x2_ASAP7_75t_L g205 ( 
.A1(n_150),
.A2(n_71),
.B1(n_44),
.B2(n_43),
.Y(n_205)
);

OA22x2_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_128),
.B1(n_127),
.B2(n_161),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_106),
.B(n_21),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_23),
.Y(n_252)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_110),
.A2(n_21),
.B1(n_19),
.B2(n_22),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_152),
.B(n_48),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_213),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_211),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_146),
.A2(n_61),
.B1(n_53),
.B2(n_56),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_215),
.B1(n_216),
.B2(n_19),
.Y(n_238)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_151),
.A2(n_30),
.B1(n_45),
.B2(n_44),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_146),
.A2(n_86),
.B1(n_83),
.B2(n_87),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_153),
.A2(n_57),
.B1(n_77),
.B2(n_76),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_148),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_222),
.B(n_171),
.C(n_181),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_192),
.A2(n_145),
.B1(n_164),
.B2(n_159),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_223),
.A2(n_228),
.B1(n_233),
.B2(n_242),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_189),
.A2(n_145),
.B1(n_112),
.B2(n_130),
.Y(n_228)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_205),
.B(n_197),
.C(n_210),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_231),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_188),
.B(n_134),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_245),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_216),
.A2(n_149),
.B1(n_165),
.B2(n_93),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_103),
.B1(n_101),
.B2(n_157),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_179),
.B1(n_195),
.B2(n_178),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_204),
.A2(n_124),
.B1(n_105),
.B2(n_109),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_173),
.B(n_77),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_38),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_255),
.B(n_218),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_257),
.A2(n_259),
.B1(n_272),
.B2(n_273),
.Y(n_301)
);

NAND2x1p5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_204),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_258),
.A2(n_267),
.B(n_284),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_191),
.B1(n_186),
.B2(n_184),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_174),
.B1(n_191),
.B2(n_215),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_260),
.A2(n_274),
.B1(n_275),
.B2(n_277),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_251),
.C(n_247),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_200),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_234),
.A2(n_191),
.B1(n_170),
.B2(n_205),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_266),
.A2(n_249),
.B(n_250),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_205),
.Y(n_267)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_225),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_191),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_278),
.C(n_229),
.Y(n_294)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_235),
.A2(n_153),
.B1(n_144),
.B2(n_142),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_142),
.B1(n_144),
.B2(n_158),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_229),
.A2(n_205),
.B1(n_157),
.B2(n_169),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_243),
.A2(n_209),
.B1(n_175),
.B2(n_177),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_158),
.B1(n_120),
.B2(n_111),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_281),
.B1(n_282),
.B2(n_225),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_227),
.A2(n_209),
.B1(n_213),
.B2(n_199),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_183),
.C(n_182),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_238),
.A2(n_120),
.B1(n_194),
.B2(n_193),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_232),
.A2(n_194),
.B1(n_193),
.B2(n_180),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_227),
.A2(n_199),
.B1(n_203),
.B2(n_171),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_225),
.B1(n_250),
.B2(n_240),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_219),
.A2(n_170),
.B(n_23),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_286),
.A2(n_281),
.B1(n_282),
.B2(n_257),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_240),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_287),
.B(n_289),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_229),
.B1(n_246),
.B2(n_245),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_291),
.A2(n_308),
.B1(n_261),
.B2(n_278),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_300),
.C(n_315),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_218),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_298),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_297),
.A2(n_303),
.B(n_306),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_256),
.B(n_253),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_253),
.C(n_254),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_305),
.B(n_230),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_267),
.A2(n_249),
.B(n_241),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_263),
.A2(n_248),
.B1(n_226),
.B2(n_254),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_272),
.B1(n_276),
.B2(n_269),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_270),
.A2(n_248),
.B1(n_226),
.B2(n_237),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_283),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_310),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_278),
.Y(n_325)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_265),
.Y(n_312)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_241),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_263),
.B1(n_260),
.B2(n_266),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_318),
.A2(n_320),
.B1(n_337),
.B2(n_344),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_266),
.B1(n_274),
.B2(n_259),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_323),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_287),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_317),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_294),
.Y(n_355)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_297),
.A3(n_294),
.B1(n_289),
.B2(n_290),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_311),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_300),
.B1(n_312),
.B2(n_310),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_268),
.Y(n_328)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_328),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_258),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_339),
.C(n_311),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_291),
.A2(n_284),
.B1(n_255),
.B2(n_273),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_230),
.B1(n_239),
.B2(n_224),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_255),
.B(n_262),
.C(n_258),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_313),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_290),
.B(n_258),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_335),
.B(n_300),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_291),
.A2(n_284),
.B1(n_285),
.B2(n_230),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_285),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_340),
.Y(n_362)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_343),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_302),
.A2(n_309),
.B1(n_292),
.B2(n_308),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_345),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_202),
.B(n_207),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_346),
.A2(n_350),
.B(n_322),
.Y(n_376)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_349),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_354),
.B(n_382),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_347),
.C(n_339),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_342),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_356),
.B(n_357),
.Y(n_400)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_338),
.A2(n_308),
.B1(n_314),
.B2(n_316),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_363),
.B1(n_370),
.B2(n_380),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_296),
.Y(n_360)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_361),
.B(n_365),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_338),
.A2(n_316),
.B1(n_303),
.B2(n_306),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_325),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_320),
.A2(n_307),
.B1(n_286),
.B2(n_299),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_369),
.A2(n_371),
.B1(n_76),
.B2(n_37),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_322),
.A2(n_304),
.B1(n_299),
.B2(n_296),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_318),
.A2(n_304),
.B1(n_244),
.B2(n_247),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_342),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_375),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_251),
.Y(n_373)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_319),
.B(n_239),
.Y(n_374)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_244),
.B(n_196),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_377),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_319),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_346),
.A2(n_244),
.B(n_198),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_378),
.B(n_379),
.Y(n_388)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_381),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_327),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_392),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_391),
.B(n_401),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_326),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_331),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_393),
.B(n_413),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_358),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_402),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_332),
.B1(n_337),
.B2(n_344),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_396),
.A2(n_398),
.B1(n_403),
.B2(n_404),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_351),
.A2(n_334),
.B1(n_335),
.B2(n_323),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_328),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_360),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_351),
.A2(n_349),
.B1(n_345),
.B2(n_343),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_351),
.A2(n_341),
.B1(n_336),
.B2(n_330),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_383),
.A2(n_341),
.B1(n_336),
.B2(n_330),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_406),
.A2(n_362),
.B1(n_368),
.B2(n_366),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_354),
.B(n_329),
.C(n_321),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_408),
.C(n_409),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_224),
.C(n_185),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_109),
.C(n_105),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_410),
.A2(n_394),
.B1(n_368),
.B2(n_353),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_31),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_374),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_124),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_376),
.C(n_383),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_417),
.C(n_422),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_363),
.C(n_365),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_418),
.A2(n_426),
.B1(n_430),
.B2(n_438),
.Y(n_449)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_400),
.A2(n_356),
.B(n_372),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_420),
.A2(n_421),
.B(n_411),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_380),
.C(n_379),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_367),
.C(n_352),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_427),
.C(n_435),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_392),
.B(n_377),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_434),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_389),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_367),
.C(n_369),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_397),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_428),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_390),
.A2(n_362),
.B1(n_371),
.B2(n_373),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_433),
.A2(n_388),
.B1(n_398),
.B2(n_403),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_370),
.C(n_378),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_405),
.A2(n_381),
.B1(n_366),
.B2(n_353),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_436),
.A2(n_27),
.B1(n_37),
.B2(n_31),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_437),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_390),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_438)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_431),
.A2(n_411),
.B(n_396),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_444),
.A2(n_447),
.B(n_15),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_416),
.A2(n_406),
.B1(n_404),
.B2(n_408),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_445),
.A2(n_451),
.B1(n_457),
.B2(n_439),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_436),
.A2(n_413),
.B(n_409),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_417),
.A2(n_435),
.B1(n_422),
.B2(n_427),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_414),
.A2(n_412),
.B(n_410),
.Y(n_453)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_453),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_454),
.A2(n_27),
.B1(n_434),
.B2(n_15),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_425),
.B(n_41),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_456),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_37),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_414),
.A2(n_31),
.B1(n_30),
.B2(n_18),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_423),
.B(n_27),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_458),
.B(n_460),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_30),
.C(n_18),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_424),
.B(n_18),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_429),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_444),
.A2(n_438),
.B(n_439),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_471),
.Y(n_497)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_470),
.A2(n_477),
.B1(n_482),
.B2(n_3),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_441),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_472),
.A2(n_455),
.B1(n_446),
.B2(n_460),
.Y(n_488)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_462),
.Y(n_473)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_0),
.Y(n_474)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_SL g475 ( 
.A1(n_449),
.A2(n_440),
.B1(n_448),
.B2(n_454),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_475),
.A2(n_445),
.B1(n_447),
.B2(n_451),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_3),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_0),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_11),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_481),
.Y(n_500)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_479),
.B(n_456),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_3),
.C(n_4),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_442),
.C(n_446),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_11),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_461),
.Y(n_482)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_484),
.B(n_488),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_442),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_490),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_496),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_467),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_11),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_491),
.B(n_499),
.Y(n_513)
);

INVx6_ASAP7_75t_L g492 ( 
.A(n_466),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_5),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_466),
.A2(n_472),
.B1(n_476),
.B2(n_482),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_495),
.A2(n_11),
.B(n_6),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_3),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_498),
.B(n_5),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_463),
.B(n_4),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_486),
.A2(n_480),
.B(n_468),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_502),
.A2(n_488),
.B1(n_514),
.B2(n_485),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_468),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_504),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_477),
.C(n_474),
.Y(n_504)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_505),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_5),
.C(n_6),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_510),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_512),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_487),
.B(n_6),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_6),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_515),
.A2(n_498),
.B(n_496),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_508),
.A2(n_514),
.B1(n_493),
.B2(n_507),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_516),
.B(n_517),
.Y(n_528)
);

AOI21x1_ASAP7_75t_SL g521 ( 
.A1(n_508),
.A2(n_500),
.B(n_494),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_521),
.A2(n_504),
.B(n_509),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_522),
.B(n_524),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_501),
.B(n_10),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_506),
.A2(n_6),
.B(n_7),
.Y(n_525)
);

AO21x1_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_526),
.B(n_513),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_8),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_529),
.A2(n_530),
.B(n_531),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_526),
.A2(n_8),
.B(n_9),
.Y(n_530)
);

AO21x1_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_8),
.B(n_9),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_521),
.A2(n_8),
.B(n_9),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_533),
.A2(n_523),
.B(n_520),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_528),
.B(n_519),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_534),
.A2(n_536),
.B(n_537),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_535),
.B(n_532),
.C(n_9),
.Y(n_538)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_538),
.Y(n_540)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_540),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_541),
.B(n_539),
.Y(n_542)
);


endmodule