module fake_netlist_5_849_n_244 (n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_36, n_25, n_18, n_27, n_42, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_48, n_2, n_31, n_23, n_13, n_3, n_49, n_6, n_39, n_244);

input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_36;
input n_25;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_49;
input n_6;
input n_39;

output n_244;

wire n_137;
wire n_210;
wire n_168;
wire n_164;
wire n_191;
wire n_91;
wire n_208;
wire n_82;
wire n_122;
wire n_194;
wire n_142;
wire n_176;
wire n_214;
wire n_140;
wire n_124;
wire n_86;
wire n_146;
wire n_136;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_237;
wire n_90;
wire n_241;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_226;
wire n_235;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_207;
wire n_240;
wire n_114;
wire n_57;
wire n_96;
wire n_189;
wire n_220;
wire n_165;
wire n_111;
wire n_229;
wire n_108;
wire n_231;
wire n_213;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_197;
wire n_107;
wire n_58;
wire n_69;
wire n_236;
wire n_116;
wire n_195;
wire n_227;
wire n_117;
wire n_233;
wire n_94;
wire n_203;
wire n_205;
wire n_113;
wire n_139;
wire n_123;
wire n_105;
wire n_80;
wire n_179;
wire n_125;
wire n_167;
wire n_128;
wire n_73;
wire n_234;
wire n_92;
wire n_149;
wire n_120;
wire n_232;
wire n_135;
wire n_156;
wire n_126;
wire n_225;
wire n_84;
wire n_202;
wire n_130;
wire n_219;
wire n_157;
wire n_79;
wire n_193;
wire n_131;
wire n_151;
wire n_173;
wire n_192;
wire n_53;
wire n_160;
wire n_198;
wire n_223;
wire n_188;
wire n_190;
wire n_201;
wire n_158;
wire n_224;
wire n_100;
wire n_62;
wire n_138;
wire n_154;
wire n_71;
wire n_228;
wire n_148;
wire n_109;
wire n_112;
wire n_212;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_185;
wire n_183;
wire n_243;
wire n_239;
wire n_175;
wire n_169;
wire n_59;
wire n_133;
wire n_238;
wire n_215;
wire n_55;
wire n_196;
wire n_99;
wire n_211;
wire n_218;
wire n_181;
wire n_54;
wire n_147;
wire n_178;
wire n_221;
wire n_67;
wire n_121;
wire n_242;
wire n_76;
wire n_200;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_161;
wire n_209;
wire n_222;
wire n_230;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_174;
wire n_186;
wire n_199;
wire n_134;
wire n_187;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_166;
wire n_206;
wire n_217;
wire n_171;
wire n_153;
wire n_145;
wire n_204;
wire n_50;
wire n_52;
wire n_88;
wire n_110;
wire n_216;

INVx2_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp67_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_15),
.Y(n_57)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_36),
.Y(n_68)
);

INVxp33_ASAP7_75t_SL g69 ( 
.A(n_18),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_0),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_1),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_3),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_3),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_63),
.B(n_4),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_58),
.A2(n_4),
.B(n_5),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_71),
.C(n_52),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_69),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_69),
.B1(n_68),
.B2(n_61),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_75),
.C(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_68),
.B1(n_61),
.B2(n_54),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_7),
.C(n_14),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_19),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_20),
.B(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_30),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_31),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_33),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_83),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_94),
.C(n_99),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_101),
.B1(n_95),
.B2(n_93),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_101),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_90),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_117),
.B(n_122),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_118),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_105),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_112),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_80),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_99),
.Y(n_151)
);

AND2x4_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_102),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

OR2x6_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_34),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_41),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_42),
.Y(n_157)
);

OAI21x1_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_133),
.B(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_138),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_136),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

AND2x4_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_149),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_149),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

AO21x2_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_158),
.B(n_156),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_157),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_125),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_154),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_154),
.Y(n_182)
);

AO21x2_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_152),
.B(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_154),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_164),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_161),
.B(n_164),
.Y(n_190)
);

AO21x2_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_152),
.B(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_167),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_170),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_128),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_179),
.Y(n_201)
);

NAND2x1p5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_181),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_182),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_180),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_186),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_202),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_191),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_191),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_191),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_207),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_209),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_190),
.Y(n_218)
);

NAND2x1_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_196),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_197),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_218),
.Y(n_227)
);

NAND2x1_ASAP7_75t_SL g228 ( 
.A(n_225),
.B(n_213),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

NAND4xp25_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_224),
.C(n_225),
.D(n_221),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_228),
.B(n_219),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_217),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

AOI221xp5_ASAP7_75t_SL g234 ( 
.A1(n_231),
.A2(n_233),
.B1(n_232),
.B2(n_211),
.C(n_129),
.Y(n_234)
);

AOI211xp5_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_152),
.B(n_184),
.C(n_136),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_235),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_136),
.C(n_186),
.Y(n_237)
);

AOI221xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_136),
.B1(n_183),
.B2(n_130),
.C(n_49),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_183),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_177),
.B1(n_153),
.B2(n_148),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_148),
.B(n_239),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_241),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_243),
.A2(n_242),
.B(n_240),
.Y(n_244)
);


endmodule