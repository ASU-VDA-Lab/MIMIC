module real_jpeg_10559_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_1),
.B(n_13),
.CON(n_12),
.SN(n_12)
);

HAxp5_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_9),
.CON(n_16),
.SN(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_1),
.A2(n_3),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g26 ( 
.A(n_1),
.B(n_3),
.Y(n_26)
);

OA21x2_ASAP7_75t_L g13 ( 
.A1(n_2),
.A2(n_14),
.B(n_15),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_14),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_2),
.A2(n_9),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g9 ( 
.A1(n_4),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_9)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

OAI221xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.C(n_24),
.Y(n_7)
);

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_8)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_20),
.B(n_21),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_20),
.Y(n_21)
);

BUFx24_ASAP7_75t_SL g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx24_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_28),
.B(n_31),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);


endmodule