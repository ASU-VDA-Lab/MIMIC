module fake_jpeg_24006_n_280 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_44),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_20),
.B1(n_33),
.B2(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_49),
.B(n_51),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_20),
.B1(n_17),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_31),
.B1(n_27),
.B2(n_34),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_30),
.B1(n_33),
.B2(n_22),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_44),
.B1(n_30),
.B2(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_57),
.A2(n_71),
.B1(n_72),
.B2(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_59),
.B(n_61),
.Y(n_108)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_63),
.B1(n_18),
.B2(n_26),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_33),
.B1(n_22),
.B2(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_0),
.Y(n_66)
);

NOR2x1_ASAP7_75t_R g97 ( 
.A(n_66),
.B(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_17),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_37),
.Y(n_78)
);

AO22x2_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_21),
.B1(n_27),
.B2(n_32),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_2),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_75),
.A2(n_101),
.B(n_102),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_37),
.C(n_41),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_85),
.B1(n_95),
.B2(n_106),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_91),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_92),
.Y(n_128)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_87),
.Y(n_111)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_41),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_57),
.B1(n_56),
.B2(n_55),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_70),
.B(n_60),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_47),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_105),
.B1(n_79),
.B2(n_83),
.Y(n_114)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_52),
.A2(n_28),
.B1(n_41),
.B2(n_3),
.Y(n_105)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_61),
.B(n_52),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_109),
.A2(n_117),
.B(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_82),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_126),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_80),
.B1(n_96),
.B2(n_104),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_1),
.B(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_77),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_130),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_73),
.B(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_134),
.A2(n_100),
.B1(n_89),
.B2(n_87),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_99),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_91),
.B1(n_106),
.B2(n_95),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_144),
.B1(n_155),
.B2(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_145),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_142),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_92),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_117),
.C(n_112),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_99),
.B1(n_86),
.B2(n_88),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_157),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_76),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_81),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_81),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_151),
.A2(n_159),
.B1(n_129),
.B2(n_115),
.Y(n_167)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_107),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_160),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_88),
.B1(n_96),
.B2(n_90),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_100),
.B1(n_89),
.B2(n_87),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_114),
.A2(n_107),
.B1(n_82),
.B2(n_7),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_163),
.B1(n_129),
.B2(n_115),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_82),
.B1(n_6),
.B2(n_8),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_134),
.B(n_120),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_158),
.B(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_132),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_140),
.B1(n_158),
.B2(n_161),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_190),
.B1(n_155),
.B2(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_177),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_187),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_185),
.C(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_179),
.B(n_180),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_119),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_135),
.B(n_131),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_5),
.B(n_8),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_145),
.A2(n_112),
.B(n_110),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_188),
.B1(n_189),
.B2(n_171),
.Y(n_214)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_195),
.B(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_162),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_201),
.C(n_211),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_166),
.A2(n_151),
.B1(n_137),
.B2(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_166),
.A2(n_159),
.B1(n_160),
.B2(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_115),
.B1(n_154),
.B2(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_122),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_185),
.B(n_16),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_172),
.Y(n_224)
);

OA21x2_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_186),
.B(n_184),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_16),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_5),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_8),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_216),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_223),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_192),
.A2(n_179),
.B1(n_187),
.B2(n_170),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_194),
.B1(n_205),
.B2(n_170),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_224),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_172),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_228),
.C(n_208),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_227),
.A2(n_196),
.B(n_169),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_181),
.C(n_169),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_180),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_234),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_205),
.B1(n_193),
.B2(n_194),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_235),
.B(n_237),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_193),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_241),
.C(n_243),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_186),
.B(n_168),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_199),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_222),
.C(n_221),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_215),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_209),
.B(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_207),
.C(n_211),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

OAI321xp33_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_229),
.A3(n_203),
.B1(n_213),
.B2(n_226),
.C(n_200),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_245),
.B(n_248),
.Y(n_255)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_249),
.B(n_202),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_220),
.C(n_228),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_252),
.C(n_230),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_224),
.C(n_175),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_176),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_247),
.Y(n_258)
);

AOI321xp33_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_237),
.A3(n_236),
.B1(n_230),
.B2(n_238),
.C(n_242),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_259),
.B(n_260),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_262),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_233),
.B1(n_190),
.B2(n_177),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_261),
.A2(n_253),
.B1(n_244),
.B2(n_245),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_191),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_265),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_219),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_173),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_9),
.B(n_10),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_259),
.C(n_175),
.Y(n_270)
);

AOI31xp33_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_191),
.B(n_212),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_13),
.Y(n_275)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_263),
.A3(n_266),
.B1(n_13),
.B2(n_14),
.C1(n_9),
.C2(n_16),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_273),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.C(n_269),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_15),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_SL g279 ( 
.A1(n_278),
.A2(n_276),
.B(n_15),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_279),
.Y(n_280)
);


endmodule