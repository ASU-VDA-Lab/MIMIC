module fake_jpeg_11753_n_336 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_50),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_38),
.Y(n_71)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_0),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_26),
.Y(n_51)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_24),
.B1(n_40),
.B2(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_58),
.A2(n_62),
.B1(n_66),
.B2(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_71),
.Y(n_117)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_21),
.B1(n_33),
.B2(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_24),
.B1(n_40),
.B2(n_33),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_63),
.A2(n_74),
.B1(n_83),
.B2(n_85),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_21),
.B1(n_33),
.B2(n_18),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_18),
.B1(n_31),
.B2(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_35),
.B1(n_32),
.B2(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_90),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_46),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_35),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_22),
.Y(n_112)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_96),
.Y(n_137)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_22),
.B1(n_32),
.B2(n_35),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_58),
.B1(n_66),
.B2(n_23),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_108),
.B(n_112),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_80),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_60),
.B(n_37),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_77),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_78),
.A2(n_32),
.B1(n_36),
.B2(n_34),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_126),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_36),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_29),
.B1(n_34),
.B2(n_37),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_25),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_28),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_75),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_81),
.B(n_26),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_87),
.B(n_81),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_106),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_159),
.B(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_151),
.B1(n_161),
.B2(n_125),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_150),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_69),
.B1(n_99),
.B2(n_67),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_69),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_26),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_156),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_64),
.Y(n_156)
);

BUFx8_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_122),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_164),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_61),
.B(n_87),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_112),
.A2(n_80),
.B1(n_89),
.B2(n_9),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_107),
.B(n_137),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_89),
.B1(n_80),
.B2(n_2),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_163),
.B(n_166),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_7),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_6),
.Y(n_166)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_10),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_11),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_0),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_174),
.Y(n_201)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_126),
.B(n_116),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_126),
.A2(n_10),
.B1(n_15),
.B2(n_3),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_154),
.B1(n_173),
.B2(n_146),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_120),
.B(n_118),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_204),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_185),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_129),
.B(n_111),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_191),
.B1(n_205),
.B2(n_154),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_109),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_198),
.C(n_202),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_186),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_190),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_118),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_130),
.C(n_123),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_126),
.B(n_134),
.C(n_107),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_102),
.C(n_132),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_141),
.A2(n_137),
.B(n_102),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_159),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_13),
.B(n_16),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_147),
.B(n_125),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_207),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_179),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_141),
.B1(n_139),
.B2(n_146),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_151),
.B1(n_161),
.B2(n_144),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_217),
.B1(n_222),
.B2(n_235),
.Y(n_243)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_174),
.B1(n_173),
.B2(n_145),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_224),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_178),
.A2(n_145),
.B1(n_140),
.B2(n_167),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_157),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_202),
.C(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_167),
.B1(n_155),
.B2(n_149),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_155),
.B1(n_106),
.B2(n_110),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_230),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_157),
.B1(n_5),
.B2(n_3),
.Y(n_230)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_178),
.A2(n_157),
.B1(n_11),
.B2(n_4),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_252),
.C(n_227),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_186),
.B(n_203),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_223),
.Y(n_266)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_177),
.C(n_206),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_195),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_257),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_213),
.A2(n_176),
.B(n_190),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_211),
.A2(n_178),
.B1(n_199),
.B2(n_194),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_256),
.A2(n_241),
.B1(n_243),
.B2(n_240),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_254),
.B1(n_250),
.B2(n_242),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_246),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_216),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_230),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_275),
.C(n_255),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_274),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_213),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_272),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_234),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_234),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_221),
.C(n_226),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_288),
.C(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_280),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_273),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_258),
.B1(n_235),
.B2(n_248),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_239),
.B(n_238),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_271),
.C(n_275),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_SL g288 ( 
.A(n_264),
.B(n_250),
.C(n_251),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_243),
.B1(n_220),
.B2(n_256),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_292),
.B1(n_259),
.B2(n_270),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_215),
.B1(n_229),
.B2(n_244),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_284),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_260),
.B(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_290),
.Y(n_312)
);

XOR2x1_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_274),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_239),
.B(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_306),
.B(n_307),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_284),
.C(n_287),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_287),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_298),
.C(n_294),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_292),
.B1(n_236),
.B2(n_238),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_310),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_298),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_187),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_189),
.B(n_196),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_318),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_296),
.B1(n_299),
.B2(n_236),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_249),
.B1(n_228),
.B2(n_212),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_197),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_308),
.B1(n_307),
.B2(n_313),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_327),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_232),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_315),
.C(n_316),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_323),
.B(n_322),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_328),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_317),
.B(n_326),
.Y(n_333)
);

OAI31xp33_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_313),
.A3(n_232),
.B(n_189),
.Y(n_334)
);

AOI21x1_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_193),
.B(n_181),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_181),
.Y(n_336)
);


endmodule