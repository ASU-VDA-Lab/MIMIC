module real_jpeg_4008_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_1),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_1),
.B(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_1),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_1),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_1),
.B(n_84),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_2),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_2),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_2),
.B(n_55),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_2),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_3),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_3),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_3),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_3),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_3),
.B(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_5),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_5),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_5),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_5),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_5),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_5),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_6),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_6),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_6),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_6),
.B(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_9),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_9),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_9),
.B(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_9),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_9),
.B(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_10),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_11),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_11),
.B(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_13),
.Y(n_189)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_14),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_14),
.Y(n_344)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_15),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_15),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_15),
.B(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_222),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_221),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_176),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_19),
.B(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_19),
.B(n_225),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_19),
.B(n_225),
.Y(n_421)
);

FAx1_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_67),
.CI(n_133),
.CON(n_19),
.SN(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_51),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_22),
.B(n_36),
.C(n_51),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_30),
.C(n_34),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_28),
.Y(n_139)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_29),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_29),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_30),
.B(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_33),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_37),
.A2(n_38),
.B1(n_187),
.B2(n_190),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_38),
.B(n_43),
.C(n_50),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_38),
.B(n_103),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_38),
.B(n_103),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g267 ( 
.A(n_40),
.Y(n_267)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_46),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_46),
.Y(n_278)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_47),
.Y(n_239)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_47),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_52),
.B(n_150),
.C(n_154),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_52),
.B(n_58),
.C(n_61),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_52),
.A2(n_65),
.B1(n_150),
.B2(n_391),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_61),
.B1(n_72),
.B2(n_76),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_60),
.A2(n_61),
.B1(n_264),
.B2(n_265),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_72),
.C(n_77),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_61),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_63),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_63),
.Y(n_340)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_63),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_98),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_68),
.B(n_99),
.C(n_121),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_82),
.C(n_96),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_69),
.B(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_77),
.B2(n_81),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_72),
.B(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_72),
.A2(n_76),
.B1(n_245),
.B2(n_246),
.Y(n_364)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_78),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_80),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_82),
.B(n_96),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_93),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_93),
.Y(n_136)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_92),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_92),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_93),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_121),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_112),
.C(n_117),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.C(n_110),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_102),
.A2(n_103),
.B1(n_110),
.B2(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_104),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_105),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_105),
.Y(n_249)
);

OR2x2_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_106),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_108),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_146),
.Y(n_145)
);

OR2x2_ASAP7_75t_SL g182 ( 
.A(n_109),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_109),
.B(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_110),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_112),
.B(n_117),
.Y(n_175)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_129),
.B2(n_131),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_124),
.B(n_129),
.C(n_132),
.Y(n_211)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_129),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_129),
.A2(n_131),
.B1(n_217),
.B2(n_220),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_130),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_157),
.C(n_174),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_134),
.B(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_149),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_135),
.B(n_149),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_137),
.B(n_411),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_145),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_138),
.A2(n_145),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_140),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_144),
.B(n_155),
.Y(n_336)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_150),
.Y(n_391)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_154),
.B(n_390),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_155),
.B(n_343),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_157),
.B(n_174),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_166),
.C(n_171),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_158),
.B(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_158),
.A2(n_159),
.B(n_162),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_166),
.B(n_171),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_172),
.B(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_206),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_191),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_181),
.A2(n_182),
.B1(n_240),
.B2(n_362),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_182),
.B(n_237),
.C(n_240),
.Y(n_236)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_184),
.Y(n_323)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_205),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_255),
.B(n_421),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_226),
.B(n_228),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_230),
.B(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_248),
.C(n_253),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_231),
.B(n_407),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.C(n_243),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_232),
.B(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_236),
.A2(n_243),
.B1(n_244),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_236),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_237),
.B(n_361),
.Y(n_360)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_240),
.Y(n_362)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_248),
.B(n_253),
.Y(n_407)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_402),
.B(n_417),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_382),
.B(n_401),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_355),
.B(n_381),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_315),
.B(n_354),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_298),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_261),
.B(n_298),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_273),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_262),
.B(n_274),
.C(n_284),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_263),
.B(n_269),
.C(n_272),
.Y(n_368)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_284),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.C(n_282),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_276),
.B(n_338),
.Y(n_337)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_300)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_285),
.B(n_289),
.C(n_297),
.Y(n_365)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_287),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_292),
.B1(n_296),
.B2(n_297),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_289),
.Y(n_296)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_314),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_299),
.B(n_351),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_301),
.A2(n_302),
.B1(n_314),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_303),
.A2(n_304),
.B1(n_310),
.B2(n_311),
.Y(n_324)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_348),
.B(n_353),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_334),
.B(n_347),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_325),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_322),
.C(n_324),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_326),
.A2(n_327),
.B1(n_331),
.B2(n_332),
.Y(n_345)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_341),
.B(n_346),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_345),
.Y(n_346)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_350),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_357),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_366),
.B2(n_367),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_358),
.B(n_368),
.C(n_369),
.Y(n_400)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_364),
.C(n_365),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_372),
.B2(n_380),
.Y(n_369)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_370),
.Y(n_380)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_378),
.B2(n_379),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_379),
.C(n_380),
.Y(n_386)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_378),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_400),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_400),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_394),
.B2(n_399),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_395),
.C(n_396),
.Y(n_412)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_389),
.C(n_392),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_392),
.B2(n_393),
.Y(n_387)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_388),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_394),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_413),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_412),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_412),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_409),
.C(n_410),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_413),
.A2(n_419),
.B(n_420),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_415),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);


endmodule