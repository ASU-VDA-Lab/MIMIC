module fake_jpeg_5256_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_31),
.B(n_33),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_19),
.Y(n_60)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_30),
.B1(n_23),
.B2(n_17),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_26),
.B1(n_24),
.B2(n_15),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_32),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_18),
.B1(n_27),
.B2(n_26),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_61),
.B1(n_63),
.B2(n_26),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2x1_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_28),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_27),
.B1(n_15),
.B2(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_27),
.B1(n_19),
.B2(n_30),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_70),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_36),
.B1(n_24),
.B2(n_15),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_77),
.B1(n_54),
.B2(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_39),
.B1(n_36),
.B2(n_37),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_72),
.A2(n_80),
.B1(n_16),
.B2(n_46),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_74),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_83),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_36),
.B1(n_17),
.B2(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_103),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_60),
.B1(n_41),
.B2(n_33),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_95),
.B1(n_96),
.B2(n_85),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_50),
.B1(n_45),
.B2(n_53),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_81),
.C(n_87),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_104),
.C(n_105),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_108),
.B1(n_76),
.B2(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_102),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_64),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_33),
.Y(n_116)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_44),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_44),
.C(n_37),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_31),
.C(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_113),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_53),
.B1(n_51),
.B2(n_62),
.Y(n_108)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_41),
.B(n_51),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_41),
.B(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_40),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_73),
.B1(n_66),
.B2(n_77),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_115),
.B(n_127),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_88),
.B(n_80),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_137),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_118),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_46),
.B1(n_31),
.B2(n_76),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_120),
.A2(n_129),
.B1(n_110),
.B2(n_94),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_122),
.B1(n_91),
.B2(n_93),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_46),
.B1(n_79),
.B2(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_56),
.B(n_21),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_91),
.A2(n_103),
.B(n_90),
.Y(n_127)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_33),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_40),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_40),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_29),
.B(n_40),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_82),
.C(n_59),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_104),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_130),
.C(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_141),
.B(n_144),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_91),
.B1(n_92),
.B2(n_98),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_127),
.B1(n_122),
.B2(n_131),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_107),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_155),
.Y(n_191)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_93),
.B1(n_111),
.B2(n_107),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_160),
.B1(n_132),
.B2(n_139),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_111),
.A3(n_107),
.B1(n_100),
.B2(n_105),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_107),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_156),
.A2(n_158),
.B(n_118),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_111),
.B(n_59),
.C(n_21),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g164 ( 
.A(n_114),
.B(n_65),
.C(n_29),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_21),
.B(n_25),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_125),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_173),
.B(n_178),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_167),
.A2(n_185),
.B1(n_25),
.B2(n_21),
.Y(n_212)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_174),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_179),
.C(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_186),
.B(n_160),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_130),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_130),
.C(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_189),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_135),
.C(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_124),
.Y(n_183)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_125),
.B1(n_124),
.B2(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_84),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_165),
.B1(n_162),
.B2(n_163),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_194),
.B1(n_197),
.B2(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_176),
.B1(n_171),
.B2(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_188),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_207),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_144),
.B1(n_164),
.B2(n_158),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_184),
.A2(n_161),
.B(n_160),
.C(n_158),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_213),
.B1(n_28),
.B2(n_3),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_147),
.B1(n_163),
.B2(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_155),
.B1(n_151),
.B2(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_151),
.B(n_1),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_215),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_128),
.B1(n_94),
.B2(n_56),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_210),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_186),
.B(n_169),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_84),
.B1(n_75),
.B2(n_65),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_65),
.C(n_75),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_178),
.C(n_28),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_28),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_219),
.B1(n_230),
.B2(n_202),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_218),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_180),
.B1(n_191),
.B2(n_167),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_179),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_224),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_182),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_233),
.C(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_178),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_224),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_12),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_196),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_0),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_28),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_213),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_247),
.C(n_2),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_242),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_220),
.B(n_233),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_221),
.A2(n_199),
.B1(n_212),
.B2(n_200),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_248),
.B1(n_2),
.B2(n_3),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_217),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_206),
.B(n_198),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_192),
.B(n_205),
.Y(n_244)
);

XOR2x2_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_205),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_249),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_211),
.C(n_215),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_222),
.A2(n_200),
.B1(n_209),
.B2(n_9),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_28),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_12),
.B(n_11),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_234),
.B(n_8),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_225),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_254),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_267),
.B1(n_8),
.B2(n_11),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_225),
.B(n_229),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_4),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_266),
.C(n_9),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_237),
.B(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_268),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_2),
.C(n_3),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_8),
.B1(n_10),
.B2(n_9),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_242),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_271),
.B(n_275),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_249),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_238),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_246),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_281),
.B(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_262),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_4),
.C(n_5),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_290),
.B1(n_281),
.B2(n_10),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_278),
.C(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_259),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_286),
.A2(n_287),
.B(n_291),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_276),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_295),
.B(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_296),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_10),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_4),
.B(n_5),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_6),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_288),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_299),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_300),
.A2(n_302),
.B(n_303),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_304),
.A2(n_297),
.B(n_301),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_306),
.A2(n_305),
.B(n_7),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_7),
.Y(n_308)
);


endmodule