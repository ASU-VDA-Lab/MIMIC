module real_jpeg_12469_n_17 (n_5, n_4, n_8, n_0, n_12, n_325, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_325;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_28),
.B1(n_30),
.B2(n_44),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_0),
.A2(n_44),
.B1(n_59),
.B2(n_63),
.Y(n_269)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_82),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_59),
.B1(n_63),
.B2(n_82),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_82),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_4),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_37),
.B1(n_59),
.B2(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_51),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_7),
.A2(n_51),
.B1(n_59),
.B2(n_63),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_8),
.A2(n_59),
.B1(n_63),
.B2(n_145),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_145),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_145),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_10),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_111),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_10),
.A2(n_59),
.B1(n_63),
.B2(n_111),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_111),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_11),
.B(n_59),
.C(n_62),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_11),
.B(n_31),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_136),
.B(n_181),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_11),
.A2(n_27),
.B(n_30),
.C(n_208),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_52),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_11),
.B(n_41),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_13),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_13),
.A2(n_59),
.B1(n_63),
.B2(n_177),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_177),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_177),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_74),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_14),
.A2(n_59),
.B1(n_63),
.B2(n_74),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_15),
.B(n_28),
.Y(n_265)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_75),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_31),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_24),
.B(n_215),
.Y(n_229)
);

NOR2x1_ASAP7_75t_R g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_26),
.A2(n_32),
.B(n_165),
.Y(n_208)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g264 ( 
.A1(n_30),
.A2(n_42),
.A3(n_48),
.B1(n_252),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_31),
.B(n_215),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_32),
.A2(n_33),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_33),
.B(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_46),
.B1(n_47),
.B2(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_42),
.A2(n_46),
.B(n_165),
.C(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_45),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_47),
.B1(n_73),
.B2(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_46),
.A2(n_144),
.B(n_146),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_46),
.A2(n_47),
.B1(n_144),
.B2(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_81),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_47),
.B(n_110),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_47),
.A2(n_108),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.C(n_72),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_68),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_80),
.C(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_79),
.B1(n_84),
.B2(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_64),
.B(n_66),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_64),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_57),
.A2(n_64),
.B1(n_104),
.B2(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_57),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_57),
.A2(n_64),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_57),
.A2(n_64),
.B1(n_140),
.B2(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_67),
.B1(n_106),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_58),
.A2(n_176),
.B(n_178),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_58),
.B(n_165),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_58),
.A2(n_178),
.B(n_257),
.Y(n_256)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_59),
.Y(n_63)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_63),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_63),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_64),
.B(n_167),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_69),
.A2(n_71),
.B1(n_86),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_69),
.A2(n_71),
.B1(n_115),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_69),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_69),
.A2(n_71),
.B1(n_228),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_69),
.A2(n_214),
.B(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_71),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_71),
.A2(n_142),
.B(n_229),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.C(n_83),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_76),
.A2(n_80),
.B1(n_119),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_80),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_84),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_153),
.B(n_321),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_148),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_123),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_92),
.B(n_123),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_112),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_113),
.C(n_118),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B(n_107),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_95),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_97),
.B1(n_107),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_98),
.A2(n_99),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_98),
.B(n_182),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_98),
.A2(n_99),
.B1(n_135),
.B2(n_269),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_99),
.B(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_114),
.B(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_117),
.A2(n_164),
.B(n_166),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_117),
.A2(n_166),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_130),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_129),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_130),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_141),
.C(n_143),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_131),
.A2(n_132),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_133),
.A2(n_138),
.B1(n_139),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_133),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_136),
.A2(n_137),
.B1(n_210),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_136),
.A2(n_137),
.B1(n_235),
.B2(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_137),
.A2(n_187),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_137),
.B(n_165),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_137),
.A2(n_195),
.B(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_141),
.B(n_143),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_147),
.B(n_250),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g321 ( 
.A1(n_148),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_149),
.B(n_152),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_315),
.B(n_320),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_303),
.B(n_314),
.Y(n_154)
);

OAI321xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_271),
.A3(n_296),
.B1(n_301),
.B2(n_302),
.C(n_325),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_244),
.B(n_270),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_222),
.B(n_243),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_203),
.B(n_221),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_183),
.B(n_202),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_170),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_161),
.B(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_175),
.C(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_180),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_191),
.B(n_201),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_189),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_196),
.B(n_200),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_193),
.B(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_205),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_216),
.C(n_220),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_209),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_224),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_236),
.B2(n_237),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_239),
.C(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_231),
.C(n_234),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_245),
.B(n_246),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_260),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_261),
.C(n_262),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_259),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_254),
.C(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_286),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_286),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_282),
.C(n_285),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_274),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_281),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_280),
.C(n_281),
.Y(n_295)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_285),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_284),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_295),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_290),
.C(n_295),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_313),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_313),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_308),
.C(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);


endmodule