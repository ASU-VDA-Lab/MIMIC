module real_aes_8784_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g410 ( .A(n_0), .Y(n_410) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_1), .A2(n_126), .B(n_129), .C(n_209), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_2), .A2(n_155), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g459 ( .A(n_3), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_4), .B(n_185), .Y(n_184) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_5), .A2(n_155), .B(n_443), .Y(n_442) );
AND2x6_ASAP7_75t_L g126 ( .A(n_6), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g222 ( .A(n_7), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_8), .B(n_39), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_9), .A2(n_154), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_10), .B(n_138), .Y(n_211) );
INVx1_ASAP7_75t_L g447 ( .A(n_11), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_12), .B(n_179), .Y(n_482) );
INVx1_ASAP7_75t_L g118 ( .A(n_13), .Y(n_118) );
INVx1_ASAP7_75t_L g494 ( .A(n_14), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_15), .A2(n_163), .B(n_244), .C(n_246), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_16), .B(n_185), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_17), .B(n_425), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_18), .B(n_155), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_19), .B(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_20), .A2(n_179), .B(n_230), .C(n_232), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_21), .B(n_185), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_22), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_23), .A2(n_165), .B(n_246), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_24), .B(n_138), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_25), .Y(n_120) );
INVx1_ASAP7_75t_L g192 ( .A(n_26), .Y(n_192) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_27), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_28), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_29), .B(n_138), .Y(n_460) );
INVx1_ASAP7_75t_L g161 ( .A(n_30), .Y(n_161) );
INVx1_ASAP7_75t_L g437 ( .A(n_31), .Y(n_437) );
INVx2_ASAP7_75t_L g124 ( .A(n_32), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_33), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_34), .A2(n_179), .B(n_180), .C(n_182), .Y(n_178) );
INVxp67_ASAP7_75t_L g164 ( .A(n_35), .Y(n_164) );
CKINVDCx14_ASAP7_75t_R g177 ( .A(n_36), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_37), .A2(n_129), .B(n_191), .C(n_195), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_38), .A2(n_126), .B(n_129), .C(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g436 ( .A(n_40), .Y(n_436) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_41), .A2(n_140), .B(n_220), .C(n_221), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_42), .B(n_138), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_43), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_44), .Y(n_157) );
INVx1_ASAP7_75t_L g228 ( .A(n_45), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g438 ( .A(n_46), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_47), .B(n_155), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_48), .A2(n_75), .B1(n_101), .B2(n_698), .C1(n_700), .C2(n_701), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_49), .A2(n_129), .B1(n_232), .B2(n_435), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_50), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_51), .Y(n_456) );
CKINVDCx14_ASAP7_75t_R g218 ( .A(n_52), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_53), .A2(n_182), .B(n_220), .C(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_54), .Y(n_506) );
INVx1_ASAP7_75t_L g444 ( .A(n_55), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_56), .A2(n_99), .B1(n_705), .B2(n_714), .C1(n_723), .C2(n_729), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_56), .A2(n_102), .B1(n_699), .B2(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_56), .Y(n_717) );
INVx1_ASAP7_75t_L g127 ( .A(n_57), .Y(n_127) );
INVx1_ASAP7_75t_L g117 ( .A(n_58), .Y(n_117) );
INVx1_ASAP7_75t_SL g181 ( .A(n_59), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_60), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_61), .B(n_185), .Y(n_234) );
INVx1_ASAP7_75t_L g133 ( .A(n_62), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_SL g424 ( .A1(n_63), .A2(n_182), .B(n_425), .C(n_426), .Y(n_424) );
INVxp67_ASAP7_75t_L g427 ( .A(n_64), .Y(n_427) );
INVx1_ASAP7_75t_L g709 ( .A(n_65), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_66), .A2(n_155), .B(n_217), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_67), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_68), .A2(n_155), .B(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_69), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_70), .Y(n_722) );
INVx1_ASAP7_75t_L g500 ( .A(n_71), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_72), .A2(n_154), .B(n_156), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_73), .Y(n_189) );
INVx1_ASAP7_75t_L g242 ( .A(n_74), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_75), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_76), .A2(n_126), .B(n_129), .C(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_77), .A2(n_155), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g245 ( .A(n_78), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_79), .B(n_162), .Y(n_471) );
INVx2_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
INVx1_ASAP7_75t_L g210 ( .A(n_81), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_82), .B(n_425), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_83), .A2(n_126), .B(n_129), .C(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g408 ( .A(n_84), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g697 ( .A(n_84), .Y(n_697) );
OR2x2_ASAP7_75t_L g713 ( .A(n_84), .B(n_704), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g128 ( .A1(n_85), .A2(n_129), .B(n_132), .C(n_142), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_86), .B(n_147), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_87), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_88), .A2(n_126), .B(n_129), .C(n_480), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_89), .Y(n_486) );
INVx1_ASAP7_75t_L g423 ( .A(n_90), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_91), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_92), .B(n_162), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_93), .B(n_113), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_94), .B(n_113), .Y(n_495) );
INVx2_ASAP7_75t_L g231 ( .A(n_95), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_96), .A2(n_155), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_97), .B(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_408), .B1(n_412), .B2(n_694), .Y(n_101) );
INVx2_ASAP7_75t_L g699 ( .A(n_102), .Y(n_699) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_342), .Y(n_102) );
NAND5xp2_ASAP7_75t_L g103 ( .A(n_104), .B(n_271), .C(n_301), .D(n_322), .E(n_328), .Y(n_103) );
AOI221xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_201), .B1(n_235), .B2(n_237), .C(n_248), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_198), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_170), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_SL g322 ( .A1(n_109), .A2(n_186), .B(n_323), .C(n_326), .Y(n_322) );
AND2x2_ASAP7_75t_L g392 ( .A(n_109), .B(n_187), .Y(n_392) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_148), .Y(n_109) );
AND2x2_ASAP7_75t_L g250 ( .A(n_110), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g254 ( .A(n_110), .B(n_251), .Y(n_254) );
OR2x2_ASAP7_75t_L g280 ( .A(n_110), .B(n_187), .Y(n_280) );
AND2x2_ASAP7_75t_L g282 ( .A(n_110), .B(n_173), .Y(n_282) );
AND2x2_ASAP7_75t_L g300 ( .A(n_110), .B(n_172), .Y(n_300) );
INVx1_ASAP7_75t_L g333 ( .A(n_110), .Y(n_333) );
INVx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g200 ( .A(n_111), .Y(n_200) );
AND2x2_ASAP7_75t_L g236 ( .A(n_111), .B(n_173), .Y(n_236) );
AND2x2_ASAP7_75t_L g389 ( .A(n_111), .B(n_187), .Y(n_389) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_119), .B(n_144), .Y(n_111) );
INVx3_ASAP7_75t_L g185 ( .A(n_112), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_112), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_112), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_SL g473 ( .A(n_112), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_113), .Y(n_174) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_113), .A2(n_421), .B(n_428), .Y(n_420) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_115), .B(n_116), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B(n_128), .Y(n_119) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_121), .A2(n_147), .B(n_189), .C(n_190), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_121), .A2(n_207), .B(n_208), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_121), .A2(n_143), .B1(n_434), .B2(n_438), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_121), .A2(n_456), .B(n_457), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g499 ( .A1(n_121), .A2(n_500), .B(n_501), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g121 ( .A(n_122), .B(n_126), .Y(n_121) );
AND2x4_ASAP7_75t_L g155 ( .A(n_122), .B(n_126), .Y(n_155) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
INVx1_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g130 ( .A(n_124), .Y(n_130) );
INVx1_ASAP7_75t_L g233 ( .A(n_124), .Y(n_233) );
INVx1_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_125), .Y(n_136) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
INVx3_ASAP7_75t_L g163 ( .A(n_125), .Y(n_163) );
INVx1_ASAP7_75t_L g425 ( .A(n_125), .Y(n_425) );
INVx4_ASAP7_75t_SL g143 ( .A(n_126), .Y(n_143) );
BUFx3_ASAP7_75t_L g195 ( .A(n_126), .Y(n_195) );
INVx5_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
AND2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
BUFx3_ASAP7_75t_L g141 ( .A(n_130), .Y(n_141) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B(n_137), .C(n_139), .Y(n_132) );
O2A1O1Ixp5_ASAP7_75t_L g209 ( .A1(n_134), .A2(n_139), .B(n_210), .C(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g435 ( .A1(n_135), .A2(n_136), .B1(n_436), .B2(n_437), .Y(n_435) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx4_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
INVx4_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
INVx2_ASAP7_75t_L g220 ( .A(n_138), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_139), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_139), .A2(n_503), .B(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g246 ( .A(n_141), .Y(n_246) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_SL g156 ( .A1(n_143), .A2(n_157), .B(n_158), .C(n_159), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_143), .A2(n_158), .B(n_177), .C(n_178), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_143), .A2(n_158), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_SL g227 ( .A1(n_143), .A2(n_158), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_143), .A2(n_158), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g422 ( .A1(n_143), .A2(n_158), .B(n_423), .C(n_424), .Y(n_422) );
O2A1O1Ixp33_ASAP7_75t_L g443 ( .A1(n_143), .A2(n_158), .B(n_444), .C(n_445), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_143), .A2(n_158), .B(n_491), .C(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
INVx1_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_146), .A2(n_478), .B(n_485), .Y(n_477) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_147), .A2(n_216), .B(n_223), .Y(n_215) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_147), .A2(n_489), .B(n_495), .Y(n_488) );
AND2x2_ASAP7_75t_L g270 ( .A(n_148), .B(n_171), .Y(n_270) );
OR2x2_ASAP7_75t_L g274 ( .A(n_148), .B(n_187), .Y(n_274) );
AND2x2_ASAP7_75t_L g299 ( .A(n_148), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g346 ( .A(n_148), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_148), .B(n_308), .Y(n_394) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_167), .Y(n_148) );
INVx1_ASAP7_75t_L g252 ( .A(n_149), .Y(n_252) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_149), .A2(n_499), .B(n_505), .Y(n_498) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_SL g467 ( .A1(n_150), .A2(n_468), .B(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_151), .A2(n_433), .B(n_439), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_151), .B(n_440), .Y(n_439) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_151), .A2(n_455), .B(n_462), .Y(n_454) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_153), .A2(n_168), .B(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_160), .B(n_166), .Y(n_159) );
OAI22xp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B1(n_164), .B2(n_165), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_162), .A2(n_192), .B(n_193), .C(n_194), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g458 ( .A1(n_162), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
INVx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_163), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_163), .B(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_163), .B(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_165), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_165), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_165), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g194 ( .A(n_166), .Y(n_194) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI322xp33_ASAP7_75t_L g395 ( .A1(n_170), .A2(n_331), .A3(n_354), .B1(n_375), .B2(n_396), .C1(n_398), .C2(n_399), .Y(n_395) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_171), .B(n_251), .Y(n_398) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_186), .Y(n_171) );
AND2x2_ASAP7_75t_L g199 ( .A(n_172), .B(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g267 ( .A(n_172), .B(n_187), .Y(n_267) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g308 ( .A(n_173), .B(n_187), .Y(n_308) );
AND2x2_ASAP7_75t_L g352 ( .A(n_173), .B(n_186), .Y(n_352) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_184), .Y(n_173) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_174), .A2(n_226), .B(n_234), .Y(n_225) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_174), .A2(n_240), .B(n_247), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_179), .B(n_181), .Y(n_180) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_183), .Y(n_483) );
OA21x2_ASAP7_75t_L g441 ( .A1(n_185), .A2(n_442), .B(n_448), .Y(n_441) );
AND2x2_ASAP7_75t_L g235 ( .A(n_186), .B(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g253 ( .A(n_186), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_186), .B(n_282), .Y(n_406) );
INVx3_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g198 ( .A(n_187), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_187), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g320 ( .A(n_187), .B(n_251), .Y(n_320) );
AND2x2_ASAP7_75t_L g347 ( .A(n_187), .B(n_282), .Y(n_347) );
OR2x2_ASAP7_75t_L g403 ( .A(n_187), .B(n_254), .Y(n_403) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_196), .Y(n_187) );
INVx1_ASAP7_75t_SL g289 ( .A(n_198), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_199), .B(n_320), .Y(n_321) );
AND2x2_ASAP7_75t_L g355 ( .A(n_199), .B(n_345), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_199), .B(n_278), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_199), .B(n_400), .Y(n_399) );
OAI31xp33_ASAP7_75t_L g373 ( .A1(n_201), .A2(n_235), .A3(n_374), .B(n_376), .Y(n_373) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_214), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_202), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g356 ( .A(n_202), .B(n_291), .Y(n_356) );
OR2x2_ASAP7_75t_L g363 ( .A(n_202), .B(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g375 ( .A(n_202), .B(n_264), .Y(n_375) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g309 ( .A(n_203), .B(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g237 ( .A(n_204), .B(n_238), .Y(n_237) );
INVx4_ASAP7_75t_L g258 ( .A(n_204), .Y(n_258) );
AND2x2_ASAP7_75t_L g295 ( .A(n_204), .B(n_239), .Y(n_295) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_212), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_205), .B(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_205), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_205), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g294 ( .A(n_214), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g364 ( .A(n_214), .Y(n_364) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_215), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g264 ( .A(n_215), .B(n_225), .Y(n_264) );
INVx2_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_215), .B(n_225), .Y(n_298) );
AND2x2_ASAP7_75t_L g305 ( .A(n_215), .B(n_261), .Y(n_305) );
BUFx3_ASAP7_75t_L g315 ( .A(n_215), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_215), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g260 ( .A(n_224), .Y(n_260) );
AND2x2_ASAP7_75t_L g268 ( .A(n_224), .B(n_258), .Y(n_268) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g238 ( .A(n_225), .B(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
INVx2_ASAP7_75t_L g461 ( .A(n_232), .Y(n_461) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_SL g275 ( .A(n_236), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_236), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_236), .B(n_345), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_237), .B(n_315), .Y(n_368) );
INVx1_ASAP7_75t_SL g402 ( .A(n_237), .Y(n_402) );
INVx1_ASAP7_75t_SL g310 ( .A(n_238), .Y(n_310) );
INVx1_ASAP7_75t_SL g261 ( .A(n_239), .Y(n_261) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_239), .Y(n_272) );
OR2x2_ASAP7_75t_L g283 ( .A(n_239), .B(n_258), .Y(n_283) );
AND2x2_ASAP7_75t_L g297 ( .A(n_239), .B(n_258), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_239), .B(n_287), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_253), .B(n_255), .C(n_266), .Y(n_248) );
AOI31xp33_ASAP7_75t_L g365 ( .A1(n_249), .A2(n_366), .A3(n_367), .B(n_368), .Y(n_365) );
AND2x2_ASAP7_75t_L g338 ( .A(n_250), .B(n_267), .Y(n_338) );
BUFx3_ASAP7_75t_L g278 ( .A(n_251), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_251), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g314 ( .A(n_251), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_251), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g269 ( .A(n_254), .Y(n_269) );
OAI222xp33_ASAP7_75t_L g378 ( .A1(n_254), .A2(n_379), .B1(n_382), .B2(n_383), .C1(n_384), .C2(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_262), .Y(n_255) );
INVx1_ASAP7_75t_L g384 ( .A(n_256), .Y(n_384) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_258), .B(n_261), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_258), .B(n_284), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_258), .B(n_259), .Y(n_354) );
INVx1_ASAP7_75t_L g405 ( .A(n_258), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_259), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g407 ( .A(n_259), .Y(n_407) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g287 ( .A(n_260), .Y(n_287) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_261), .Y(n_330) );
AOI32xp33_ASAP7_75t_L g266 ( .A1(n_262), .A2(n_267), .A3(n_268), .B1(n_269), .B2(n_270), .Y(n_266) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_264), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g341 ( .A(n_264), .Y(n_341) );
OR2x2_ASAP7_75t_L g382 ( .A(n_264), .B(n_283), .Y(n_382) );
INVx1_ASAP7_75t_L g318 ( .A(n_265), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_267), .B(n_278), .Y(n_303) );
INVx3_ASAP7_75t_L g312 ( .A(n_267), .Y(n_312) );
AOI322xp5_ASAP7_75t_L g328 ( .A1(n_267), .A2(n_312), .A3(n_329), .B1(n_331), .B2(n_334), .C1(n_338), .C2(n_339), .Y(n_328) );
AND2x2_ASAP7_75t_L g304 ( .A(n_268), .B(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_L g381 ( .A(n_268), .Y(n_381) );
A2O1A1O1Ixp25_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B(n_276), .C(n_284), .D(n_285), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_272), .B(n_315), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OAI221xp5_ASAP7_75t_L g285 ( .A1(n_274), .A2(n_286), .B1(n_289), .B2(n_290), .C(n_293), .Y(n_285) );
INVx1_ASAP7_75t_SL g400 ( .A(n_274), .Y(n_400) );
AOI21xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B(n_283), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_278), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI221xp5_ASAP7_75t_SL g370 ( .A1(n_280), .A2(n_364), .B1(n_371), .B2(n_372), .C(n_373), .Y(n_370) );
OAI222xp33_ASAP7_75t_L g401 ( .A1(n_281), .A2(n_402), .B1(n_403), .B2(n_404), .C1(n_406), .C2(n_407), .Y(n_401) );
AND2x2_ASAP7_75t_L g359 ( .A(n_282), .B(n_345), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_282), .A2(n_297), .B(n_344), .Y(n_371) );
INVx1_ASAP7_75t_L g385 ( .A(n_282), .Y(n_385) );
INVx2_ASAP7_75t_SL g288 ( .A(n_283), .Y(n_288) );
AND2x2_ASAP7_75t_L g291 ( .A(n_284), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_SL g325 ( .A(n_287), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_287), .B(n_297), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_288), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_288), .B(n_298), .Y(n_327) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21xp5_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_296), .B(n_299), .Y(n_293) );
INVx1_ASAP7_75t_SL g311 ( .A(n_295), .Y(n_311) );
AND2x2_ASAP7_75t_L g358 ( .A(n_295), .B(n_341), .Y(n_358) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g397 ( .A(n_297), .B(n_315), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_298), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g383 ( .A(n_299), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_304), .B1(n_306), .B2(n_313), .C(n_316), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B1(n_311), .B2(n_312), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_310), .A2(n_317), .B1(n_319), .B2(n_321), .Y(n_316) );
OR2x2_ASAP7_75t_L g387 ( .A(n_311), .B(n_315), .Y(n_387) );
OR2x2_ASAP7_75t_L g390 ( .A(n_311), .B(n_325), .Y(n_390) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_332), .A2(n_387), .B1(n_388), .B2(n_390), .C(n_391), .Y(n_386) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND3xp33_ASAP7_75t_SL g342 ( .A(n_343), .B(n_357), .C(n_369), .Y(n_342) );
AOI222xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_348), .B1(n_350), .B2(n_353), .C1(n_355), .C2(n_356), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_345), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g367 ( .A(n_347), .Y(n_367) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_360), .B2(n_362), .C(n_365), .Y(n_357) );
INVx1_ASAP7_75t_L g372 ( .A(n_358), .Y(n_372) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp33_ASAP7_75t_L g391 ( .A1(n_362), .A2(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NOR5xp2_ASAP7_75t_L g369 ( .A(n_370), .B(n_378), .C(n_386), .D(n_395), .E(n_401), .Y(n_369) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_SL g698 ( .A1(n_408), .A2(n_413), .B1(n_694), .B2(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g696 ( .A(n_409), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g704 ( .A(n_409), .Y(n_704) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_SL g413 ( .A(n_414), .B(n_631), .Y(n_413) );
NOR4xp25_ASAP7_75t_L g414 ( .A(n_415), .B(n_561), .C(n_592), .D(n_611), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g415 ( .A(n_416), .B(n_519), .C(n_534), .D(n_552), .Y(n_415) );
AOI222xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_464), .B1(n_496), .B2(n_507), .C1(n_512), .C2(n_514), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_449), .Y(n_417) );
INVx1_ASAP7_75t_L g575 ( .A(n_418), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_429), .Y(n_418) );
AND2x2_ASAP7_75t_L g450 ( .A(n_419), .B(n_441), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_419), .B(n_453), .Y(n_604) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g511 ( .A(n_420), .B(n_431), .Y(n_511) );
AND2x2_ASAP7_75t_L g520 ( .A(n_420), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g546 ( .A(n_420), .Y(n_546) );
AND2x2_ASAP7_75t_L g567 ( .A(n_420), .B(n_431), .Y(n_567) );
BUFx2_ASAP7_75t_L g590 ( .A(n_420), .Y(n_590) );
AND2x2_ASAP7_75t_L g614 ( .A(n_420), .B(n_432), .Y(n_614) );
AND2x2_ASAP7_75t_L g678 ( .A(n_420), .B(n_441), .Y(n_678) );
AND2x2_ASAP7_75t_L g579 ( .A(n_429), .B(n_510), .Y(n_579) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_430), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_441), .Y(n_430) );
OR2x2_ASAP7_75t_L g539 ( .A(n_431), .B(n_454), .Y(n_539) );
AND2x2_ASAP7_75t_L g551 ( .A(n_431), .B(n_510), .Y(n_551) );
BUFx2_ASAP7_75t_L g683 ( .A(n_431), .Y(n_683) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g452 ( .A(n_432), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g533 ( .A(n_432), .B(n_454), .Y(n_533) );
AND2x2_ASAP7_75t_L g586 ( .A(n_432), .B(n_441), .Y(n_586) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_432), .Y(n_622) );
AND2x2_ASAP7_75t_L g509 ( .A(n_441), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_SL g521 ( .A(n_441), .Y(n_521) );
INVx2_ASAP7_75t_L g532 ( .A(n_441), .Y(n_532) );
BUFx2_ASAP7_75t_L g556 ( .A(n_441), .Y(n_556) );
AND2x2_ASAP7_75t_SL g613 ( .A(n_441), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AOI332xp33_ASAP7_75t_L g534 ( .A1(n_450), .A2(n_535), .A3(n_539), .B1(n_540), .B2(n_544), .B3(n_547), .C1(n_548), .C2(n_550), .Y(n_534) );
NAND2x1_ASAP7_75t_L g619 ( .A(n_450), .B(n_510), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_450), .B(n_524), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_SL g552 ( .A1(n_451), .A2(n_553), .B(n_556), .C(n_557), .Y(n_552) );
AND2x2_ASAP7_75t_L g691 ( .A(n_451), .B(n_532), .Y(n_691) );
INVx3_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g588 ( .A(n_452), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g593 ( .A(n_452), .B(n_590), .Y(n_593) );
INVx1_ASAP7_75t_L g524 ( .A(n_453), .Y(n_524) );
AND2x2_ASAP7_75t_L g627 ( .A(n_453), .B(n_586), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_453), .B(n_567), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_453), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_453), .B(n_545), .Y(n_653) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g510 ( .A(n_454), .Y(n_510) );
OAI31xp33_ASAP7_75t_L g692 ( .A1(n_464), .A2(n_613), .A3(n_620), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
AND2x2_ASAP7_75t_L g496 ( .A(n_465), .B(n_497), .Y(n_496) );
NAND2x1_ASAP7_75t_SL g515 ( .A(n_465), .B(n_516), .Y(n_515) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_465), .Y(n_602) );
AND2x2_ASAP7_75t_L g607 ( .A(n_465), .B(n_518), .Y(n_607) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_466), .A2(n_520), .B(n_522), .C(n_525), .Y(n_519) );
OR2x2_ASAP7_75t_L g536 ( .A(n_466), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g549 ( .A(n_466), .Y(n_549) );
AND2x2_ASAP7_75t_L g555 ( .A(n_466), .B(n_498), .Y(n_555) );
INVx2_ASAP7_75t_L g573 ( .A(n_466), .Y(n_573) );
AND2x2_ASAP7_75t_L g584 ( .A(n_466), .B(n_538), .Y(n_584) );
AND2x2_ASAP7_75t_L g616 ( .A(n_466), .B(n_574), .Y(n_616) );
AND2x2_ASAP7_75t_L g620 ( .A(n_466), .B(n_543), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_466), .B(n_475), .Y(n_625) );
AND2x2_ASAP7_75t_L g659 ( .A(n_466), .B(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_466), .B(n_562), .Y(n_693) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_473), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_475), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g601 ( .A(n_475), .Y(n_601) );
AND2x2_ASAP7_75t_L g663 ( .A(n_475), .B(n_584), .Y(n_663) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_487), .Y(n_475) );
OR2x2_ASAP7_75t_L g517 ( .A(n_476), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g527 ( .A(n_476), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_476), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g635 ( .A(n_476), .Y(n_635) );
AND2x2_ASAP7_75t_L g652 ( .A(n_476), .B(n_498), .Y(n_652) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_487), .Y(n_543) );
AND2x2_ASAP7_75t_L g572 ( .A(n_477), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g583 ( .A(n_477), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_477), .B(n_538), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_484), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_483), .Y(n_480) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g497 ( .A(n_488), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g518 ( .A(n_488), .Y(n_518) );
AND2x2_ASAP7_75t_L g574 ( .A(n_488), .B(n_538), .Y(n_574) );
INVx1_ASAP7_75t_L g676 ( .A(n_496), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_497), .Y(n_680) );
INVx2_ASAP7_75t_L g538 ( .A(n_498), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_509), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_509), .B(n_614), .Y(n_672) );
OR2x2_ASAP7_75t_L g513 ( .A(n_510), .B(n_511), .Y(n_513) );
INVx1_ASAP7_75t_SL g565 ( .A(n_510), .Y(n_565) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_516), .A2(n_569), .B1(n_571), .B2(n_575), .C(n_576), .Y(n_568) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g596 ( .A(n_517), .B(n_560), .Y(n_596) );
INVx2_ASAP7_75t_L g528 ( .A(n_518), .Y(n_528) );
INVx1_ASAP7_75t_L g554 ( .A(n_518), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_518), .B(n_538), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_518), .B(n_541), .Y(n_648) );
INVx1_ASAP7_75t_L g656 ( .A(n_518), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_520), .B(n_524), .Y(n_570) );
AND2x4_ASAP7_75t_L g545 ( .A(n_521), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g658 ( .A(n_524), .B(n_614), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_527), .B(n_559), .Y(n_558) );
INVxp67_ASAP7_75t_L g666 ( .A(n_528), .Y(n_666) );
INVxp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g566 ( .A(n_532), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g638 ( .A(n_532), .B(n_614), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_532), .B(n_551), .Y(n_644) );
AOI322xp5_ASAP7_75t_L g598 ( .A1(n_533), .A2(n_567), .A3(n_574), .B1(n_599), .B2(n_602), .C1(n_603), .C2(n_605), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_533), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g664 ( .A(n_536), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
INVx2_ASAP7_75t_L g541 ( .A(n_538), .Y(n_541) );
INVx1_ASAP7_75t_L g600 ( .A(n_538), .Y(n_600) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_539), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g636 ( .A(n_541), .B(n_549), .Y(n_636) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g548 ( .A(n_543), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g591 ( .A(n_543), .B(n_584), .Y(n_591) );
AND2x2_ASAP7_75t_L g595 ( .A(n_543), .B(n_555), .Y(n_595) );
OAI21xp33_ASAP7_75t_SL g605 ( .A1(n_544), .A2(n_606), .B(n_608), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_544), .A2(n_676), .B1(n_677), .B2(n_679), .Y(n_675) );
INVx3_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g550 ( .A(n_545), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_545), .B(n_565), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_547), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g687 ( .A(n_554), .Y(n_687) );
INVx4_ASAP7_75t_L g560 ( .A(n_555), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_555), .B(n_582), .Y(n_630) );
INVx1_ASAP7_75t_SL g642 ( .A(n_556), .Y(n_642) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g655 ( .A(n_560), .B(n_656), .Y(n_655) );
OAI211xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_563), .B(n_568), .C(n_585), .Y(n_561) );
OAI221xp5_ASAP7_75t_SL g681 ( .A1(n_563), .A2(n_601), .B1(n_680), .B2(n_682), .C(n_684), .Y(n_681) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_565), .B(n_678), .Y(n_677) );
OAI31xp33_ASAP7_75t_L g657 ( .A1(n_566), .A2(n_643), .A3(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g597 ( .A(n_567), .Y(n_597) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g647 ( .A(n_572), .Y(n_647) );
AND2x2_ASAP7_75t_L g660 ( .A(n_574), .B(n_583), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_580), .Y(n_576) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_584), .B(n_687), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B(n_591), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI221xp5_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B1(n_596), .B2(n_597), .C(n_598), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_593), .A2(n_662), .B(n_664), .C(n_667), .Y(n_661) );
CKINVDCx16_ASAP7_75t_R g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_596), .B(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g623 ( .A(n_604), .Y(n_623) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g609 ( .A(n_607), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g651 ( .A(n_607), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI211xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B(n_617), .C(n_626), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_615), .A2(n_625), .B1(n_689), .B2(n_690), .C(n_692), .Y(n_688) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B1(n_621), .B2(n_624), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_628), .B(n_629), .Y(n_626) );
INVx1_ASAP7_75t_SL g689 ( .A(n_628), .Y(n_689) );
INVxp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR4xp25_ASAP7_75t_L g631 ( .A(n_632), .B(n_661), .C(n_681), .D(n_688), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .B(n_639), .C(n_657), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_645), .C(n_649), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g668 ( .A(n_646), .Y(n_668) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
OR2x2_ASAP7_75t_L g679 ( .A(n_647), .B(n_680), .Y(n_679) );
OAI21xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B(n_654), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_673), .C(n_675), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_678), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2x2_ASAP7_75t_L g703 ( .A(n_697), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_711), .Y(n_706) );
NOR2xp33_ASAP7_75t_SL g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_SL g728 ( .A(n_708), .Y(n_728) );
INVx1_ASAP7_75t_L g727 ( .A(n_710), .Y(n_727) );
OA21x2_ASAP7_75t_L g730 ( .A1(n_710), .A2(n_728), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_713), .Y(n_720) );
BUFx2_ASAP7_75t_L g731 ( .A(n_713), .Y(n_731) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B(n_721), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_720), .B(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
endmodule