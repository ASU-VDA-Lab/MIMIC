module fake_jpeg_671_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_22),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_68),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_49),
.Y(n_110)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx12_ASAP7_75t_R g111 ( 
.A(n_63),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_SL g64 ( 
.A1(n_30),
.A2(n_1),
.B(n_3),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_28),
.C(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_4),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_12),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_75),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_12),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_80),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_83),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_20),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_88),
.Y(n_131)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_4),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_86),
.B(n_5),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_32),
.B1(n_23),
.B2(n_21),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_118),
.Y(n_146)
);

OR2x2_ASAP7_75t_SL g162 ( 
.A(n_97),
.B(n_133),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_31),
.B1(n_23),
.B2(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_98),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_31),
.B(n_40),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_100),
.B(n_103),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_18),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_57),
.A2(n_45),
.B1(n_42),
.B2(n_38),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_136),
.B1(n_91),
.B2(n_125),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_54),
.A2(n_28),
.B1(n_38),
.B2(n_35),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_115),
.A2(n_122),
.B1(n_93),
.B2(n_91),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_75),
.B(n_19),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_56),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_58),
.A2(n_35),
.B1(n_40),
.B2(n_33),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_37),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_62),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_128),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_55),
.B(n_26),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_33),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_70),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_88),
.A2(n_80),
.B1(n_74),
.B2(n_87),
.Y(n_136)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_37),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_143),
.B(n_144),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_5),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_145),
.B(n_154),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_125),
.B1(n_127),
.B2(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_71),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_150),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_6),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_152),
.A2(n_160),
.B1(n_113),
.B2(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_130),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_172),
.B1(n_101),
.B2(n_113),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_159),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_103),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_8),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_89),
.A2(n_9),
.B1(n_63),
.B2(n_115),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_9),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_110),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_168),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_114),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_92),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_114),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_89),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_174),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_104),
.A2(n_136),
.B1(n_121),
.B2(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_92),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_96),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_146),
.A2(n_107),
.B1(n_108),
.B2(n_96),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_196),
.B1(n_150),
.B2(n_178),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_147),
.B(n_150),
.Y(n_213)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_137),
.B1(n_138),
.B2(n_99),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_192),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_111),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_200),
.C(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_101),
.B1(n_108),
.B2(n_146),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_152),
.B1(n_170),
.B2(n_168),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_166),
.C(n_141),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_162),
.B(n_159),
.C(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_140),
.B(n_142),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_204),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_174),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_223),
.B(n_190),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_221),
.B1(n_225),
.B2(n_199),
.Y(n_249)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_218),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_156),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_150),
.B1(n_175),
.B2(n_177),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_224),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_149),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_179),
.B1(n_165),
.B2(n_139),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_164),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_231),
.C(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_186),
.B(n_188),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_186),
.B(n_188),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_183),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_233),
.Y(n_252)
);

CKINVDCx11_ASAP7_75t_R g233 ( 
.A(n_193),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_195),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_185),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_235),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_241),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_194),
.C(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_215),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_196),
.B1(n_202),
.B2(n_189),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_245),
.B(n_240),
.Y(n_263)
);

NAND2x1_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_190),
.Y(n_246)
);

A2O1A1O1Ixp25_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_219),
.B(n_218),
.C(n_225),
.D(n_216),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_221),
.B1(n_219),
.B2(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_193),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_247),
.Y(n_261)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_255),
.Y(n_272)
);

XNOR2x2_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_251),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_252),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_259),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_211),
.Y(n_259)
);

OA21x2_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_212),
.B(n_213),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_244),
.B(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_264),
.B(n_266),
.Y(n_276)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_267),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_220),
.B1(n_207),
.B2(n_210),
.Y(n_266)
);

AOI221xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_201),
.B1(n_210),
.B2(n_207),
.C(n_203),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_269),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_262),
.C(n_241),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_277),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_239),
.Y(n_277)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_246),
.B(n_249),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g288 ( 
.A1(n_280),
.A2(n_256),
.B(n_266),
.C(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_268),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_260),
.B(n_254),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_283),
.A2(n_288),
.B(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_250),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_270),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_242),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_268),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_245),
.B(n_242),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_274),
.C(n_275),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_261),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_269),
.B1(n_265),
.B2(n_236),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_272),
.B1(n_290),
.B2(n_253),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_295),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_276),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_280),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_288),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_253),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_297),
.B(n_295),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_308),
.B(n_303),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_296),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_309),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_305),
.B(n_238),
.Y(n_310)
);

OAI221xp5_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_288),
.B1(n_238),
.B2(n_203),
.C(n_201),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_313),
.B(n_311),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);


endmodule