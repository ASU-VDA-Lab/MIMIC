module real_jpeg_16348_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_0),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_36),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_36),
.B1(n_149),
.B2(n_153),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_3),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_3),
.A2(n_46),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_3),
.A2(n_46),
.B1(n_136),
.B2(n_139),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_46),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_5),
.Y(n_249)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_7),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_226),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_225),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_178),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_14),
.B(n_178),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_122),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_47),
.B1(n_120),
.B2(n_121),
.Y(n_15)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_16),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_26),
.B1(n_34),
.B2(n_43),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_25),
.B(n_26),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_19),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_20),
.Y(n_161)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_26),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_26)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_28),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_28),
.Y(n_211)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_30),
.Y(n_165)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_36),
.B1(n_73),
.B2(n_77),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_35),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_35),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_35),
.B(n_251),
.C(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_35),
.B(n_176),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_35),
.B(n_235),
.Y(n_268)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_36),
.B(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_80),
.B1(n_81),
.B2(n_119),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_71),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_58),
.Y(n_49)
);

NAND2x1_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_59),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_50),
.A2(n_58),
.B1(n_72),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_50),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_55),
.Y(n_253)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_58),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

AO22x2_ASAP7_75t_L g233 ( 
.A1(n_71),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_233)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_80),
.A2(n_81),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_R g281 ( 
.A(n_80),
.B(n_233),
.C(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_105),
.B1(n_111),
.B2(n_112),
.Y(n_81)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_96),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B1(n_91),
.B2(n_94),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_111),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_156),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_130),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_124),
.A2(n_181),
.B1(n_182),
.B2(n_185),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_130),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_130),
.B(n_261),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B(n_141),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_142),
.B1(n_148),
.B2(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_138),
.Y(n_257)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_148),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_172),
.B2(n_173),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_167),
.B2(n_171),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_172),
.A2(n_173),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_173),
.B(n_186),
.C(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_173),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_173),
.B(n_268),
.Y(n_269)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_186),
.C(n_192),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_179),
.A2(n_180),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_184),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_184),
.B(n_245),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_186),
.A2(n_239),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_186),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_186),
.A2(n_192),
.B1(n_276),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_220),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_220),
.Y(n_237)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_196),
.A3(n_199),
.B1(n_205),
.B2(n_212),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_280),
.B(n_286),
.Y(n_227)
);

OAI21x1_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_242),
.B(n_279),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_230),
.B(n_238),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_233),
.B1(n_246),
.B2(n_258),
.Y(n_245)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_233),
.B(n_258),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

AOI21x1_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_271),
.B(n_278),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_259),
.B(n_270),
.Y(n_243)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_267),
.B(n_269),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_272),
.B(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);


endmodule