module real_aes_9421_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_874, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_874;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g191 ( .A(n_0), .B(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g525 ( .A(n_1), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_2), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_3), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_4), .B(n_506), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_5), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_6), .B(n_198), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_7), .Y(n_184) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_8), .B(n_87), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_9), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_10), .B(n_171), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_11), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_12), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_13), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_14), .B(n_187), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_15), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_16), .B(n_174), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_17), .B(n_216), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_18), .B(n_187), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_19), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_20), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_21), .B(n_198), .Y(n_231) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_22), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_23), .B(n_171), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_24), .B(n_153), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_25), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_26), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_27), .B(n_153), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_28), .B(n_216), .Y(n_580) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_29), .Y(n_145) );
OAI21xp33_ASAP7_75t_L g503 ( .A1(n_30), .A2(n_190), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_31), .B(n_171), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_32), .B(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_33), .B(n_169), .Y(n_168) );
NAND2xp33_ASAP7_75t_SL g151 ( .A(n_34), .B(n_147), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_35), .B(n_171), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_36), .B(n_235), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_37), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_38), .B(n_144), .Y(n_278) );
INVx1_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
OAI21x1_ASAP7_75t_L g138 ( .A1(n_40), .A2(n_70), .B(n_139), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_41), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_42), .B(n_171), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_43), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_44), .B(n_235), .Y(n_234) );
AND2x6_ASAP7_75t_L g158 ( .A(n_45), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_46), .B(n_135), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_47), .A2(n_83), .B1(n_506), .B2(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_48), .B(n_135), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_49), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_50), .B(n_165), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_51), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_52), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_53), .Y(n_543) );
INVx1_ASAP7_75t_L g159 ( .A(n_54), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_55), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_56), .B(n_221), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_57), .A2(n_123), .B1(n_124), .B2(n_486), .Y(n_122) );
INVxp33_ASAP7_75t_SL g486 ( .A(n_57), .Y(n_486) );
XOR2x1_ASAP7_75t_L g489 ( .A(n_57), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_58), .B(n_507), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_59), .B(n_507), .Y(n_565) );
NAND2xp33_ASAP7_75t_L g146 ( .A(n_60), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_61), .B(n_235), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_62), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_63), .B(n_165), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_64), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g101 ( .A(n_65), .B(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g535 ( .A(n_66), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_67), .B(n_153), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_68), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_69), .B(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_71), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_72), .B(n_187), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_73), .B(n_216), .Y(n_229) );
INVx1_ASAP7_75t_L g529 ( .A(n_74), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_75), .B(n_235), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_76), .Y(n_600) );
BUFx10_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
INVx1_ASAP7_75t_L g594 ( .A(n_78), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_79), .B(n_187), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_80), .B(n_171), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_81), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_82), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_84), .B(n_165), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_85), .B(n_187), .Y(n_228) );
INVx1_ASAP7_75t_L g538 ( .A(n_86), .Y(n_538) );
INVx2_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
OR2x2_ASAP7_75t_L g105 ( .A(n_89), .B(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_L g120 ( .A(n_89), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_89), .B(n_107), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_90), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_91), .B(n_169), .Y(n_276) );
INVx1_ASAP7_75t_L g102 ( .A(n_92), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_93), .B(n_198), .Y(n_206) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_94), .B(n_501), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_95), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_96), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_96), .B(n_868), .Y(n_867) );
NAND2xp33_ASAP7_75t_L g604 ( .A(n_97), .B(n_165), .Y(n_604) );
AOI21xp5_ASAP7_75t_SL g98 ( .A1(n_99), .A2(n_110), .B(n_861), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_103), .Y(n_100) );
INVx4_ASAP7_75t_L g866 ( .A(n_101), .Y(n_866) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx4_ASAP7_75t_L g847 ( .A(n_104), .Y(n_847) );
INVx5_ASAP7_75t_L g851 ( .A(n_104), .Y(n_851) );
OR2x2_ASAP7_75t_SL g863 ( .A(n_104), .B(n_864), .Y(n_863) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g872 ( .A(n_105), .Y(n_872) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x6_ASAP7_75t_L g113 ( .A(n_107), .B(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
OAI221xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_116), .B1(n_843), .B2(n_852), .C(n_855), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g859 ( .A(n_114), .B(n_860), .Y(n_859) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx12f_ASAP7_75t_L g854 ( .A(n_115), .Y(n_854) );
NOR2x1p5_ASAP7_75t_L g865 ( .A(n_115), .B(n_866), .Y(n_865) );
AOI21x1_ASAP7_75t_L g871 ( .A1(n_115), .A2(n_866), .B(n_872), .Y(n_871) );
AOI21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_487), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVxp67_ASAP7_75t_L g488 ( .A(n_119), .Y(n_488) );
BUFx8_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g844 ( .A(n_124), .B(n_845), .Y(n_844) );
NAND2x1p5_ASAP7_75t_L g124 ( .A(n_125), .B(n_407), .Y(n_124) );
NOR2x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_331), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_301), .Y(n_126) );
AOI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_209), .B1(n_237), .B2(n_268), .C(n_281), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_161), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g360 ( .A(n_131), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_131), .B(n_359), .Y(n_425) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g309 ( .A(n_132), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g382 ( .A(n_132), .B(n_248), .Y(n_382) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g284 ( .A(n_133), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_133), .B(n_248), .Y(n_346) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_133), .Y(n_387) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g269 ( .A(n_134), .B(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_134), .Y(n_354) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_140), .B(n_160), .Y(n_134) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_135), .A2(n_226), .B(n_234), .Y(n_225) );
INVx2_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g208 ( .A(n_136), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_136), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx5_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g193 ( .A(n_138), .Y(n_193) );
OAI21x1_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_150), .B(n_156), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_146), .C(n_148), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_143), .A2(n_544), .B1(n_550), .B2(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g174 ( .A(n_144), .Y(n_174) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_144), .A2(n_171), .B1(n_183), .B2(n_184), .Y(n_182) );
INVx2_ASAP7_75t_L g506 ( .A(n_144), .Y(n_506) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_145), .Y(n_147) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_145), .Y(n_154) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx1_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
INVx2_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
INVx2_ASAP7_75t_L g502 ( .A(n_147), .Y(n_502) );
INVx2_ASAP7_75t_L g504 ( .A(n_147), .Y(n_504) );
INVx2_ASAP7_75t_L g507 ( .A(n_147), .Y(n_507) );
INVx2_ASAP7_75t_SL g155 ( .A(n_148), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_148), .A2(n_168), .B(n_170), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_148), .A2(n_215), .B(n_217), .Y(n_214) );
INVx2_ASAP7_75t_SL g233 ( .A(n_148), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_148), .A2(n_514), .B(n_515), .Y(n_513) );
CKINVDCx6p67_ASAP7_75t_R g566 ( .A(n_148), .Y(n_566) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx12f_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
INVx5_ASAP7_75t_L g202 ( .A(n_149), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_155), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_153), .B(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_153), .B(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_L g611 ( .A(n_153), .Y(n_611) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
INVx2_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
INVx2_ASAP7_75t_L g254 ( .A(n_154), .Y(n_254) );
INVx2_ASAP7_75t_L g544 ( .A(n_154), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_155), .A2(n_173), .B(n_175), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_155), .A2(n_158), .B(n_182), .C(n_185), .Y(n_181) );
AOI21x1_ASAP7_75t_L g218 ( .A1(n_155), .A2(n_219), .B(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_155), .A2(n_517), .B(n_518), .Y(n_516) );
OAI21x1_ASAP7_75t_L g213 ( .A1(n_156), .A2(n_214), .B(n_218), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_156), .A2(n_252), .B(n_256), .Y(n_251) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_156), .A2(n_513), .B(n_516), .Y(n_512) );
INVx2_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
INVx8_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g601 ( .A1(n_157), .A2(n_235), .B(n_602), .Y(n_601) );
INVx8_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OAI21x1_ASAP7_75t_SL g195 ( .A1(n_158), .A2(n_196), .B(n_203), .Y(n_195) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_158), .A2(n_227), .B(n_230), .Y(n_226) );
AOI21xp33_ASAP7_75t_L g539 ( .A1(n_158), .A2(n_236), .B(n_537), .Y(n_539) );
INVx1_ASAP7_75t_L g547 ( .A(n_158), .Y(n_547) );
INVx1_ASAP7_75t_L g614 ( .A(n_158), .Y(n_614) );
INVx1_ASAP7_75t_SL g484 ( .A(n_161), .Y(n_484) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_179), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_162), .B(n_329), .Y(n_363) );
BUFx2_ASAP7_75t_L g385 ( .A(n_162), .Y(n_385) );
AND2x2_ASAP7_75t_L g400 ( .A(n_162), .B(n_243), .Y(n_400) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx3_ASAP7_75t_L g294 ( .A(n_163), .Y(n_294) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g248 ( .A(n_164), .Y(n_248) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_177), .Y(n_164) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_165), .A2(n_181), .B(n_191), .Y(n_180) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_165), .A2(n_251), .B(n_260), .Y(n_250) );
OAI21x1_ASAP7_75t_L g272 ( .A1(n_165), .A2(n_273), .B(n_280), .Y(n_272) );
INVx2_ASAP7_75t_L g498 ( .A(n_165), .Y(n_498) );
NOR2x1p5_ASAP7_75t_SL g613 ( .A(n_165), .B(n_614), .Y(n_613) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_172), .B(n_176), .Y(n_166) );
INVx2_ASAP7_75t_L g527 ( .A(n_171), .Y(n_527) );
INVx2_ASAP7_75t_L g577 ( .A(n_171), .Y(n_577) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_176), .A2(n_274), .B(n_277), .Y(n_273) );
AO31x2_ASAP7_75t_L g497 ( .A1(n_176), .A2(n_498), .A3(n_499), .B(n_508), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_176), .A2(n_563), .B(n_567), .Y(n_562) );
OAI21x1_ASAP7_75t_SL g573 ( .A1(n_176), .A2(n_574), .B(n_579), .Y(n_573) );
AND2x2_ASAP7_75t_L g405 ( .A(n_179), .B(n_211), .Y(n_405) );
AND2x2_ASAP7_75t_L g481 ( .A(n_179), .B(n_307), .Y(n_481) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_194), .Y(n_179) );
INVx3_ASAP7_75t_L g243 ( .A(n_180), .Y(n_243) );
INVx2_ASAP7_75t_L g305 ( .A(n_180), .Y(n_305) );
AND2x2_ASAP7_75t_L g320 ( .A(n_180), .B(n_266), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_188), .B(n_190), .Y(n_185) );
INVx5_ASAP7_75t_L g216 ( .A(n_187), .Y(n_216) );
OR2x2_ASAP7_75t_L g596 ( .A(n_187), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g258 ( .A(n_189), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_190), .A2(n_204), .B(n_206), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_190), .A2(n_500), .B1(n_503), .B2(n_505), .Y(n_499) );
BUFx2_ASAP7_75t_L g530 ( .A(n_190), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_190), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_190), .B(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g578 ( .A(n_190), .Y(n_578) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_192), .A2(n_195), .B(n_207), .Y(n_194) );
BUFx4f_ASAP7_75t_L g222 ( .A(n_192), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_192), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_L g561 ( .A(n_192), .Y(n_561) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g236 ( .A(n_193), .Y(n_236) );
INVx3_ASAP7_75t_L g242 ( .A(n_194), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_200), .C(n_202), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_198), .A2(n_527), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g201 ( .A(n_199), .Y(n_201) );
INVx2_ASAP7_75t_L g221 ( .A(n_201), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_202), .A2(n_228), .B(n_229), .Y(n_227) );
O2A1O1Ixp5_ASAP7_75t_L g256 ( .A1(n_202), .A2(n_257), .B(n_258), .C(n_259), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_202), .A2(n_278), .B(n_279), .Y(n_277) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_202), .A2(n_542), .B(n_546), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_202), .A2(n_568), .B(n_569), .Y(n_567) );
INVx1_ASAP7_75t_L g582 ( .A(n_202), .Y(n_582) );
INVx2_ASAP7_75t_L g533 ( .A(n_205), .Y(n_533) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x6_ASAP7_75t_L g439 ( .A(n_210), .B(n_440), .Y(n_439) );
OAI33xp33_ASAP7_75t_L g482 ( .A1(n_210), .A2(n_305), .A3(n_309), .B1(n_483), .B2(n_484), .B3(n_485), .Y(n_482) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_211), .B(n_376), .Y(n_429) );
INVx1_ASAP7_75t_L g452 ( .A(n_211), .Y(n_452) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_224), .Y(n_211) );
AND2x2_ASAP7_75t_L g239 ( .A(n_212), .B(n_225), .Y(n_239) );
BUFx2_ASAP7_75t_L g375 ( .A(n_212), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_222), .B(n_223), .Y(n_212) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_213), .A2(n_222), .B(n_223), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_216), .A2(n_533), .B1(n_534), .B2(n_535), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_216), .A2(n_506), .B1(n_607), .B2(n_608), .Y(n_606) );
OAI21x1_ASAP7_75t_L g511 ( .A1(n_222), .A2(n_512), .B(n_519), .Y(n_511) );
OAI21x1_ASAP7_75t_SL g572 ( .A1(n_222), .A2(n_573), .B(n_583), .Y(n_572) );
AND2x2_ASAP7_75t_L g262 ( .A(n_224), .B(n_242), .Y(n_262) );
INVx1_ASAP7_75t_L g300 ( .A(n_224), .Y(n_300) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_224), .Y(n_319) );
NOR2xp67_ASAP7_75t_L g356 ( .A(n_224), .B(n_297), .Y(n_356) );
INVx1_ASAP7_75t_L g373 ( .A(n_224), .Y(n_373) );
INVx1_ASAP7_75t_L g402 ( .A(n_224), .Y(n_402) );
AND2x2_ASAP7_75t_L g413 ( .A(n_224), .B(n_366), .Y(n_413) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_233), .A2(n_253), .B(n_255), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_233), .A2(n_275), .B(n_276), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_233), .A2(n_610), .B(n_611), .C(n_612), .Y(n_609) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_236), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_236), .B(n_594), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_244), .B1(n_249), .B2(n_261), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_239), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g336 ( .A(n_239), .Y(n_336) );
AND2x2_ASAP7_75t_L g364 ( .A(n_239), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g390 ( .A(n_239), .B(n_323), .Y(n_390) );
AND2x2_ASAP7_75t_L g427 ( .A(n_239), .B(n_338), .Y(n_427) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_241), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_242), .Y(n_323) );
AND2x2_ASAP7_75t_L g338 ( .A(n_242), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_SL g366 ( .A(n_242), .Y(n_366) );
INVx1_ASAP7_75t_L g376 ( .A(n_242), .Y(n_376) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_242), .Y(n_418) );
AND2x2_ASAP7_75t_L g265 ( .A(n_243), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g339 ( .A(n_243), .Y(n_339) );
AND2x2_ASAP7_75t_L g365 ( .A(n_243), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g349 ( .A(n_245), .B(n_330), .Y(n_349) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g455 ( .A(n_246), .B(n_283), .Y(n_455) );
INVx1_ASAP7_75t_L g468 ( .A(n_246), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
INVx2_ASAP7_75t_L g392 ( .A(n_247), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_247), .B(n_284), .Y(n_437) );
BUFx2_ASAP7_75t_L g462 ( .A(n_247), .Y(n_462) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g359 ( .A(n_249), .Y(n_359) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g288 ( .A(n_250), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x4_ASAP7_75t_L g306 ( .A(n_262), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g313 ( .A(n_262), .Y(n_313) );
AND2x2_ASAP7_75t_L g454 ( .A(n_262), .B(n_419), .Y(n_454) );
AND2x2_ASAP7_75t_L g476 ( .A(n_262), .B(n_304), .Y(n_476) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x6_ASAP7_75t_L g458 ( .A(n_264), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g355 ( .A(n_265), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g449 ( .A(n_265), .B(n_413), .Y(n_449) );
AND2x4_ASAP7_75t_L g299 ( .A(n_266), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_SL g307 ( .A(n_266), .Y(n_307) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_R g419 ( .A(n_267), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_268), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g479 ( .A(n_268), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_269), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_269), .B(n_327), .Y(n_396) );
AOI322xp5_ASAP7_75t_L g397 ( .A1(n_269), .A2(n_351), .A3(n_398), .B1(n_401), .B2(n_403), .C1(n_405), .C2(n_406), .Y(n_397) );
INVx1_ASAP7_75t_L g310 ( .A(n_270), .Y(n_310) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g289 ( .A(n_271), .Y(n_289) );
AND2x2_ASAP7_75t_L g316 ( .A(n_271), .B(n_287), .Y(n_316) );
INVx1_ASAP7_75t_L g353 ( .A(n_271), .Y(n_353) );
AND2x2_ASAP7_75t_L g370 ( .A(n_271), .B(n_288), .Y(n_370) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI21xp33_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_290), .B(n_295), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_282), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
OR2x2_ASAP7_75t_L g362 ( .A(n_283), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g448 ( .A(n_283), .B(n_370), .Y(n_448) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g335 ( .A(n_284), .B(n_310), .Y(n_335) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g291 ( .A(n_286), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g441 ( .A(n_286), .B(n_385), .Y(n_441) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g325 ( .A(n_287), .Y(n_325) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g329 ( .A(n_288), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_289), .Y(n_330) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g314 ( .A(n_293), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g334 ( .A(n_293), .B(n_335), .Y(n_334) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_293), .B(n_369), .Y(n_368) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_293), .B(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g327 ( .A(n_294), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g406 ( .A(n_294), .B(n_359), .Y(n_406) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
OR2x2_ASAP7_75t_L g432 ( .A(n_296), .B(n_318), .Y(n_432) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g483 ( .A(n_299), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_308), .B(n_311), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g312 ( .A(n_304), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g451 ( .A(n_304), .B(n_452), .Y(n_451) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_305), .B(n_373), .Y(n_404) );
INVx2_ASAP7_75t_L g395 ( .A(n_307), .Y(n_395) );
BUFx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g434 ( .A(n_309), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_309), .B(n_462), .Y(n_461) );
NAND2xp67_ASAP7_75t_SL g485 ( .A(n_309), .B(n_392), .Y(n_485) );
OAI222xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_314), .B2(n_317), .C1(n_324), .C2(n_326), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_314), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g426 ( .A(n_315), .Y(n_426) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g386 ( .A(n_316), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
BUFx3_ASAP7_75t_L g341 ( .A(n_318), .Y(n_341) );
NAND2x1_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g412 ( .A(n_320), .B(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
NAND2x1_ASAP7_75t_L g326 ( .A(n_327), .B(n_330), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_327), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g472 ( .A(n_327), .B(n_421), .Y(n_472) );
INVx1_ASAP7_75t_L g478 ( .A(n_327), .Y(n_478) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_357), .C(n_377), .Y(n_331) );
AOI322xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_336), .A3(n_337), .B1(n_340), .B2(n_342), .C1(n_347), .C2(n_355), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_334), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g421 ( .A(n_335), .Y(n_421) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_335), .Y(n_435) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g447 ( .A(n_338), .B(n_399), .Y(n_447) );
AND2x2_ASAP7_75t_L g372 ( .A(n_339), .B(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_341), .A2(n_458), .B1(n_461), .B2(n_463), .Y(n_460) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AOI222xp33_ASAP7_75t_L g409 ( .A1(n_349), .A2(n_410), .B1(n_412), .B2(n_414), .C1(n_416), .C2(n_420), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_351), .B(n_392), .Y(n_415) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g391 ( .A(n_352), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_355), .A2(n_358), .B1(n_361), .B2(n_364), .C(n_367), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g446 ( .A(n_360), .B(n_370), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_363), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g480 ( .A(n_363), .Y(n_480) );
INVx2_ASAP7_75t_L g440 ( .A(n_365), .Y(n_440) );
AND2x2_ASAP7_75t_L g465 ( .A(n_365), .B(n_419), .Y(n_465) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_371), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g381 ( .A(n_370), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g473 ( .A(n_370), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_372), .Y(n_378) );
AND2x4_ASAP7_75t_L g416 ( .A(n_372), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx2_ASAP7_75t_L g399 ( .A(n_375), .Y(n_399) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_375), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_388), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx2_ASAP7_75t_L g443 ( .A(n_386), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B1(n_393), .B2(n_396), .C(n_397), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_392), .A2(n_457), .B(n_460), .Y(n_456) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_402), .B(n_418), .Y(n_459) );
INVx1_ASAP7_75t_L g411 ( .A(n_405), .Y(n_411) );
INVxp67_ASAP7_75t_L g463 ( .A(n_406), .Y(n_463) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_408), .B(n_444), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_422), .C(n_430), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_421), .B(n_468), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_426), .B(n_427), .C(n_428), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_429), .B(n_443), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B1(n_438), .B2(n_441), .C(n_442), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .C(n_436), .Y(n_433) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g471 ( .A(n_440), .Y(n_471) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_445), .B(n_456), .C(n_464), .D(n_475), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B1(n_448), .B2(n_449), .C(n_450), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B(n_455), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_469), .B2(n_472), .C1(n_473), .C2(n_874), .Y(n_464) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_479), .B2(n_481), .C(n_482), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2x1p5_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
NOR2x1p5_ASAP7_75t_L g490 ( .A(n_491), .B(n_766), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_719), .Y(n_491) );
NOR4xp25_ASAP7_75t_L g492 ( .A(n_493), .B(n_630), .C(n_661), .D(n_695), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_553), .B(n_621), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AOI322xp5_ASAP7_75t_L g733 ( .A1(n_495), .A2(n_622), .A3(n_644), .B1(n_734), .B2(n_735), .C1(n_736), .C2(n_737), .Y(n_733) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_520), .Y(n_495) );
INVx1_ASAP7_75t_L g678 ( .A(n_496), .Y(n_678) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_510), .Y(n_496) );
INVx2_ASAP7_75t_L g626 ( .A(n_497), .Y(n_626) );
INVx2_ASAP7_75t_SL g642 ( .A(n_497), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_497), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g671 ( .A(n_497), .B(n_627), .Y(n_671) );
INVx1_ASAP7_75t_L g687 ( .A(n_497), .Y(n_687) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_506), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
AND2x2_ASAP7_75t_L g645 ( .A(n_510), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g690 ( .A(n_510), .Y(n_690) );
AND2x2_ASAP7_75t_L g706 ( .A(n_510), .B(n_674), .Y(n_706) );
AND2x2_ASAP7_75t_L g718 ( .A(n_510), .B(n_540), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_510), .B(n_660), .Y(n_773) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_510), .Y(n_823) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx3_ASAP7_75t_L g627 ( .A(n_511), .Y(n_627) );
BUFx3_ASAP7_75t_L g806 ( .A(n_520), .Y(n_806) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_540), .Y(n_520) );
OR2x2_ASAP7_75t_L g629 ( .A(n_521), .B(n_540), .Y(n_629) );
INVx2_ASAP7_75t_L g640 ( .A(n_521), .Y(n_640) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g646 ( .A(n_522), .Y(n_646) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_531), .B(n_539), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_528), .B(n_530), .Y(n_523) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_536), .B(n_537), .Y(n_531) );
AO21x1_ASAP7_75t_L g589 ( .A1(n_536), .A2(n_590), .B(n_593), .Y(n_589) );
AOI21x1_ASAP7_75t_L g595 ( .A1(n_536), .A2(n_596), .B(n_598), .Y(n_595) );
AND2x4_ASAP7_75t_L g641 ( .A(n_540), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g648 ( .A(n_540), .Y(n_648) );
INVx2_ASAP7_75t_SL g674 ( .A(n_540), .Y(n_674) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_540), .Y(n_677) );
AND2x2_ASAP7_75t_L g794 ( .A(n_540), .B(n_640), .Y(n_794) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_548), .B(n_552), .Y(n_540) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_615), .Y(n_553) );
NOR2xp67_ASAP7_75t_L g554 ( .A(n_555), .B(n_584), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_555), .B(n_686), .C(n_688), .Y(n_685) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g817 ( .A(n_556), .B(n_783), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_556), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_571), .Y(n_557) );
INVx2_ASAP7_75t_L g655 ( .A(n_558), .Y(n_655) );
AND2x2_ASAP7_75t_L g712 ( .A(n_558), .B(n_618), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_558), .B(n_603), .Y(n_759) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g634 ( .A(n_559), .Y(n_634) );
OAI21x1_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_562), .B(n_570), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B(n_566), .Y(n_563) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_566), .A2(n_606), .B(n_609), .C(n_613), .Y(n_605) );
AND2x4_ASAP7_75t_L g700 ( .A(n_571), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g710 ( .A(n_571), .B(n_603), .Y(n_710) );
INVx1_ASAP7_75t_L g765 ( .A(n_571), .Y(n_765) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g618 ( .A(n_572), .Y(n_618) );
AOI21x1_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_578), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B(n_582), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_584), .A2(n_833), .B1(n_835), .B2(n_836), .C(n_838), .Y(n_832) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g824 ( .A(n_585), .B(n_653), .Y(n_824) );
AND2x2_ASAP7_75t_L g840 ( .A(n_585), .B(n_712), .Y(n_840) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_603), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_586), .B(n_620), .Y(n_623) );
INVx2_ASAP7_75t_L g732 ( .A(n_586), .Y(n_732) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_587), .Y(n_715) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g617 ( .A(n_588), .Y(n_617) );
BUFx3_ASAP7_75t_L g652 ( .A(n_588), .Y(n_652) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_595), .B(n_601), .Y(n_588) );
INVxp67_ASAP7_75t_L g602 ( .A(n_593), .Y(n_602) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g620 ( .A(n_603), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_603), .B(n_617), .Y(n_657) );
INVx1_ASAP7_75t_L g665 ( .A(n_603), .Y(n_665) );
INVx1_ASAP7_75t_L g701 ( .A(n_603), .Y(n_701) );
HB1xp67_ASAP7_75t_SL g725 ( .A(n_603), .Y(n_725) );
INVx1_ASAP7_75t_L g763 ( .A(n_603), .Y(n_763) );
AND2x4_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_615), .A2(n_622), .B(n_624), .Y(n_621) );
AND2x4_ASAP7_75t_SL g615 ( .A(n_616), .B(n_619), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g664 ( .A(n_617), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g743 ( .A(n_617), .Y(n_743) );
INVx2_ASAP7_75t_L g635 ( .A(n_618), .Y(n_635) );
AND2x4_ASAP7_75t_L g653 ( .A(n_618), .B(n_633), .Y(n_653) );
BUFx2_ASAP7_75t_L g667 ( .A(n_618), .Y(n_667) );
AND2x2_ASAP7_75t_L g730 ( .A(n_618), .B(n_620), .Y(n_730) );
INVx1_ASAP7_75t_L g736 ( .A(n_619), .Y(n_736) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g681 ( .A(n_620), .B(n_633), .Y(n_681) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g791 ( .A(n_623), .B(n_792), .Y(n_791) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_628), .Y(n_624) );
AND2x4_ASAP7_75t_SL g658 ( .A(n_625), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_625), .B(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_SL g727 ( .A(n_625), .B(n_673), .Y(n_727) );
AOI32xp33_ASAP7_75t_L g776 ( .A1(n_625), .A2(n_638), .A3(n_754), .B1(n_777), .B2(n_778), .Y(n_776) );
INVxp67_ASAP7_75t_L g807 ( .A(n_625), .Y(n_807) );
AND2x4_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x4_ASAP7_75t_L g717 ( .A(n_626), .B(n_640), .Y(n_717) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_627), .Y(n_637) );
AND2x4_ASAP7_75t_L g745 ( .A(n_628), .B(n_671), .Y(n_745) );
AND2x4_ASAP7_75t_L g748 ( .A(n_628), .B(n_637), .Y(n_748) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g811 ( .A(n_629), .B(n_650), .Y(n_811) );
OAI21xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_636), .B(n_643), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_631), .B(n_731), .Y(n_818) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI31xp33_ASAP7_75t_L g711 ( .A1(n_632), .A2(n_712), .A3(n_713), .B(n_716), .Y(n_711) );
OR4x1_ASAP7_75t_L g772 ( .A(n_632), .B(n_773), .C(n_774), .D(n_775), .Y(n_772) );
AND2x2_ASAP7_75t_L g777 ( .A(n_632), .B(n_731), .Y(n_777) );
AND2x4_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g709 ( .A(n_633), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_633), .B(n_715), .Y(n_714) );
BUFx2_ASAP7_75t_L g792 ( .A(n_633), .Y(n_792) );
INVx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x4_ASAP7_75t_L g668 ( .A(n_634), .B(n_652), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
OR2x2_ASAP7_75t_L g750 ( .A(n_637), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g801 ( .A(n_637), .Y(n_801) );
AND2x2_ASAP7_75t_L g839 ( .A(n_637), .B(n_673), .Y(n_839) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g694 ( .A(n_639), .Y(n_694) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g734 ( .A(n_641), .B(n_645), .Y(n_734) );
INVx2_ASAP7_75t_L g751 ( .A(n_641), .Y(n_751) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_641), .Y(n_760) );
AND2x2_ASAP7_75t_L g837 ( .A(n_641), .B(n_694), .Y(n_837) );
INVx1_ASAP7_75t_L g705 ( .A(n_642), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_649), .B1(n_654), .B2(n_658), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx2_ASAP7_75t_L g660 ( .A(n_646), .Y(n_660) );
AND2x2_ASAP7_75t_L g673 ( .A(n_646), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g684 ( .A(n_646), .B(n_651), .Y(n_684) );
INVx1_ASAP7_75t_L g774 ( .A(n_647), .Y(n_774) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
AND2x2_ASAP7_75t_L g754 ( .A(n_650), .B(n_700), .Y(n_754) );
AND2x2_ASAP7_75t_L g771 ( .A(n_650), .B(n_730), .Y(n_771) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_653), .A2(n_683), .B1(n_685), .B2(n_691), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_653), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_SL g735 ( .A(n_653), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_653), .B(n_692), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_654), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AND2x4_ASAP7_75t_L g663 ( .A(n_655), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g702 ( .A(n_655), .Y(n_702) );
AND2x2_ASAP7_75t_L g784 ( .A(n_655), .B(n_710), .Y(n_784) );
INVx1_ASAP7_75t_L g809 ( .A(n_655), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_656), .B(n_712), .Y(n_797) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g804 ( .A(n_657), .Y(n_804) );
INVx1_ASAP7_75t_L g778 ( .A(n_659), .Y(n_778) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_660), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g780 ( .A(n_660), .B(n_705), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_669), .B1(n_675), .B2(n_679), .C(n_682), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx2_ASAP7_75t_L g692 ( .A(n_664), .Y(n_692) );
AOI322xp5_ASAP7_75t_L g813 ( .A1(n_666), .A2(n_670), .A3(n_722), .B1(n_814), .B2(n_816), .C1(n_817), .C2(n_818), .Y(n_813) );
AND2x4_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AND2x4_ASAP7_75t_L g680 ( .A(n_667), .B(n_681), .Y(n_680) );
OR2x6_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g723 ( .A(n_671), .B(n_676), .Y(n_723) );
AND2x2_ASAP7_75t_L g793 ( .A(n_671), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_671), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g830 ( .A(n_671), .Y(n_830) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g800 ( .A(n_673), .B(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g770 ( .A(n_675), .Y(n_770) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g697 ( .A(n_677), .Y(n_697) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI31xp33_ASAP7_75t_L g795 ( .A1(n_680), .A2(n_796), .A3(n_798), .B(n_800), .Y(n_795) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_681), .Y(n_737) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g693 ( .A(n_686), .Y(n_693) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g722 ( .A(n_689), .B(n_717), .Y(n_722) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .C(n_694), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_703), .B2(n_707), .C(n_711), .Y(n_695) );
INVx1_ASAP7_75t_L g755 ( .A(n_696), .Y(n_755) );
OR2x2_ASAP7_75t_L g829 ( .A(n_697), .B(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_699), .B(n_732), .Y(n_785) );
AND2x4_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
BUFx2_ASAP7_75t_L g789 ( .A(n_700), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
AND2x2_ASAP7_75t_L g816 ( .A(n_706), .B(n_717), .Y(n_816) );
AND2x4_ASAP7_75t_L g842 ( .A(n_706), .B(n_780), .Y(n_842) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx2_ASAP7_75t_L g744 ( .A(n_710), .Y(n_744) );
BUFx2_ASAP7_75t_L g841 ( .A(n_712), .Y(n_841) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g799 ( .A(n_714), .B(n_744), .Y(n_799) );
INVx1_ASAP7_75t_L g783 ( .A(n_715), .Y(n_783) );
AND2x2_ASAP7_75t_SL g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NOR3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_738), .C(n_752), .Y(n_719) );
OAI221xp5_ASAP7_75t_SL g720 ( .A1(n_721), .A2(n_724), .B1(n_726), .B2(n_728), .C(n_733), .Y(n_720) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_722), .A2(n_757), .B1(n_760), .B2(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OR2x6_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g758 ( .A(n_732), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_735), .B(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_746), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_745), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g775 ( .A(n_742), .Y(n_775) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_743), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g827 ( .A(n_743), .Y(n_827) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g752 ( .A(n_753), .B(n_756), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NAND4xp75_ASAP7_75t_L g766 ( .A(n_767), .B(n_786), .C(n_812), .D(n_831), .Y(n_766) );
NOR2x1_ASAP7_75t_L g767 ( .A(n_768), .B(n_779), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .C(n_776), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g835 ( .A(n_784), .Y(n_835) );
NOR2x1_ASAP7_75t_L g786 ( .A(n_787), .B(n_802), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_795), .Y(n_787) );
OAI21xp33_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B(n_793), .Y(n_788) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g815 ( .A(n_794), .Y(n_815) );
AND2x2_ASAP7_75t_L g834 ( .A(n_794), .B(n_801), .Y(n_834) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_805), .B1(n_807), .B2(n_808), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_806), .B(n_822), .Y(n_821) );
NAND2x1_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_819), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_824), .B1(n_825), .B2(n_828), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_839), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_838) );
OAI21xp33_ASAP7_75t_L g861 ( .A1(n_843), .A2(n_862), .B(n_867), .Y(n_861) );
AOI21xp5_ASAP7_75t_SL g843 ( .A1(n_844), .A2(n_846), .B(n_848), .Y(n_843) );
INVx5_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx6_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_853), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_SL g856 ( .A(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx12f_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
BUFx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx6_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
endmodule