module fake_jpeg_7679_n_303 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_40),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_0),
.C(n_1),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_21),
.B(n_30),
.C(n_19),
.Y(n_44)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_26),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_27),
.B1(n_20),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_63),
.B1(n_25),
.B2(n_18),
.Y(n_82)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_27),
.B1(n_20),
.B2(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_37),
.A2(n_40),
.B1(n_18),
.B2(n_22),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_22),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_79),
.B(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_41),
.B1(n_42),
.B2(n_36),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_90),
.B1(n_55),
.B2(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_42),
.B1(n_43),
.B2(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_84),
.B1(n_52),
.B2(n_51),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_42),
.B1(n_39),
.B2(n_36),
.Y(n_72)
);

AO22x2_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_55),
.B1(n_58),
.B2(n_51),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_43),
.C(n_39),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_94),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_82),
.B1(n_56),
.B2(n_47),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_24),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_26),
.B1(n_22),
.B2(n_25),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_39),
.B1(n_17),
.B2(n_31),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_50),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_46),
.A2(n_19),
.B1(n_31),
.B2(n_17),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_41),
.B1(n_28),
.B2(n_23),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_52),
.B(n_58),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_39),
.B1(n_23),
.B2(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_1),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_66),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_33),
.C(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_95),
.B(n_96),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_106),
.B(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_60),
.B1(n_73),
.B2(n_83),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_91),
.B1(n_84),
.B2(n_24),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_65),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_74),
.B(n_13),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_118),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_61),
.B(n_24),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_48),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_61),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_1),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_56),
.B1(n_60),
.B2(n_33),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_90),
.B1(n_69),
.B2(n_70),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_70),
.B1(n_86),
.B2(n_73),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_131),
.B(n_109),
.C(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_144),
.B1(n_148),
.B2(n_105),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_76),
.C(n_94),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_141),
.C(n_103),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_89),
.B1(n_81),
.B2(n_71),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_130),
.B1(n_140),
.B2(n_147),
.Y(n_164)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_136),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_79),
.B1(n_70),
.B2(n_93),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_119),
.Y(n_152)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_145),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_79),
.B1(n_93),
.B2(n_87),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_79),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_13),
.C(n_16),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_110),
.A2(n_91),
.B1(n_33),
.B2(n_24),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_33),
.B1(n_24),
.B2(n_29),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_102),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_161),
.C(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

XNOR2x2_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_105),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_157),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_159),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_117),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_154),
.B1(n_173),
.B2(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_121),
.B1(n_114),
.B2(n_103),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_85),
.B1(n_11),
.B2(n_12),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_128),
.B1(n_139),
.B2(n_140),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_129),
.A2(n_104),
.B(n_99),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_138),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_169),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_134),
.A2(n_129),
.B(n_143),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_172),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_108),
.B(n_109),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_112),
.B(n_109),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_116),
.Y(n_196)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_132),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_113),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_144),
.C(n_147),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_120),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_180),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_179),
.B(n_3),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_122),
.B1(n_111),
.B2(n_109),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_202),
.B1(n_164),
.B2(n_153),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_177),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_159),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_194),
.C(n_198),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_148),
.C(n_109),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_85),
.C(n_116),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_118),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_204),
.C(n_10),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_85),
.B1(n_33),
.B2(n_29),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_169),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_2),
.C(n_3),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_167),
.B(n_162),
.Y(n_216)
);

AOI211xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_171),
.B(n_172),
.C(n_168),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_208),
.B1(n_217),
.B2(n_7),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_200),
.B(n_157),
.Y(n_211)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_215),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_181),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_185),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_216),
.B(n_220),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_174),
.B1(n_156),
.B2(n_170),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_228),
.B1(n_187),
.B2(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_157),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_10),
.B(n_15),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_221),
.A2(n_224),
.B(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_184),
.B(n_2),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_205),
.B(n_190),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_2),
.B(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_226),
.A2(n_229),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_204),
.C(n_192),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_186),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_182),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_240),
.C(n_244),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_202),
.B1(n_189),
.B2(n_194),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_230),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_238),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_221),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_201),
.C(n_7),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_239),
.C(n_242),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_212),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_6),
.C(n_7),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_6),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_236),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_216),
.C(n_220),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_226),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_251),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_223),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_222),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_260),
.C(n_262),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_256),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_211),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_261),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_227),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_244),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_225),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_219),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_263),
.B(n_248),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_257),
.C(n_261),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_237),
.C(n_231),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_243),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_234),
.C(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_208),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_285),
.C(n_271),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_228),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_245),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_284),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_249),
.B1(n_252),
.B2(n_240),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_9),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

AOI221xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_279),
.B1(n_285),
.B2(n_283),
.C(n_269),
.Y(n_287)
);

NAND2x1_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_14),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_264),
.B(n_269),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_16),
.B(n_14),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_11),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_15),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_13),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_294),
.B(n_297),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_296),
.C(n_292),
.Y(n_298)
);

AOI31xp33_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_291),
.A3(n_287),
.B(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_294),
.B(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_15),
.Y(n_303)
);


endmodule