module fake_jpeg_23831_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_1),
.B(n_3),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_0),
.C(n_5),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_17),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_16),
.Y(n_24)
);

OA21x2_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_2),
.B(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_20),
.Y(n_26)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_14),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_29),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_12),
.C(n_17),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_24),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_25),
.C(n_13),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_19),
.B1(n_21),
.B2(n_16),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_16),
.B1(n_8),
.B2(n_11),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_25),
.C(n_20),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_9),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_8),
.B(n_13),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_9),
.C(n_6),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_9),
.B(n_11),
.C(n_37),
.Y(n_41)
);


endmodule