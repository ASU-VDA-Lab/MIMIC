module fake_jpeg_29905_n_544 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_544);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_544;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_59),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_33),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_70),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_17),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_101),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_27),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_99),
.Y(n_134)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_96),
.Y(n_160)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g137 ( 
.A(n_102),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_30),
.B(n_46),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_112),
.B(n_138),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_120),
.B(n_128),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_80),
.B(n_27),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_43),
.B1(n_53),
.B2(n_47),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_153),
.B1(n_105),
.B2(n_49),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_71),
.B(n_30),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_82),
.A2(n_28),
.B1(n_21),
.B2(n_40),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_139),
.B(n_163),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_54),
.B(n_28),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_63),
.B(n_21),
.Y(n_144)
);

BUFx2_ASAP7_75t_R g150 ( 
.A(n_85),
.Y(n_150)
);

INVx2_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_155),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_84),
.A2(n_47),
.B1(n_29),
.B2(n_45),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_103),
.B1(n_102),
.B2(n_40),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_154),
.A2(n_79),
.B1(n_22),
.B2(n_38),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_90),
.A2(n_46),
.B(n_50),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_90),
.A2(n_50),
.B(n_45),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_47),
.Y(n_179)
);

HAxp5_ASAP7_75t_SL g163 ( 
.A(n_105),
.B(n_33),
.CON(n_163),
.SN(n_163)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_210),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_169),
.A2(n_209),
.B1(n_213),
.B2(n_216),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_130),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_170),
.Y(n_230)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_172),
.Y(n_264)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_174),
.Y(n_261)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_178),
.B(n_180),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_179),
.A2(n_221),
.B(n_182),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_116),
.B(n_48),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

CKINVDCx12_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

INVx6_ASAP7_75t_SL g238 ( 
.A(n_184),
.Y(n_238)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_71),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_186),
.B(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_108),
.B(n_41),
.Y(n_187)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_41),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_189),
.B(n_196),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_190),
.B(n_224),
.Y(n_274)
);

BUFx16f_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_137),
.A2(n_76),
.B1(n_97),
.B2(n_62),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_48),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_202),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_19),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_111),
.B(n_19),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_68),
.B1(n_49),
.B2(n_81),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_109),
.Y(n_205)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_111),
.A2(n_49),
.B1(n_65),
.B2(n_106),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_129),
.B(n_93),
.C(n_32),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_107),
.Y(n_260)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_215),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_49),
.B1(n_34),
.B2(n_38),
.Y(n_213)
);

CKINVDCx12_ASAP7_75t_R g214 ( 
.A(n_166),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_217),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_134),
.B(n_34),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

CKINVDCx12_ASAP7_75t_R g218 ( 
.A(n_166),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_222),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_131),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_223),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_166),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_148),
.B(n_22),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_158),
.A2(n_66),
.B1(n_75),
.B2(n_69),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_127),
.B1(n_122),
.B2(n_140),
.Y(n_265)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_161),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_226),
.A2(n_143),
.B1(n_140),
.B2(n_57),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_164),
.B1(n_165),
.B2(n_132),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_227),
.A2(n_258),
.B1(n_267),
.B2(n_273),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_228),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_L g229 ( 
.A1(n_216),
.A2(n_165),
.B1(n_115),
.B2(n_136),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_240),
.B1(n_265),
.B2(n_268),
.Y(n_278)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_180),
.B(n_153),
.CI(n_133),
.CON(n_237),
.SN(n_237)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_237),
.B(n_51),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_177),
.A2(n_219),
.B1(n_190),
.B2(n_195),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_125),
.B(n_152),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_247),
.B(n_260),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_219),
.A2(n_171),
.B1(n_147),
.B2(n_198),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_201),
.A2(n_147),
.B1(n_115),
.B2(n_55),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_199),
.A2(n_67),
.B1(n_61),
.B2(n_143),
.Y(n_273)
);

OA22x2_ASAP7_75t_SL g275 ( 
.A1(n_237),
.A2(n_183),
.B1(n_193),
.B2(n_200),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_275),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_276),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_211),
.B1(n_208),
.B2(n_226),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_277),
.A2(n_291),
.B1(n_308),
.B2(n_229),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_178),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_279),
.B(n_281),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_238),
.Y(n_280)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_203),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_286),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_203),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_285),
.B(n_299),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_212),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_243),
.A2(n_200),
.B1(n_272),
.B2(n_254),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_287),
.A2(n_310),
.B1(n_217),
.B2(n_192),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_295),
.Y(n_339)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_181),
.B1(n_174),
.B2(n_207),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_227),
.B(n_210),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_292),
.A2(n_122),
.B(n_266),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_293),
.B(n_297),
.Y(n_334)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_294),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_223),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_261),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_296),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_270),
.Y(n_297)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_301),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_245),
.B(n_232),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_236),
.B(n_185),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_305),
.Y(n_335)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_247),
.B(n_191),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_304),
.Y(n_343)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g305 ( 
.A(n_228),
.B(n_176),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_250),
.B(n_220),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_237),
.B(n_220),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_316),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_243),
.A2(n_170),
.B1(n_206),
.B2(n_205),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_247),
.B(n_170),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_253),
.B(n_14),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_257),
.B(n_191),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_313),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_230),
.B(n_175),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_273),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_246),
.B(n_14),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_249),
.B(n_172),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_234),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_234),
.C(n_244),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_246),
.C(n_271),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_329),
.C(n_346),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_302),
.A2(n_262),
.B1(n_263),
.B2(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_235),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_323),
.B(n_283),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_259),
.B1(n_267),
.B2(n_266),
.Y(n_325)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_325),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_235),
.C(n_251),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_340),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_331),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_278),
.A2(n_188),
.B1(n_248),
.B2(n_251),
.Y(n_336)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_286),
.C(n_299),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_304),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_307),
.B1(n_277),
.B2(n_291),
.Y(n_338)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_275),
.A2(n_173),
.B1(n_248),
.B2(n_242),
.Y(n_340)
);

OAI32xp33_ASAP7_75t_L g341 ( 
.A1(n_295),
.A2(n_242),
.A3(n_231),
.B1(n_141),
.B2(n_264),
.Y(n_341)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_341),
.Y(n_387)
);

INVx13_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_288),
.A2(n_231),
.B1(n_264),
.B2(n_70),
.Y(n_344)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_197),
.C(n_77),
.Y(n_346)
);

O2A1O1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_309),
.A2(n_77),
.B(n_197),
.C(n_51),
.Y(n_351)
);

O2A1O1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_351),
.A2(n_289),
.B(n_314),
.C(n_306),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_278),
.A2(n_51),
.B1(n_3),
.B2(n_4),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g358 ( 
.A1(n_323),
.A2(n_305),
.B(n_282),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_L g422 ( 
.A1(n_358),
.A2(n_359),
.B(n_324),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_363),
.B(n_380),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_305),
.C(n_293),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_365),
.B(n_374),
.C(n_379),
.Y(n_402)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_354),
.Y(n_366)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_366),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_334),
.B(n_315),
.Y(n_367)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_384),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_312),
.Y(n_371)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_319),
.B(n_280),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_372),
.B(n_375),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_298),
.Y(n_373)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_316),
.C(n_300),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_322),
.B(n_294),
.Y(n_375)
);

OAI32xp33_ASAP7_75t_L g376 ( 
.A1(n_339),
.A2(n_275),
.A3(n_292),
.B1(n_297),
.B2(n_308),
.Y(n_376)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_376),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_298),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_390),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_347),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_378),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_292),
.C(n_275),
.Y(n_379)
);

CKINVDCx10_ASAP7_75t_R g381 ( 
.A(n_349),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_381),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_304),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_389),
.Y(n_393)
);

INVx6_ASAP7_75t_SL g384 ( 
.A(n_353),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_339),
.A2(n_310),
.B(n_296),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_351),
.B(n_343),
.Y(n_394)
);

A2O1A1O1Ixp25_ASAP7_75t_L g389 ( 
.A1(n_333),
.A2(n_294),
.B(n_296),
.C(n_276),
.D(n_301),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_338),
.B(n_51),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_345),
.B1(n_326),
.B2(n_327),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_392),
.A2(n_401),
.B1(n_408),
.B2(n_388),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_394),
.B(n_398),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_348),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_397),
.B(n_399),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_344),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_348),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_328),
.Y(n_400)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_400),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_391),
.A2(n_370),
.B1(n_387),
.B2(n_363),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_328),
.Y(n_407)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_370),
.A2(n_345),
.B1(n_326),
.B2(n_318),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_419),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_333),
.Y(n_412)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_412),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_365),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_413),
.B(n_354),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_343),
.Y(n_414)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_414),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_387),
.A2(n_321),
.B1(n_329),
.B2(n_341),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_417),
.A2(n_357),
.B1(n_361),
.B2(n_376),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_366),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_360),
.B(n_332),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_421),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_332),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_422),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_346),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_3),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_364),
.C(n_368),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_435),
.C(n_440),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_405),
.A2(n_364),
.B(n_385),
.Y(n_426)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_429),
.B(n_443),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_416),
.B(n_384),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_432),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_395),
.B(n_324),
.Y(n_432)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_409),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_434),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_357),
.C(n_355),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_437),
.A2(n_439),
.B1(n_401),
.B2(n_408),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_417),
.A2(n_361),
.B1(n_362),
.B2(n_383),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_355),
.C(n_390),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_403),
.A2(n_362),
.B1(n_385),
.B2(n_389),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_398),
.B1(n_423),
.B2(n_411),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_331),
.C(n_352),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_448),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_404),
.B(n_2),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_447),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_404),
.B(n_2),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_415),
.B(n_2),
.Y(n_448)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_449),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_397),
.B(n_3),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_446),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_445),
.A2(n_396),
.B(n_412),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_454),
.A2(n_456),
.B(n_467),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_455),
.A2(n_460),
.B1(n_429),
.B2(n_441),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_445),
.A2(n_396),
.B(n_403),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_459),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_393),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_439),
.A2(n_392),
.B1(n_394),
.B2(n_418),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_460),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_444),
.A2(n_414),
.B1(n_400),
.B2(n_407),
.Y(n_462)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_462),
.Y(n_475)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_398),
.B1(n_423),
.B2(n_409),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_465),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_445),
.A2(n_393),
.B(n_410),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_433),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_469),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_438),
.Y(n_469)
);

XOR2x2_ASAP7_75t_L g470 ( 
.A(n_438),
.B(n_428),
.Y(n_470)
);

XNOR2x1_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_442),
.Y(n_481)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_466),
.B(n_427),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_484),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_480),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_454),
.A2(n_456),
.B(n_467),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_491),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_489),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_463),
.B(n_425),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_435),
.C(n_440),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_486),
.C(n_490),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_428),
.C(n_437),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_447),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_450),
.Y(n_490)
);

INVx13_ASAP7_75t_L g491 ( 
.A(n_469),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_479),
.A2(n_455),
.B1(n_451),
.B2(n_471),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_493),
.A2(n_476),
.B1(n_490),
.B2(n_489),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_479),
.A2(n_452),
.B1(n_434),
.B2(n_472),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_496),
.A2(n_499),
.B1(n_482),
.B2(n_8),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_470),
.C(n_461),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_498),
.C(n_500),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_458),
.C(n_453),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_475),
.A2(n_488),
.B1(n_487),
.B2(n_453),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_406),
.C(n_5),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_483),
.A2(n_4),
.B(n_5),
.Y(n_501)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_477),
.A2(n_13),
.B(n_5),
.Y(n_502)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_502),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_12),
.C(n_6),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_503),
.B(n_6),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_487),
.B(n_4),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_506),
.B(n_7),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_481),
.A2(n_4),
.B(n_6),
.Y(n_507)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_507),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_514),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_492),
.A2(n_491),
.B(n_477),
.Y(n_509)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_509),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_478),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_511),
.B(n_515),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_517),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_7),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_505),
.A2(n_7),
.B(n_8),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_498),
.A2(n_7),
.B(n_9),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_493),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_525),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_504),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_494),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_526),
.B(n_529),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_494),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_510),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_532),
.B(n_534),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_525),
.A2(n_500),
.B(n_519),
.Y(n_533)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_528),
.B(n_527),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_523),
.B(n_512),
.Y(n_534)
);

AOI322xp5_ASAP7_75t_L g539 ( 
.A1(n_536),
.A2(n_11),
.A3(n_12),
.B1(n_495),
.B2(n_503),
.C1(n_504),
.C2(n_535),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_SL g537 ( 
.A1(n_530),
.A2(n_524),
.B(n_518),
.C(n_521),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_531),
.C(n_514),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_538),
.B(n_539),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_540),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_541),
.A2(n_11),
.B1(n_495),
.B2(n_523),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_11),
.Y(n_543)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_543),
.Y(n_544)
);


endmodule