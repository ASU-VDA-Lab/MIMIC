module real_jpeg_16095_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_7),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_1),
.B(n_114),
.Y(n_113)
);

AOI22x1_ASAP7_75t_L g119 ( 
.A1(n_1),
.A2(n_3),
.B1(n_120),
.B2(n_124),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_1),
.B(n_138),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_2),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_3),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_3),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_3),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_3),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_3),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_4),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_4),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_4),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_4),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_4),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_4),
.B(n_334),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_6),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_6),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_6),
.B(n_68),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_6),
.B(n_114),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_8),
.B(n_54),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_9),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_9),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_9),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_9),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_9),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_9),
.B(n_294),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_10),
.Y(n_329)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_11),
.Y(n_116)
);

BUFx4f_ASAP7_75t_L g156 ( 
.A(n_11),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_54),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_13),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_13),
.B(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_13),
.B(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_14),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_14),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_17),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_17),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_17),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_17),
.B(n_123),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_18),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_18),
.Y(n_150)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_210),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_172),
.B(n_207),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_25),
.B(n_173),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_102),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_64),
.C(n_85),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_27),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_45),
.C(n_56),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_29),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_30),
.B(n_39),
.C(n_43),
.Y(n_129)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_45),
.B(n_56),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_46),
.B(n_52),
.Y(n_232)
);

NOR2x1_ASAP7_75t_R g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_50),
.Y(n_336)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_55),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.C(n_62),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_57),
.A2(n_60),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_57),
.Y(n_219)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_60),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_60),
.B(n_306),
.C(n_308),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_60),
.A2(n_220),
.B1(n_308),
.B2(n_309),
.Y(n_321)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_62),
.B(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_64),
.B(n_85),
.Y(n_175)
);

XOR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_73),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_66),
.B(n_71),
.C(n_73),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_70),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.C(n_82),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_74),
.A2(n_82),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_74),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_78),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_79),
.B(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx13_ASAP7_75t_SL g180 ( 
.A(n_82),
.Y(n_180)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_84),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_86),
.B(n_91),
.C(n_100),
.Y(n_146)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_89),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_96),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_96),
.A2(n_100),
.B1(n_227),
.B2(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_100),
.B(n_223),
.C(n_227),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_144),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_130),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_118),
.C(n_129),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_105),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_113),
.C(n_117),
.Y(n_132)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_118),
.A2(n_119),
.B1(n_129),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_119),
.A2(n_182),
.B(n_190),
.Y(n_181)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_128),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_130)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_134),
.A2(n_135),
.B1(n_200),
.B2(n_201),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_197),
.C(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

XOR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_157),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_155),
.Y(n_292)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_156),
.Y(n_254)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_204),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_204),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_196),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_181),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_272),
.C(n_277),
.Y(n_271)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_197),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_198),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_198),
.A2(n_315),
.B1(n_316),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_237),
.B(n_343),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_235),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_213),
.B(n_235),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_233),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_233),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.C(n_231),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_232),
.Y(n_244)
);

XOR2x2_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_262),
.B(n_342),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_260),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_241),
.B(n_260),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_257),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_243),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_257),
.B1(n_258),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.C(n_250),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

AO22x1_ASAP7_75t_SL g296 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_255),
.Y(n_297)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_284),
.B(n_341),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g341 ( 
.A(n_264),
.B(n_268),
.Y(n_341)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.C(n_280),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_277),
.Y(n_288)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21x1_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_300),
.B(n_340),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_298),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_298),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.C(n_296),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_290),
.B1(n_296),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_293),
.Y(n_307)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_333),
.Y(n_332)
);

AOI21x1_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_312),
.B(n_339),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_305),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_307),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_322),
.B(n_338),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_319),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_332),
.B(n_337),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_330),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_330),
.Y(n_337)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);


endmodule