module fake_jpeg_26432_n_132 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVxp67_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_26),
.Y(n_29)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_27),
.B(n_10),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_15),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_14),
.C(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_46),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_34),
.B(n_29),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_20),
.B1(n_11),
.B2(n_16),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_26),
.B1(n_27),
.B2(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_37),
.B1(n_43),
.B2(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_54),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_70),
.B1(n_26),
.B2(n_30),
.Y(n_87)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_65),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_45),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_71),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_37),
.B1(n_34),
.B2(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_60),
.B1(n_26),
.B2(n_30),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_74),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_76),
.B(n_25),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_19),
.C(n_18),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_12),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_80),
.B1(n_63),
.B2(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_19),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_52),
.B(n_15),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_21),
.C(n_25),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_91),
.C(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_12),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_21),
.C(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_93),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_67),
.C(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_96),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_76),
.B1(n_69),
.B2(n_63),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_64),
.B1(n_30),
.B2(n_14),
.Y(n_98)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_101),
.B(n_100),
.Y(n_108)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_14),
.B(n_25),
.Y(n_101)
);

OA21x2_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_85),
.B(n_91),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_84),
.C(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_25),
.B1(n_21),
.B2(n_3),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_95),
.B(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_92),
.C(n_99),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_113),
.C(n_114),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_105),
.B1(n_109),
.B2(n_21),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_1),
.C(n_5),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_9),
.C(n_2),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_9),
.C(n_3),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_21),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_1),
.B(n_3),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_8),
.C(n_4),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_125),
.Y(n_126)
);

OAI221xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_119),
.C(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_127),
.B(n_6),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_8),
.Y(n_132)
);


endmodule