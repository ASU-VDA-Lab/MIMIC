module fake_jpeg_3465_n_441 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_64),
.Y(n_115)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_27),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g171 ( 
.A(n_59),
.Y(n_171)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_16),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_61),
.A2(n_80),
.B(n_86),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_72),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_77),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_17),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_30),
.B(n_12),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_2),
.B(n_3),
.Y(n_86)
);

BUFx6f_ASAP7_75t_SL g87 ( 
.A(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_29),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_93),
.Y(n_127)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_90),
.Y(n_178)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_28),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_R g95 ( 
.A(n_21),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_95),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_3),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_100),
.Y(n_136)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_32),
.B(n_3),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_20),
.C(n_43),
.Y(n_150)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_105),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_107),
.Y(n_145)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_111),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_55),
.B1(n_33),
.B2(n_41),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_33),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_113),
.Y(n_158)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_56),
.A2(n_21),
.B1(n_53),
.B2(n_45),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_117),
.A2(n_123),
.B1(n_134),
.B2(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_121),
.B(n_151),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_54),
.B1(n_48),
.B2(n_51),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_60),
.A2(n_55),
.B1(n_48),
.B2(n_46),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g238 ( 
.A1(n_125),
.A2(n_154),
.B1(n_165),
.B2(n_169),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_45),
.B1(n_42),
.B2(n_40),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_59),
.A2(n_33),
.B1(n_46),
.B2(n_41),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_135),
.A2(n_140),
.B1(n_141),
.B2(n_147),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_58),
.A2(n_26),
.B1(n_34),
.B2(n_53),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_68),
.A2(n_34),
.B1(n_42),
.B2(n_40),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_96),
.A2(n_39),
.B1(n_36),
.B2(n_20),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_142),
.A2(n_160),
.B1(n_174),
.B2(n_175),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_39),
.B1(n_36),
.B2(n_20),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_150),
.B(n_174),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_4),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_20),
.B1(n_7),
.B2(n_8),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_5),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_155),
.B(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_69),
.B(n_5),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_159),
.B(n_176),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_109),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_65),
.A2(n_9),
.B1(n_11),
.B2(n_84),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_81),
.A2(n_90),
.B1(n_75),
.B2(n_91),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_110),
.A2(n_9),
.B1(n_11),
.B2(n_75),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_103),
.B(n_11),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_106),
.A2(n_11),
.B1(n_71),
.B2(n_95),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_71),
.A2(n_63),
.B1(n_82),
.B2(n_83),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_101),
.A2(n_98),
.B1(n_61),
.B2(n_77),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_80),
.A2(n_21),
.B1(n_32),
.B2(n_25),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_150),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_59),
.A2(n_21),
.B1(n_27),
.B2(n_55),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_125),
.B1(n_146),
.B2(n_131),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_115),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_187),
.Y(n_286)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_127),
.B(n_119),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_189),
.B(n_211),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_192),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_179),
.A2(n_121),
.B1(n_151),
.B2(n_155),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_193),
.A2(n_204),
.B1(n_215),
.B2(n_217),
.Y(n_280)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_199),
.Y(n_246)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_197),
.Y(n_273)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_137),
.A2(n_116),
.B1(n_156),
.B2(n_138),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_205),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_209),
.Y(n_247)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

OR2x4_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_158),
.Y(n_208)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_203),
.B(n_216),
.C(n_193),
.Y(n_254)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_120),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_214),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_163),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_145),
.B(n_174),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_234),
.B(n_221),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_146),
.A2(n_161),
.B(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_213),
.B(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_116),
.A2(n_164),
.B1(n_148),
.B2(n_161),
.Y(n_217)
);

BUFx12_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_218),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_138),
.B(n_156),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_132),
.A2(n_164),
.B1(n_149),
.B2(n_143),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_230),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_128),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_224),
.Y(n_258)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_153),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_225),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_168),
.B(n_143),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_226),
.B(n_231),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_233),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_228),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_229),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_149),
.A2(n_168),
.B1(n_118),
.B2(n_122),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_114),
.B(n_120),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_114),
.B(n_118),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_232),
.B(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_166),
.Y(n_244)
);

INVx13_ASAP7_75t_L g235 ( 
.A(n_128),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_139),
.B(n_152),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_152),
.A2(n_174),
.B1(n_139),
.B2(n_166),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_188),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_131),
.B(n_177),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_239),
.B(n_240),
.Y(n_284)
);

CKINVDCx6p67_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

CKINVDCx12_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_200),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_270),
.C(n_278),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_264),
.B1(n_243),
.B2(n_247),
.Y(n_295)
);

NOR2x1_ASAP7_75t_R g311 ( 
.A(n_254),
.B(n_256),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_266),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g260 ( 
.A1(n_212),
.A2(n_219),
.B(n_221),
.C(n_186),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_260),
.B(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_204),
.B(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_281),
.Y(n_293)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_191),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_219),
.A2(n_186),
.B(n_191),
.C(n_238),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_238),
.C(n_209),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_227),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_185),
.C(n_229),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_207),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_225),
.B(n_183),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_218),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_205),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_287),
.B(n_302),
.Y(n_338)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g289 ( 
.A(n_250),
.B(n_205),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_310),
.Y(n_325)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_251),
.Y(n_291)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_251),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_294),
.Y(n_339)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_295),
.A2(n_297),
.B1(n_298),
.B2(n_317),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_255),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_252),
.A2(n_227),
.B1(n_235),
.B2(n_201),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_278),
.A2(n_187),
.B1(n_197),
.B2(n_201),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_304),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_280),
.A2(n_218),
.B1(n_247),
.B2(n_260),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_303),
.A2(n_309),
.B1(n_279),
.B2(n_261),
.Y(n_330)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_254),
.B(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_305),
.B(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_259),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_308),
.Y(n_336)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

AO22x1_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_268),
.B1(n_258),
.B2(n_267),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_257),
.A2(n_269),
.B(n_242),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_318),
.B(n_320),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_254),
.B(n_276),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_253),
.Y(n_329)
);

OA22x2_ASAP7_75t_L g315 ( 
.A1(n_280),
.A2(n_266),
.B1(n_243),
.B2(n_270),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_275),
.B(n_271),
.C(n_262),
.Y(n_327)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_319),
.B1(n_272),
.B2(n_245),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_244),
.A2(n_257),
.B1(n_282),
.B2(n_284),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_259),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_249),
.B(n_245),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_282),
.A2(n_242),
.B1(n_274),
.B2(n_271),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_287),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_323),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_268),
.B(n_258),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_324),
.A2(n_332),
.B(n_343),
.Y(n_365)
);

AO21x1_ASAP7_75t_L g354 ( 
.A1(n_327),
.A2(n_328),
.B(n_330),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_277),
.B1(n_261),
.B2(n_279),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_344),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_253),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_337),
.C(n_291),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_307),
.A2(n_277),
.B(n_262),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_246),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_295),
.A2(n_273),
.B1(n_275),
.B2(n_286),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_340),
.A2(n_296),
.B1(n_300),
.B2(n_310),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_313),
.A2(n_246),
.B(n_265),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_289),
.A2(n_265),
.B(n_273),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_263),
.B(n_286),
.Y(n_346)
);

AOI221xp5_ASAP7_75t_L g369 ( 
.A1(n_346),
.A2(n_263),
.B1(n_288),
.B2(n_294),
.C(n_344),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_303),
.A2(n_263),
.B1(n_293),
.B2(n_304),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_347),
.A2(n_306),
.B1(n_293),
.B2(n_320),
.Y(n_359)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_339),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_348),
.B(n_351),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_349),
.A2(n_360),
.B1(n_366),
.B2(n_369),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_333),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_334),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_355),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_353),
.A2(n_324),
.B(n_343),
.Y(n_374)
);

AO22x1_ASAP7_75t_L g355 ( 
.A1(n_327),
.A2(n_299),
.B1(n_311),
.B2(n_317),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_364),
.Y(n_371)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_362),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_359),
.A2(n_335),
.B1(n_323),
.B2(n_333),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_321),
.A2(n_298),
.B1(n_315),
.B2(n_292),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_312),
.C(n_315),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_367),
.C(n_336),
.Y(n_376)
);

AOI322xp5_ASAP7_75t_SL g362 ( 
.A1(n_338),
.A2(n_308),
.A3(n_318),
.B1(n_309),
.B2(n_312),
.C1(n_315),
.C2(n_316),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_368),
.Y(n_379)
);

XNOR2x2_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_312),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_315),
.B1(n_296),
.B2(n_290),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_326),
.B(n_337),
.C(n_331),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_341),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_329),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_372),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_364),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_373),
.A2(n_374),
.B1(n_382),
.B2(n_365),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_377),
.C(n_378),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_335),
.C(n_345),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_360),
.C(n_350),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_365),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_385),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_366),
.A2(n_323),
.B1(n_325),
.B2(n_346),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_345),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_359),
.Y(n_394)
);

NOR3xp33_ASAP7_75t_SL g385 ( 
.A(n_348),
.B(n_325),
.C(n_338),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_SL g386 ( 
.A(n_353),
.B(n_322),
.C(n_327),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_386),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_371),
.B(n_355),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_394),
.C(n_401),
.Y(n_403)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_389),
.Y(n_402)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_383),
.Y(n_390)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_351),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_391),
.B(n_392),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_382),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_397),
.A2(n_380),
.B1(n_384),
.B2(n_327),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_373),
.A2(n_349),
.B1(n_328),
.B2(n_330),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_399),
.B(n_400),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_352),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_371),
.B(n_350),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_406),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_396),
.A2(n_354),
.B(n_374),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_397),
.A2(n_375),
.B1(n_386),
.B2(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_408),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_391),
.A2(n_354),
.B(n_357),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_400),
.A2(n_357),
.B1(n_327),
.B2(n_354),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_394),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_332),
.B(n_377),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_412),
.A2(n_407),
.B(n_405),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_398),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_416),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_398),
.C(n_393),
.Y(n_416)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_417),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_378),
.C(n_376),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_418),
.B(n_420),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_419),
.A2(n_411),
.B(n_410),
.Y(n_427)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

BUFx24_ASAP7_75t_SL g421 ( 
.A(n_409),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_389),
.C(n_342),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_415),
.A2(n_404),
.B1(n_412),
.B2(n_408),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_428),
.Y(n_433)
);

INVx11_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_368),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_427),
.A2(n_415),
.B(n_416),
.Y(n_430)
);

BUFx4f_ASAP7_75t_SL g429 ( 
.A(n_422),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_432),
.C(n_427),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_393),
.C(n_403),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_431),
.B(n_422),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_436),
.B1(n_432),
.B2(n_425),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_423),
.C(n_433),
.Y(n_437)
);

AOI21xp33_ASAP7_75t_SL g439 ( 
.A1(n_437),
.A2(n_438),
.B(n_424),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_437),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_426),
.Y(n_441)
);


endmodule