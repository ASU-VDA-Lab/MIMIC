module fake_jpeg_23135_n_240 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_240);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_28),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_29),
.B1(n_22),
.B2(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_55),
.B1(n_61),
.B2(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_29),
.B1(n_26),
.B2(n_30),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_54),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_29),
.B1(n_26),
.B2(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_15),
.B1(n_28),
.B2(n_17),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_18),
.B1(n_19),
.B2(n_17),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_32),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_72),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_73),
.B1(n_38),
.B2(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_78),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_76),
.B(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_32),
.C(n_41),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_43),
.C(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_41),
.B1(n_36),
.B2(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_34),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_21),
.B1(n_36),
.B2(n_27),
.Y(n_83)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_56),
.B1(n_62),
.B2(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_93),
.B1(n_97),
.B2(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_90),
.B(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_38),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_31),
.B(n_16),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_96),
.B(n_84),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_56),
.B1(n_53),
.B2(n_36),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_60),
.C(n_39),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_73),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_39),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_106),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_39),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_103),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_101),
.C(n_92),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_69),
.B1(n_76),
.B2(n_74),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_115),
.B1(n_127),
.B2(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_67),
.B1(n_71),
.B2(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_118),
.B(n_123),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_30),
.B(n_27),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_124),
.B(n_104),
.Y(n_140)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_82),
.B1(n_72),
.B2(n_39),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_89),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_149),
.B1(n_146),
.B2(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_147),
.C(n_150),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_133),
.B(n_25),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_102),
.A3(n_106),
.B1(n_97),
.B2(n_100),
.C1(n_104),
.C2(n_63),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_47),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_64),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_146),
.B1(n_144),
.B2(n_138),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_100),
.B(n_103),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_144),
.B(n_145),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_87),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_113),
.B(n_115),
.Y(n_145)
);

AND2x4_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_103),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_0),
.B(n_2),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_108),
.B1(n_109),
.B2(n_87),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_103),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_86),
.B1(n_82),
.B2(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_159),
.B1(n_131),
.B2(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_157),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_120),
.C(n_128),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_150),
.C(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_64),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_47),
.B1(n_25),
.B2(n_63),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_162),
.B1(n_167),
.B2(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_47),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_149),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_139),
.B(n_141),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_160),
.B(n_144),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_175),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_151),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_180),
.B(n_182),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_141),
.C(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_185),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_133),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_139),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_187),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_135),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_181),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_200),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_191),
.B1(n_196),
.B2(n_190),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_154),
.B1(n_155),
.B2(n_161),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_184),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_175),
.C(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_187),
.A2(n_163),
.B(n_155),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_201),
.B(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_166),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_161),
.B(n_156),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_203),
.B(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_204),
.B(n_198),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_207),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_171),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_170),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_209),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_154),
.C(n_172),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_211),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_183),
.B(n_159),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_165),
.B1(n_173),
.B2(n_168),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_212),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_204),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_0),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_2),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_2),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_3),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_210),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_207),
.B1(n_4),
.B2(n_5),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_227),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_226),
.A3(n_225),
.B1(n_219),
.B2(n_217),
.C1(n_221),
.C2(n_12),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_217),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_6),
.C2(n_12),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_235),
.A3(n_229),
.B1(n_9),
.B2(n_11),
.C1(n_13),
.C2(n_8),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_13),
.C2(n_231),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_11),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_236),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_13),
.Y(n_240)
);


endmodule