module fake_jpeg_18058_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx4_ASAP7_75t_SL g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_1),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_11),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_2),
.B(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_21),
.B1(n_13),
.B2(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_12),
.B(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_8),
.B1(n_7),
.B2(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_19),
.A2(n_8),
.B1(n_3),
.B2(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_27),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_24),
.Y(n_38)
);

BUFx24_ASAP7_75t_SL g39 ( 
.A(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_32),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_44),
.B(n_45),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_31),
.B(n_23),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_30),
.C(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

AOI21x1_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_47),
.B(n_41),
.Y(n_49)
);


endmodule