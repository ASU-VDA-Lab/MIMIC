module real_jpeg_19243_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_332, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_332;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_176;
wire n_215;
wire n_166;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_0),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_95),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_95),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_0),
.A2(n_40),
.B1(n_41),
.B2(n_95),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_23),
.B1(n_44),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_1),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_85),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_85),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_85),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_91),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_91),
.Y(n_251)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_5),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_97),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_97),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_6),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_29),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_16),
.B(n_44),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_100),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_78),
.B1(n_81),
.B2(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_6),
.B(n_55),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_31),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_7),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_7),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_60),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_60),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_255)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_11),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_102),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_102),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_102),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_63),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_63),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_63),
.Y(n_274)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_51),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_14),
.A2(n_31),
.A3(n_41),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_16),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_16),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

BUFx3_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_325),
.B(n_328),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_68),
.B(n_324),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_21),
.B(n_34),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_21),
.B(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_21),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_27),
.Y(n_28)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_24),
.B(n_100),
.CON(n_99),
.SN(n_99)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_26),
.A2(n_29),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_26),
.A2(n_29),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_26),
.A2(n_29),
.B(n_32),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_31),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_28),
.A2(n_30),
.B1(n_99),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_30),
.B(n_100),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_64),
.C(n_66),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_35),
.A2(n_36),
.B1(n_320),
.B2(n_322),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_47),
.C(n_56),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_37),
.A2(n_291),
.B1(n_292),
.B2(n_294),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_37),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_37),
.A2(n_47),
.B1(n_294),
.B2(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_43),
.B(n_46),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_38),
.A2(n_43),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_38),
.A2(n_43),
.B1(n_84),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_38),
.A2(n_43),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_38),
.A2(n_43),
.B1(n_152),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_38),
.A2(n_43),
.B1(n_174),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_38),
.A2(n_43),
.B1(n_90),
.B2(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_38),
.A2(n_43),
.B1(n_86),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_38),
.A2(n_43),
.B1(n_228),
.B2(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_38),
.A2(n_43),
.B1(n_46),
.B2(n_261),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_40),
.B(n_51),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_41),
.A2(n_42),
.B(n_100),
.C(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_43),
.B(n_100),
.Y(n_155)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_45),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_47),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_49),
.A2(n_54),
.B(n_55),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_55),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_49),
.A2(n_55),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_53),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_53),
.B1(n_96),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_50),
.A2(n_53),
.B1(n_126),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_50),
.A2(n_53),
.B1(n_110),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_50),
.A2(n_53),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_56),
.A2(n_57),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_61),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_58),
.A2(n_61),
.B1(n_108),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_58),
.A2(n_61),
.B1(n_235),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_66),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_317),
.B(n_323),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_286),
.A3(n_309),
.B1(n_315),
.B2(n_316),
.C(n_332),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_265),
.B(n_285),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_241),
.B(n_264),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_132),
.B(n_217),
.C(n_240),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_117),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_74),
.B(n_117),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_103),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_76),
.B(n_87),
.C(n_103),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_77),
.B(n_83),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_79),
.B1(n_116),
.B2(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_78),
.A2(n_81),
.B1(n_142),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_78),
.A2(n_144),
.B1(n_161),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_78),
.A2(n_131),
.B1(n_161),
.B2(n_176),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_78),
.A2(n_82),
.B1(n_161),
.B2(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_78),
.A2(n_81),
.B(n_226),
.Y(n_259)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.C(n_98),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_105),
.B(n_111),
.C(n_112),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_109),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_115),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_129),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_124),
.B(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_128),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_216),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_211),
.B(n_215),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_197),
.B(n_210),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_178),
.B(n_196),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_166),
.B(n_177),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_153),
.B(n_165),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_145),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_149),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_158),
.B(n_164),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_173),
.C(n_175),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B1(n_194),
.B2(n_195),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_198),
.B(n_199),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_207),
.C(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_219),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_239),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_229),
.B2(n_230),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_230),
.C(n_239),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_233),
.C(n_238),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_238),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_243),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_263),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_256),
.B2(n_257),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_257),
.C(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_249),
.C(n_253),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_251),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_259),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_259),
.A2(n_277),
.B1(n_280),
.B2(n_333),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_283),
.B2(n_284),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_276),
.C(n_284),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B(n_275),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_274),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_288),
.C(n_299),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_275),
.A2(n_288),
.B1(n_289),
.B2(n_314),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_275),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_301),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_301),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_289)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_295),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_295),
.A2(n_298),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_303),
.C(n_308),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_299),
.A2(n_300),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_319),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_320),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule