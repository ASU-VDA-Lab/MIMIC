module fake_jpeg_21456_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_20),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_68),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_45),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_58),
.B1(n_52),
.B2(n_57),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_91),
.B1(n_95),
.B2(n_53),
.Y(n_99)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_93),
.Y(n_98)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_61),
.B1(n_47),
.B2(n_54),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_51),
.B(n_50),
.C(n_44),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_61),
.B1(n_53),
.B2(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_65),
.B1(n_62),
.B2(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_97),
.B(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_106),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_19),
.B1(n_41),
.B2(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_0),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_18),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_14),
.B1(n_36),
.B2(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_1),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_2),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_105),
.Y(n_120)
);

OAI322xp33_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_122),
.A3(n_123),
.B1(n_23),
.B2(n_42),
.C1(n_32),
.C2(n_31),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_104),
.B1(n_101),
.B2(n_105),
.Y(n_121)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_112),
.B(n_119),
.C(n_115),
.D(n_117),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_13),
.B(n_34),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.C(n_121),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_113),
.B1(n_9),
.B2(n_30),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_8),
.C(n_29),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_24),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_12),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_2),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_3),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_3),
.C(n_4),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);


endmodule