module fake_jpeg_24516_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_18),
.B1(n_13),
.B2(n_20),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_19),
.B1(n_14),
.B2(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_29),
.A2(n_24),
.B(n_17),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_1),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_42),
.B(n_16),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_45),
.B1(n_17),
.B2(n_15),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_43),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_32),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_25),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_21),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_15),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_30),
.C(n_3),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_54),
.C(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_23),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_22),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_59),
.B1(n_63),
.B2(n_46),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_2),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_16),
.B1(n_3),
.B2(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_34),
.B1(n_42),
.B2(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_70),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_75),
.B1(n_63),
.B2(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_47),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_81),
.C(n_73),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_70),
.C(n_49),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_83),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_71),
.B(n_59),
.Y(n_85)
);

AOI222xp33_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_72),
.B1(n_49),
.B2(n_54),
.C1(n_58),
.C2(n_61),
.Y(n_86)
);

NAND4xp25_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.C(n_78),
.D(n_81),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_46),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_88),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_92),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_60),
.B1(n_67),
.B2(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_11),
.C(n_7),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_90),
.B1(n_96),
.B2(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_100),
.Y(n_102)
);


endmodule