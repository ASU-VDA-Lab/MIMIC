module real_jpeg_17455_n_19 (n_17, n_8, n_0, n_141, n_2, n_132, n_139, n_142, n_10, n_137, n_9, n_12, n_135, n_134, n_6, n_136, n_133, n_11, n_14, n_131, n_138, n_7, n_18, n_3, n_5, n_4, n_1, n_140, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_141;
input n_2;
input n_132;
input n_139;
input n_142;
input n_10;
input n_137;
input n_9;
input n_12;
input n_135;
input n_134;
input n_6;
input n_136;
input n_133;
input n_11;
input n_14;
input n_131;
input n_138;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_140;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_0),
.B(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_1),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_4),
.B(n_73),
.C(n_98),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_5),
.B(n_77),
.C(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_6),
.B(n_57),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_7),
.A2(n_75),
.B(n_85),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_10),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_14),
.B(n_42),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_16),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_16),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_17),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_SL g106 ( 
.A1(n_18),
.A2(n_54),
.A3(n_67),
.B1(n_70),
.B2(n_107),
.C1(n_109),
.C2(n_142),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_23),
.B(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_79),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_121),
.B(n_127),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_36),
.B(n_119),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_30),
.B(n_35),
.Y(n_120)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_112),
.B(n_116),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI31xp67_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_47),
.A3(n_72),
.B(n_103),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR3xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.C(n_60),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_62),
.C(n_108),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_60),
.A3(n_104),
.B1(n_105),
.B2(n_106),
.C(n_141),
.Y(n_103)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_92),
.C(n_93),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.C(n_81),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_131),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_132),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_133),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_134),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_135),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_136),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_137),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_138),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_139),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_140),
.Y(n_99)
);


endmodule