module fake_jpeg_19757_n_202 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_3),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_18),
.B1(n_15),
.B2(n_27),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_31),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_50),
.B1(n_43),
.B2(n_47),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_27),
.B1(n_14),
.B2(n_24),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_27),
.B1(n_18),
.B2(n_21),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_60),
.B1(n_69),
.B2(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_54),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_24),
.B(n_22),
.Y(n_53)
);

BUFx24_ASAP7_75t_SL g86 ( 
.A(n_53),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_21),
.B1(n_25),
.B2(n_15),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_25),
.B1(n_16),
.B2(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_13),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx2_ASAP7_75t_SL g65 ( 
.A(n_41),
.Y(n_65)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_16),
.B(n_1),
.C(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_13),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_0),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_87),
.Y(n_103)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_80),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_46),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_16),
.B(n_48),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_88),
.B(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_48),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_16),
.B(n_41),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_2),
.C(n_4),
.Y(n_112)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_70),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_77),
.A2(n_71),
.B(n_69),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_80),
.B(n_75),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_98),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_69),
.B1(n_68),
.B2(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_111),
.B1(n_114),
.B2(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_55),
.C(n_54),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_73),
.C(n_97),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_106),
.B(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_110),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_70),
.B1(n_61),
.B2(n_45),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_113),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_4),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_5),
.B(n_6),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_73),
.B(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_88),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_134),
.C(n_101),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_132),
.B(n_136),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_81),
.B1(n_90),
.B2(n_91),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_127),
.B1(n_98),
.B2(n_109),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_84),
.B1(n_78),
.B2(n_79),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_79),
.B(n_96),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_115),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_78),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_105),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_78),
.B(n_79),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_141),
.B1(n_149),
.B2(n_126),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_143),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_144),
.B1(n_118),
.B2(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_98),
.C(n_99),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_122),
.C(n_127),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_112),
.B1(n_102),
.B2(n_116),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_7),
.B(n_10),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_151),
.B(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_146),
.C(n_149),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_126),
.B1(n_135),
.B2(n_130),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_165),
.B1(n_148),
.B2(n_153),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_140),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_172),
.C(n_173),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_152),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_143),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_141),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_155),
.B(n_154),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_177),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_163),
.B(n_157),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_136),
.B(n_123),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_179),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_156),
.C(n_121),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_184),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_131),
.B1(n_121),
.B2(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_131),
.B1(n_133),
.B2(n_11),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_188),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_133),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_182),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_184),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_190),
.C(n_182),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_R g196 ( 
.A(n_193),
.B(n_187),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_196),
.A2(n_79),
.B(n_10),
.C(n_11),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.C(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_199),
.B(n_7),
.Y(n_200)
);

NAND2x1p5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_12),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_12),
.Y(n_202)
);


endmodule