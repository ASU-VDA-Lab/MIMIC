module real_jpeg_3147_n_16 (n_5, n_4, n_8, n_0, n_12, n_272, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_272;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_166;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_205;
wire n_61;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_37),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_1),
.A2(n_37),
.B1(n_70),
.B2(n_71),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_1),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_52),
.B1(n_59),
.B2(n_60),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_52),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_70),
.B1(n_71),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_3),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_125),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_125),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_125),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_5),
.A2(n_70),
.B1(n_71),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_76),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_76),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_76),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_70),
.B1(n_71),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_155),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_155),
.Y(n_215)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_33),
.B1(n_70),
.B2(n_71),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_11),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_12),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_12),
.B(n_31),
.C(n_46),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_12),
.B(n_28),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_12),
.B(n_96),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_12),
.B(n_59),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_12),
.A2(n_59),
.B(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_12),
.B(n_78),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_12),
.A2(n_70),
.B(n_242),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_14),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_50),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_108),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_80),
.B2(n_81),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.C(n_67),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_22),
.A2(n_23),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_26),
.A2(n_38),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_31),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_27),
.A2(n_29),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_27),
.A2(n_86),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_27),
.A2(n_35),
.B(n_148),
.Y(n_232)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_28),
.B(n_36),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_28),
.A2(n_38),
.B1(n_120),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_38),
.B1(n_144),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_28),
.A2(n_38),
.B1(n_186),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_29),
.A2(n_86),
.B(n_121),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_31),
.B(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_39),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_40),
.A2(n_51),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_40),
.A2(n_48),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_40),
.A2(n_94),
.B(n_100),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_95),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_41),
.A2(n_96),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_41),
.A2(n_96),
.B1(n_171),
.B2(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_41),
.A2(n_99),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_44),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_43),
.B(n_55),
.Y(n_207)
);

CKINVDCx6p67_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_44),
.B(n_176),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_44),
.A2(n_56),
.A3(n_59),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_48),
.A2(n_49),
.B(n_102),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_53),
.B(n_67),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B(n_62),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_54),
.B(n_144),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_54),
.A2(n_65),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_54),
.A2(n_65),
.B1(n_150),
.B2(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_66)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_60),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_59),
.B(n_71),
.C(n_73),
.Y(n_145)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_72),
.B(n_143),
.C(n_145),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_63),
.B(n_105),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_64),
.A2(n_105),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_65),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_75),
.B(n_77),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_68),
.A2(n_74),
.B1(n_75),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_68),
.A2(n_74),
.B1(n_124),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_68),
.A2(n_74),
.B1(n_154),
.B2(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_71),
.B(n_144),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_97),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_92),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_84),
.A2(n_85),
.B1(n_93),
.B2(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_119),
.B(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_103),
.B(n_107),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_103),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_105),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_114),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_109),
.B(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_114),
.A2(n_115),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.C(n_126),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_117),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_118),
.B(n_122),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_126),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_159),
.B(n_270),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_156),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_133),
.B(n_156),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.C(n_139),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_134),
.B(n_137),
.Y(n_254)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_139),
.B(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.C(n_153),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_140),
.B(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_149),
.B(n_153),
.Y(n_258)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI321xp33_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_252),
.A3(n_262),
.B1(n_268),
.B2(n_269),
.C(n_272),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_235),
.B(n_251),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_217),
.B(n_234),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_199),
.B(n_216),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_180),
.B(n_198),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_173),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_173),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_170),
.C(n_201),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_192),
.B(n_197),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_187),
.B(n_191),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_190),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_202),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_210),
.C(n_213),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_233),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_233),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_230),
.C(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_237),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_246),
.B2(n_247),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_248),
.C(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_244),
.C(n_245),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.C(n_261),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_257),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);


endmodule