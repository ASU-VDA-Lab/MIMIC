module fake_jpeg_7077_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_25),
.Y(n_32)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2x1p5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_10),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_15),
.C(n_13),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_31),
.Y(n_53)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_48),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_48),
.B1(n_39),
.B2(n_42),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_33),
.C(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_29),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_65),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_67),
.C(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_52),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_43),
.C(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_76),
.A2(n_45),
.B(n_18),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_86),
.B1(n_20),
.B2(n_50),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_28),
.B(n_18),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_85),
.B(n_69),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_49),
.B(n_11),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_38),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_91),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_85),
.B(n_19),
.C(n_10),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_78),
.B1(n_23),
.B2(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_78),
.B1(n_23),
.B2(n_26),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_25),
.C(n_10),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_89),
.B1(n_93),
.B2(n_82),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_101),
.C(n_102),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_92),
.B(n_19),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_98),
.B(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_3),
.C(n_4),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_9),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_3),
.B(n_7),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_1),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_103),
.C(n_107),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_1),
.B(n_2),
.Y(n_110)
);


endmodule