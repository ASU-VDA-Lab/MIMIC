module fake_jpeg_8065_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_39),
.Y(n_60)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_7),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_34),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_50),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_21),
.B1(n_25),
.B2(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_63),
.B1(n_31),
.B2(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_19),
.B1(n_31),
.B2(n_18),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_39),
.A2(n_21),
.B1(n_35),
.B2(n_32),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_35),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_79),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_21),
.B1(n_35),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_83),
.B1(n_84),
.B2(n_52),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_62),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_40),
.C(n_46),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_44),
.A3(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_22),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_39),
.B1(n_44),
.B2(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_33),
.B1(n_17),
.B2(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_91),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_40),
.B(n_37),
.C(n_36),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_92),
.B1(n_53),
.B2(n_52),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_39),
.B1(n_30),
.B2(n_22),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_20),
.B1(n_29),
.B2(n_59),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_97),
.Y(n_127)
);

AOI22x1_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_62),
.B1(n_22),
.B2(n_28),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_70),
.B(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_102),
.B1(n_117),
.B2(n_85),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_69),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_77),
.C(n_65),
.Y(n_142)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_114),
.Y(n_129)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_80),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_111),
.Y(n_134)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_40),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_59),
.B1(n_28),
.B2(n_30),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_113),
.B1(n_100),
.B2(n_96),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_128),
.B1(n_140),
.B2(n_141),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_SL g121 ( 
.A(n_118),
.B(n_73),
.C(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_77),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_76),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_135),
.C(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_70),
.B1(n_82),
.B2(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_130),
.B(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_75),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_138),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_76),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_75),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_115),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_36),
.C(n_37),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_152),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_155),
.B(n_162),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_103),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_156),
.C(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_127),
.B1(n_139),
.B2(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_153),
.B1(n_160),
.B2(n_64),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_72),
.B1(n_78),
.B2(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_138),
.B(n_134),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_46),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_40),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_72),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_90),
.B1(n_61),
.B2(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_65),
.B(n_64),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_116),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_125),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_34),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.C(n_37),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_129),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_1),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_121),
.C(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_184),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_141),
.B(n_142),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_7),
.B(n_14),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_141),
.B1(n_109),
.B2(n_61),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_188),
.B1(n_145),
.B2(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_182),
.C(n_183),
.Y(n_190)
);

OAI321xp33_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_30),
.A3(n_28),
.B1(n_37),
.B2(n_110),
.C(n_34),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_181),
.A2(n_162),
.B(n_165),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_65),
.C(n_55),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_55),
.C(n_28),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_55),
.C(n_2),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_166),
.C(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_7),
.B1(n_15),
.B2(n_3),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_157),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_192),
.C(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_193),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_160),
.B1(n_143),
.B2(n_167),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_174),
.B(n_4),
.C(n_5),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_156),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_150),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.C(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_150),
.C(n_148),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_171),
.B1(n_187),
.B2(n_169),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_201),
.A2(n_173),
.B(n_187),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_205),
.Y(n_211)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_1),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_186),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_210),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_2),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_190),
.C(n_198),
.Y(n_222)
);

INVxp33_ASAP7_75t_SL g214 ( 
.A(n_200),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_206),
.Y(n_223)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_190),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_172),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_189),
.C(n_192),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_170),
.B1(n_179),
.B2(n_168),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_201),
.B1(n_194),
.B2(n_179),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_202),
.B1(n_205),
.B2(n_199),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_224),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_229),
.C(n_207),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_223),
.A2(n_9),
.B(n_4),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_216),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_230),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_209),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_207),
.C(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_2),
.C(n_6),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_211),
.C(n_219),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_233),
.B(n_234),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_210),
.Y(n_233)
);

NAND4xp25_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_217),
.C(n_208),
.D(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_238),
.C(n_9),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_222),
.B1(n_4),
.B2(n_5),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_240),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_244),
.C(n_12),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_243)
);

AOI21x1_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_14),
.B(n_16),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_11),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_237),
.B(n_236),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_247),
.C(n_245),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_243),
.B1(n_240),
.B2(n_16),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_249),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_250),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_235),
.B(n_251),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_252),
.Y(n_255)
);


endmodule