module fake_jpeg_18906_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_45),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_27),
.B1(n_29),
.B2(n_17),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_32),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_60),
.C(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_25),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_27),
.B1(n_29),
.B2(n_17),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_46),
.B1(n_18),
.B2(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_29),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_18),
.B1(n_16),
.B2(n_22),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_70),
.B(n_77),
.Y(n_133)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_72),
.B(n_80),
.Y(n_134)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_82),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_21),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_104),
.Y(n_125)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_21),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_96),
.Y(n_135)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_43),
.B1(n_40),
.B2(n_50),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_106),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_49),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_43),
.B1(n_40),
.B2(n_50),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_45),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_45),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_50),
.B1(n_93),
.B2(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_127),
.B1(n_81),
.B2(n_26),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_132),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_43),
.B1(n_16),
.B2(n_22),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_102),
.B1(n_86),
.B2(n_95),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_23),
.B1(n_22),
.B2(n_24),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_26),
.B(n_34),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_140),
.B(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_37),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_73),
.B(n_37),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_45),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_92),
.C(n_107),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_150),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_98),
.B(n_74),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_142),
.A2(n_170),
.B(n_155),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_74),
.B(n_1),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_152),
.B(n_35),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_145),
.A2(n_121),
.B1(n_116),
.B2(n_114),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_146),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_169),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_102),
.B1(n_86),
.B2(n_89),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_156),
.B1(n_157),
.B2(n_168),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_154),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_23),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_76),
.B1(n_109),
.B2(n_72),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_132),
.B1(n_137),
.B2(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_160),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_21),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_35),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_108),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_121),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_85),
.B1(n_26),
.B2(n_34),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_108),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_20),
.B(n_24),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_115),
.A2(n_45),
.B1(n_31),
.B2(n_14),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_146),
.B1(n_168),
.B2(n_144),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_114),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_118),
.B(n_113),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_183),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_182),
.B1(n_192),
.B2(n_28),
.Y(n_218)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_187),
.CI(n_36),
.CON(n_219),
.SN(n_219)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_196),
.B(n_19),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_121),
.B1(n_128),
.B2(n_113),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_128),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_186),
.B(n_197),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_150),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_201),
.B1(n_0),
.B2(n_2),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_116),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_190),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_143),
.A2(n_45),
.B1(n_36),
.B2(n_31),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_204),
.B1(n_28),
.B2(n_19),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_142),
.A2(n_35),
.B(n_30),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_21),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_104),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_36),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_31),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_200),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_149),
.A2(n_35),
.B1(n_28),
.B2(n_30),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_154),
.B(n_170),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_162),
.A2(n_158),
.B1(n_145),
.B2(n_160),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_141),
.C(n_148),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_210),
.C(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_161),
.C(n_165),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_212),
.A2(n_227),
.B(n_229),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_171),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_172),
.C(n_36),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_172),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_218),
.A2(n_220),
.B1(n_221),
.B2(n_226),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_222),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_36),
.C(n_31),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_231),
.B1(n_186),
.B2(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_36),
.C(n_30),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_192),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_175),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_230),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_19),
.B(n_1),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_189),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_9),
.B1(n_7),
.B2(n_6),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_233),
.A2(n_184),
.B1(n_178),
.B2(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_248),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_188),
.B1(n_185),
.B2(n_184),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_181),
.B(n_196),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_240),
.B(n_229),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_207),
.A2(n_183),
.B(n_185),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_188),
.B1(n_205),
.B2(n_195),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_241),
.A2(n_233),
.B(n_211),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_205),
.B1(n_174),
.B2(n_182),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_212),
.B(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_217),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_208),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_249),
.B(n_221),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_202),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.Y(n_267)
);

XOR2x2_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_202),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_226),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_254),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_9),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_214),
.Y(n_256)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_256),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_206),
.C(n_215),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_261),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_216),
.C(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_225),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_266),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_218),
.C(n_214),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_273),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_0),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_276),
.C(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

INVxp33_ASAP7_75t_SL g277 ( 
.A(n_275),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_236),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_292),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_253),
.C(n_250),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_243),
.C(n_247),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_243),
.C(n_235),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_284),
.B(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_235),
.C(n_251),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_239),
.C(n_254),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_266),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_279),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_3),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_305),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_265),
.B(n_262),
.C(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_268),
.B1(n_277),
.B2(n_270),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_302),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_271),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_262),
.C(n_273),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_4),
.C(n_5),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_2),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_283),
.B(n_292),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_3),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_314),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_299),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_312),
.Y(n_323)
);

OAI21x1_ASAP7_75t_SL g322 ( 
.A1(n_316),
.A2(n_308),
.B(n_310),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

XOR2x2_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_314),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_315),
.B(n_294),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_321),
.B(n_317),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_326),
.C(n_309),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_295),
.C(n_293),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_293),
.B(n_4),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_5),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g332 ( 
.A(n_331),
.Y(n_332)
);


endmodule