module fake_jpeg_3862_n_126 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_0),
.C(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_17),
.B1(n_14),
.B2(n_15),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_28),
.B(n_25),
.C(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_37),
.B1(n_20),
.B2(n_19),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_16),
.B1(n_11),
.B2(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_13),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_28),
.C(n_23),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_55),
.C(n_42),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_51),
.B(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_52),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_27),
.B(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_39),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_26),
.C(n_32),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_42),
.B(n_39),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_59),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_44),
.B1(n_49),
.B2(n_33),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_74),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_67),
.CI(n_62),
.CON(n_80),
.SN(n_80)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_43),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_45),
.B1(n_44),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_35),
.B1(n_43),
.B2(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_43),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_60),
.B1(n_35),
.B2(n_61),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_48),
.C(n_32),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_85),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_77),
.B(n_69),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_84),
.Y(n_96)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_76),
.C(n_78),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_18),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.C(n_82),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_74),
.C(n_79),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_84),
.B1(n_86),
.B2(n_83),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_5),
.B(n_2),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_18),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_20),
.B1(n_18),
.B2(n_13),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_13),
.C(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_0),
.B(n_10),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_10),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_103),
.A2(n_94),
.B1(n_93),
.B2(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_107),
.B(n_100),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_113),
.C(n_108),
.Y(n_118)
);

NAND2x1p5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_95),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_97),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_117),
.C(n_118),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_4),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_7),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_111),
.A3(n_112),
.B1(n_114),
.B2(n_8),
.C1(n_10),
.C2(n_7),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_123),
.B(n_124),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);


endmodule