module fake_jpeg_8533_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_2),
.Y(n_6)
);

BUFx16f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_2),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx3_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_15),
.Y(n_25)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_13),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_8),
.B(n_9),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_7),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_18),
.B(n_19),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_0),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_1),
.B(n_4),
.C(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_13),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_17),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_26),
.B(n_27),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_31),
.C(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_19),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.C(n_25),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_32),
.B1(n_23),
.B2(n_27),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_18),
.B1(n_26),
.B2(n_28),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_26),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_36),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_37),
.B(n_26),
.Y(n_41)
);


endmodule